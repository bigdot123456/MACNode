`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xt0wYsn/6fbWgi0rcu6s0lgJuPL6i3wa1sSA1WUPIYIhViX5ilE0YO1v6Gj+lXGN9UHZ9rMsOuqr
5+TQKKHmqw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MttwRJ/LALdvinGSt+dl1xLchlNnj+9rZbGEoXfSjsdj4FY9ArFVWoH7La6DbwUvGlc8rU2ExXAR
qC4YnDf9WhoM1EvGDx46vnY3iEIGI4SUwSvIWehzTuhM96hE3STIIMrplGe23MqJOQiWHe717LRR
9aCefpMwaZ5QVtEr14Y=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qTjP/9EKQGFGCkxYTmYgbEE3rQ2DvUlBREwY3Y4SYe1BkUHeSJHFIKdth0S+wG3+yGHA4qIlXvEo
cpB2KUs2W3d/i6VK9ddJ0Zzf4qefbCT0q6FDQw6YK/ZFu58DTVKyQKeOFV1FGf08rkjFMSEuo4iA
OUiMizfbIqZ2ottdb8BobrSS5vk+yMm+S/Cw527dtx7McN7XMi1/hA9Hd/0pLXFQtvw38pPcZEuh
XSUnZCola7yPVrgVK1ekrezImxAiH2WhQNXatmaDpqmV9aEwGWEYlupZTYcstIsIdtgA8dOD5UoV
2Daga4S1L69lRB4EKtAvVX5uoN3sOEOuUN/tWQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ezRXVbvbBTrGkGToYe+fJABRb3pZc4QV3hOwosYfIu5n5mFnW+J7bSuvgEPCbXdbf/M6lYh9t7SH
a5VszFFQo4OGMkZXi9WP+o9bkbquuG0vaj9FGv7OWK/rHyC2WBE7yFCQ06xU4oPMA7Nc1+UZ2zOB
ScDuhzzFqnsSFdAdD45aWXGU5Ao2398hUeXfoJzYU+1dbQds3Zl3j6x/4ykQVvNL64OOQc8f8OXs
Xr5VfjeV6nQ7QoRYRHBaodPjMbYo/XwblLC9hq44vJxvpcUl59i+gDSp72WZVPYnDeax9seQNJR9
TEt/uGD0sSAhWmxi9eceM++JmHtweuwVEMvPbQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QkIHwzuHGa2pwYKKO/dfwPg+/jaJw/AhvO9i02+CYmlgbpOAygYY9f/5h5WAdkDuV7bGadPJFKWr
cGoWmQdOgnSJtU+Uh+3FrcumwE7Q7lnCOBh3Awij1E5NJa5oIyOXzLWbZebQ9zWfNYbvc/FXdOkl
Py/mojjZbKCpdb05hbTkUgWbNj7pQ/qXN74iQCTByhIgXLfv7zxCDPZ8oGg1sbiY2TlqGrzkvfVB
yb7pdl8XYCxYR0FNJYEEUwpOjeDBiTbLsE5lppfPrTzHLv7fnSJAgo8RZJrQcxyXZ9DYA38e2udR
gGqAIiS7/l+Tsst6Wrrem/ODNL/6DRFt+oRs6A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ktSCUKMz98r+/gdhtr3qnXHmjqvUL1LEQ/qtNXkrYj5dqH0ZaMSVS+eJ9RSy+hE4CSN3HG4fQJzJ
WWSnikBQ9NOs4p14CYs5/x0DfOyzNOdlNNWnctXJDEjyINpmDOdaQsjs3xdP//OarFBdIBpllpwx
dkEh31aj9PT/n5Xa8BQ=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cBTW4nvIl3B0gOpjT7XQg08WgPz4imwj/8MtM3x7T3NqiLgKiQQzdGX7INeYPb1+30E64wyv6x+G
J/ZZ1ncPVpSUKIyIGNE+9ssNr3Bdo/0c2MdsEzrKgD6Yo4tP0hH4O3Qw9HbnZ6VPizRxV/m59JeC
RicHdeU7ucwMCe3Ks2m61l6nYW0Oz/RVCIR3pua2g9rv+p6JLb8bMV/ejshxiSet9ccKTmsteEq4
WG3Flnx85GPOvEuWk8zbW1tFPVd7uTUaUFSB2+9XwrVV9qYVCgAiLITe+fhhai5OEruUV6/O/ALK
hHPUIkwugRDpY7bcTDSRC8WBa4gXpu/jGLGzRg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Wzig0NT8mk50CYBIvYxqOTEK0lZ7HDov7kE3SxkChwfoutr2tD0hy6XMtSKNhnSHeNImuvYN7ZxW
+C2xB9sjbBJY8ANkftxhYDz0WI/TsRlh7c0EwCSrkXhJro7gP8CPqjVGu1t+BnXwrUzd9uThXNON
JVW+iRxnwRC3xVjHoT2yQe1AybbKoDb9DAJvsjPR/vQO1xPBbNFp+EZPpRWXRrML3ZWa4lP3OzUn
CbDO7vMPiAc7hI/ZY4x53AwWtbp9yrXaT5ThAESnVfC6hG+kpjyvcX6sKbBP9zToEeNmI6UntGdN
mv1ZMe6KfbVajJ+BcpjKz1z9Im+kK8ovmX+85A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1167584)
`protect data_block
VMmFQmPQaQ6KvWzZoMQ42AAfNs3QGhZZwBNhc910esYckcvkJ6zzCPL2s5Ss8HbJKTBPhFS6Asg8
1O+kcRTaBU6YoYcfcDT6ZI6z/CUfWKmMRXl6ch46KFkeeH63gnXOr3fzjY/CWavC55elQBwEotrr
77+Ey1ojOD5NJSt7V6XwR4spBWbJYOw4xrHtvIqnE01Dxj2Ai2R8u/NAUSiEjXFDvP6b5HzkU49V
q9CLoImlxkwIVWbaCpMR4K2I8ClNd0qva9+spBvzyzV5/KTOGhD2O3ML1FCoVOxvkFNj+qKQhO47
7eqYb82faSV0/o3dMYzNds0MEVVh+pH0gxkMth0cAUDyuEDI0X+jRyBrZA+P+Diywsp9XvpYqTxn
Blan1mc2AAVvvAyE40wRLGym6CqVnOYstCLYn6pTSNQf4rpfR8xjDs74apdRLxFCF8/M0CHZCA8J
53bRpB87QLN6RDeO1zHqLLXFQO/MzVpxy2BpQ5rbJshwxhW/pkN/uRLRQDxT2IwrtCuSFZVwyxSB
Q6V62bjUe9rERRwDzMKoHO5WafRjKqibBIa1X+Ym9MEQQtonBt3DoKg2EnCceoRd1Q1xdhXii6Wv
yshb6+7V40X6KaV6njHjA2vvG4d7Whp2QhYoLXae/+RQs9IMOv+fs0X1PODyLxVYXQfvrE7cGYlS
oPKa4PupwEjKrwfRrfDj0GU8REEfocxvAOQjwh0appgx0PkSsZvPHotkIJQ61coqhNri4/HW21jP
kvkRZ/nwFd6Nf7QqDXP5bUyS/8LsvwY4HwF7NV76b6u4rO/7TfQt6YHScZxU0zB6zuCDLt78+3bY
kV5xqOpCqy7Mjl7lAHZ4ev9muOOjYcVdl+vwDud19Z/uqn7Grho5FDKIHfXWQ7asb+13BS6357X7
3BawCnj4nyAP/tmNd5ppj/CNGslkudQO3fl09C3u/ihY+kXNPPb9QKmP7FpOZmkJw2znuWMAGGXe
ApaYRyW0sN6eTqxONZUtsPLv0cbZtTVbDlN4p3BCAyNtwCJNuPnx2pV5z1mcv7JswA3ziEgzuRxo
hlBoc3cmTrZAHJ5mVYPYtYFDLI1/XUq4Qo/5vC0RrtmZwd1qk7uoutlrMUXPNjKgUOeFyVcRTLij
0DBx+M4/HbORb5znZ4iLpo+85WFMLitl1KcGu5zPuFdnIuPuUMzBpfAAAZZ7cB56HNYKNlYRIKjU
2DMpJYpKhHAxIJ9yZemzrfaSx0xyJ0hEoEY3GPxKqw3C2j3PlJQ4HORyCaNR8d5MqG94Hmk6vEcG
ZEspx8Cb3DlfyEzMczlPcrIYiTmSmVgP3ykA8HNUa37Iuuu6OPwOfKmNKj2l9HKBc9y9+SvewTGU
2nkc5lSvPH7TiSl2OIHzKdfEVw55CvmaChccVz2JP2H1bfzMibVPKuENLTSYX93opGI36UrO6d56
cdyA2fChV8KHxRB4R5LMXBAdVjAyKrHMrVidS4lp6ZCvL/CfgQRWLX1m0eju0fFOg50GBgXi1msR
TyxAkucg2/5FKPDEKTzZXCzs3NTsY39InCwxmC8eE907J2/e0Ia9RTKqQYmor+lbL81uI8H+mz2A
sKH4YzumRqbP/mpFsAZE92P207Nb7byT9vuFUW2CGMXdtABZJjVZPZQLAaag11VNsRQvM2xBicDK
Me8leSoJNaVy6xxpwrOFFefescOH/vQAyEqVjOtRHkJxEYexSX6gpc3MZ+Hr88nBOS7R/ugYmfVN
5fFZOQzDVNICVgnNwKo1g+IKUGOqZUiN+DpThZNv/tarKdoSdgfCfdlM7aC5T10rEKEH3H0MLVu5
ZGSEE7D8kUUNs4ZBzZv+GMkG8zF9Nff0yjdUlQGs03g8uxr333WqHIJna8AfJ9D9gCtEJg6CuS7n
KR3fZz8lCqNy97XK3xhzTYuBret2mPJZHMg2YIEymu7l7YRYf6hhxhf7AioXU+Pk6zSLPy9XyNGB
loprWCub0ke4378YYza6zOJyjupF5HLEa/SVLKOUMCg3vEpXHLyaIYhhOOtD7og3CGgPeaB/Kj4f
j24Y/eDFaHQcoqlWWWJQkLAqo04ld3IjipR41RfMsOg7s2mfdUhcn8EAFdo5ht0iwXQ2xmeRxMuz
E7d6G46VWuGI4mPPZQFUICFbWhxGW5zOZVVOejpSus+ppJkKEUF/TwcR4oWmZ/YTbJd9ohVFZcBo
zHAhpJVkskeHPrJsDpqLzSrid0z9Ll0sgr/C2mKxL3eI66kBeIk+lVHVB3vUOsrYNXpZ3QERtVfz
iBXeurz+nH2pK2p+6/8CxmJIJ8CLxSDQkSmyqODFfYWGrvuLdvmL4azVjjyjTcXpGiLtwYhP+W00
Boi1qdzOk9gs3oMPsamcX+DVDIJaFYkXSUkfDPgKqzh6RBXWUlXYI+ZR0DKtG/GZB+Uczb5FGS5C
sjxqPfkFQm9kaxvm5C4AUaM0bb0gOanqMNDOeOVIYF+564ockr8BpllSh9TEiSlk2WQhzF7Kw1rZ
vD1oHJq3avW7fpv/EDBzaEXjNUjgDDUgtsxKqnJpBuA13wJOuxBhP+kHEmJlBcuLecGUtZJXP5SH
rJn7FIQe5V0LU0ngQ9R1PGGvRO/UZVvvagYmuj0UrgsTCCUYcotKeodqmVL8CHYcpXpFo9OqbW71
09eQHN+wtC5+LBIm3AMkpPZEpQK3ZknmTWkrOC9JW8gfd1wuPPXpXvF+Qp+gA2AjeA3XXvlU5SUX
zsqPM/TZnMRvNaGnKftz3nNSf0eYQYWgTzRK1LZFlT7BCerYqX/W6enNRfnRp78ij6nK17FD0HLj
7uucHHYcjLvFf28exWneDDudsryjFjmEVbFiKSzQUjaYnUaAPE+o3pxwKNlid2fhEFeLxcVmcaq+
jeyxxXKQ0s2EcXQWJQuCc9zF7c7Rtup1nU/O2i/cPJCxV+dNs4K0f5xGx/MrbKgIh9lPIcGCnqPh
ez/hJ5k3Xb/CT4xoh3XRopHXglk//YLF3N2ADZ0i8psh6cQXqVF1+T40D/ilCGMdLvLwkRIUYZUH
O3f8iXihorq6l2LyNwXdp+amDoazfU7a8C3tgJekZHQfUo5HLVCxaO/OSYGYGguJyAhIXfv/VW3l
2rtEb8SLC2hQb/+LlA3kzKPhOB9gs2bZ0VpAvdMBNMw7aOiZC49io24eM2SaDvYbSYxA8t1jXSK1
y770OgYmhEaYLHda3R8n7BhNv4eGr3aQpLgCEv6fQ9MX5yE1MBmudgKTm5UahJVK8qXBj4/iQoOg
rIL9kC1ko5x3SgxS4xiKuvV9S99tztrfOi3rzmhTVK0Z+1Tck+sDk6XE3GP/lZ5+pGaiNmeHsOD+
ZjinrlDTk6cdNTW90O1a/DwMBjRZ2RlC8wnmFB63kP8yHKspRuee8d1NxywawWnze182XZ0BuuVc
On7+w9K7dhhctzbKhjNvtXbPMkdJoM/G4/H8QNR/O931or2uOa5jJ0SfDYCSoR6jruURe63iNWyD
zkF5iLgrK//fqcXF+Tf+4l+5HbTh/eEERB7rrBijcLmaa4RogZD9+mFZbixkGE89F/3ASROeywMt
5RY8tl2Gz0vG3rMrRjjyjKKuNLFXwPbqvpz8odpCFGa5zNLWQbz2YFLJpKmKZqLVBoq96vj0fdwn
9gjTGanzmdUEWk93tBssAeciAapzCjO5J0M1XyfE06Yt2gt40HUjlqIZBetwsWfqEYXpOGfakxaM
EQ9TE4K9k5M89YqlJiQaIBRspJfgQdSYUgkjvY1CcCGb8G/YmA4ViujjFqm5MGSzsl0meUjZ3t9S
vod5uhiK3Nc/uQgAFlxayEBou7K2Qe1zwAjC0jVU8XR9NC7WG+Glomj/EHJH+VU8uqEoMobQdytY
xKGZlBFj+HIsJZmkiLZhflXvVBR8rM5h8uFKXEafLLBKmHhvo/4qzyf2htOplWQ4xiRKBQQcxIkU
xTAQ6+h3dJIA3NoyTuSgn2c2HyNQB408qOsEz0EylYSmRm2/XL+ZmCChp6PoTiy3MqrWQ8n26vp8
Jybvspi1CzSCLxXzRHLBydgRtJjXpc6qPWCCmMUMldTq9P7KB3JS7Gt4z2GiCEAdmyHRe+o/VbSo
ZbLB5qS6Ypz2KCR1NgBHdAYxGku909Ijw4J8w28iVokM6xfw7AB0AN+03DkY6PUOotNXHCoOgGc0
/8bzRqlFv4O+BLmyhM2m0LSAHTa9C0x8aVG/LwfU5oUaflryEwCOZCk/CYA94pYGWytOJkJq82bZ
jlSklX2FleZWlU8bt++F2b5YS2F6EQ9xfV3aFit0jwDnKt2pbKah/1t7Jg7HX2RunB9RmVWFWSi0
j94J5Fxk+QUV6FjGkWk1nEpg5zy9DiwdGfvhPEnBCYpTRLUsrY8MWR456tADrzw8H6tJN6ni8ncO
7mOW4xAef4/f8amu7VxbmDCZFwrVXxAUnrMYBy/d6YVdMTHQSUXI/W+bawpWbeAMGWffELDNaU9e
aJq9+rCK0zOhz24qiaHoCbOE/UiDKFQlnhTD64C2/OfDBzt9vPV/IVeftbpajzGRCnCFNsMVX7Z1
YIryEvHfZTf+WwDB4lcp3E6bRNknCtBek8fQZ3H19/FBxsguPhLDaa78wAALbclfiKlW/IlDC+y5
b1qkLMkcpmGLM63vBy8Wo1qEf56MP6WwHMXzwhutzUNNNxqpYqJ1zH2AbVkEDcLNDd5IQlzxceWL
SIonWD4f4iG26JqSTAav7jFD3NhD+FIPB1O+0piAQ3AEQM5qeJfudI1XqCvuh9klMn3R10jiJeGd
PS0hyhYxaWDoiXX8tOnTWX1t3Ix+RV5UhrYd9ZgJ9YXIJ0R0PZLJkl3VLMbLveoF/yd28OhENgmZ
0qGUUQ0ZlTjy1qn1FbgYvJeLNnBM/8xmq++4ipkdf2zQYvnY8mLpoCbi5wyLpa5w3CkF8Z6ON2Z1
Mqo9VuCPZ7+su4ayuryVXPKKjoG1aF/wOE8rdV2cQOgkmP5gwScy2fE3o050dhtG0PGiTjyfOzWw
5grQpLEpOaPDo1jLAnhDTSDepgJjSljbXm0vKlwH0trbAkUOe6kP6idWToUPUuNt7WxSl4t4AVqT
tKln49t8vA+l05YSC60LWABNqsbKI9u1KJndjXGoMD07dynMx1Yxe82oJieKi+585O2PAWgoxPE4
GQ38blxNgdTgdma/hqEyxw6Resitx/kcKenuVY1UHxn8ArDnhO7Ge/iNvum0OYEA6w/HSF/scPqx
DiBrWncRF0z2xrihUtf8r30B8cJ6JqToY3BYtWLBEuqRRQWhyiaeVU9YgTFDjh7MSIm1f9vLcpV6
s4jo8WvN5Trx+fB6KhwWlQ3ZUzy/uMS21a8R/6ohhOUi9Ab/Fzh1TJd/4K8PfBty6Pbov2swml6z
E5mqG05DMCAaueDmcY7PL+5jm08vvlozhOEXwlqFDnUZsw0G6PLMGft5NteVWbBr5VRcKytwua1w
WLY624T+8XKFMaP23v6Dm5d6FazUOBjN97/mxpKF8JAnBiHVeKDGNbJ1iPyHbnqlNkWWSo3rRgqn
wYjnuCvFGpMaeT1ORvZuJba7rOqRaaKo2B8ZkmSWoklnd+Au8iuoBvXY89zZYV3l9nqPU+AfFyK6
WMHYh3hJ+SxIYMN7R40we0gJL0ZJv7H+DZvHxneyHIUYnyIWRHMSzosWqI/AFHt2nGPaONk24vhW
3HKMneT3jP27V8GQjwS7J6dmf8X9MKwLyLcQxMGu8ZX4Rh0txNBas8CvKa/4GkPJIMafuWO15X4Y
fHpK7O8yadoIG8jQdDFm0pjpVgS1MOASLXn/ptobAjg7cmdLvi6DCCaX/MDkHfIQVNw40FPz5lRR
LEtCYM82sbkcX2GUVliePPsFZ2WUk1cCymNwQetdirvcZutH7iz3GMzZYRjLahnnG2GynNHtKDC3
DcPK5qz77mVDIG+adSJ9fV8Jta4uZAp8B4ff2B+in/Ibm/JJPKTCsK0w3bdGkFPpBfLg15BucCzk
1jg8haojD9IKwPttA1UgRZ8fYyYIuvRa79yyLfMP3qKT/9YAyQV/pU9yrvGKpgJN4Wc1TZQLnqqj
hE9u1yqLJ3HumWeMeECzKmo3u+le3FBErsZEJSRwt5JcOEKRvBlD2UJipD3MsFWFp3+i7pPV4uhX
5gtKHfVKwdynlLrGw2v48E4PumjTZ2TM4lqWg3euwuPxRbMJ/g9dRcP6ZeTA1NVuRxsFOwMv6ssU
w7jV8VjJxqOoiTzYv2HkpYmB9Yu1tcr3DdmRsTwLzKvqT7SIrdwN4WROFGSxIFu+ze8Ph46DQAnz
vOpKnRp6fvTOZP3gNcaLG+FdlF3gzqFREnVD8pEdQ2Eluts98ubioDp9N7D818VD33JTQD1S+H/c
60PZsMY55XuWnOgJ8K+xIBaD8n/dbgOvbObyLmibONmphEXhrTiSRCsEqXXJqdRllMDd644+X8Nb
KaLTwBza3JgvlK5cfTXKDPdhWv6awx9x1NeWzG2Cx1ll5d2M3mIIsohS6YE4kSQkOxX/nTpxUTPA
pago22la2sIkLNDrpka9ufYy3pQc8eBLxPHcXV7ymgshGTHbrqisARxfM0Ivf+1HQvVwhgpvbJrX
ItT2VNg1VQJjzi/guuuVns0cZl2NjYbtMmGZbYnAcCPFcTy3GvLtx8FKnr8IE8xHimDZUC2ZBCUA
urguvTcXULQCXKWS4GmVitASFjMSCpD6Or6OcF2IqKDxsQnABbxoZGfxPLg/F+erd5fJmHPS85Yo
W6jEZCNkJA3YY7NQfGu+YuDARrXkhBnxGlU/qGv853Mg+6rL+GaxEJTw60zLH2bFtAtkmG82MyPX
D/IRDHAASj1dNBPgyGytNC+WWG5TkEWD31ffdth2aJJy4nHY1H+j3Gmd5J8z5mpqhqhq/Tb9Mg1Q
6lcWozG8MJy86LGimnJ+mu+ZbVqaVrOrDbgUt59pr8STLLmUVxS8MH6qdNuzfUllRGQr6jJr8Fy1
tgkuRVcVfoOFU9Kc/x+0usmOA4isdCgXpvbl+xEZtP94jrDlL5t1JF7A654G8bWr5t9PICqLObYK
N1XLNxQR9Z0af3w9hvMebtx/Jp0dJvZbrFujL8nYFNnH+rcx5P/LuQeK4nvyNH/nkJ62Ki0WI01V
V0p2T7NHJcF6awGOlQHhugn/RXYBgFZH9GN54ELAkdtAUt8QvjI8HxN4Fbu0oVxCo31Hx4ZIJEi0
kA4+v/Lq6f+hNE4BCcXLLKWqdVQ6OvFqrjb2EK6gcR7xgdWLD2VYmQMeT8+xUr5LeZ8VVak407p3
m+Qj47BmnU3l8JbnC81T4ZCS5F+LaQVKz11uPKzK+bLz6oawS/EFqQI1IkV/qM+DNtq7Wfq+UDkN
Jv+NNtIISo4PNAo0PNcpkNxOBcKYLz6TRbyWFzcX2D+l0FWS4jBSS+UByK0b26Fktoi3RdAmrJs4
bP9fIE4RH/yPHyB/0ASSJ2KAjMIihA1FtWcKbJW+HMu4+qi6gh3lbax6rpkGe2x9xg3+lLJZVdzr
lnpsteso2peZ8REdA1a35/+TBDBpBYtoujlYH5M1jLLrN2RuBRSxBLWFueje3E2pwrFoHAmnBkn2
McwPGljFb2nHCRJSkJ951St7t7kkY/7KrvPyiMDmoT+QgGiCHgf8S8S0xJsJr+aeLUO/9ml/fw+x
l/x8yr8vo4RqQEi9asYml/xkQ/5sb7NFa327zrLWBNbtoTZ7qseKJUEs7BD2CEzcC5ROnL4Jh578
Yz4SFGcISemoHvBXsZm/n4TNfixwMjI0QAeYqBzC3DLm0d3JYuVWldEmpl+Yyn7RZaA/M89xI59B
ILnAS5KwrIyzcUGEyL8ZfRt2kw4ow6jsZe2qN/gbHzbYfpNKS3oQPVx3uBPR8To2BUt9PqQQFmrf
BBJW096rwV5MtUhZOkRo9MQJ9E6ITfPvun8VQGtLAWIGTF5/rYb3r4dDKdq0xfIvNH6e7Cpg33kP
sjverHqjWiyTN19Rc8KwtqUfD5KroXvRDZgu4H+6a6TfoMhNUWIBR8MgAhzKX4GhoM1G0c1pqfLk
/slrr9KroGqugPjl+VjuPhAu3g3fAInOoOcpmIBDcBaJGfGr8MfPptt3ZyhGy+bhziUSM+S1ehDE
SyvaNMulamCQkkPlWTAG8l2qfqMy2VfkkF3iWu3HvSa2UaFot/LOXLnI9hL465yQnn3pCxLCU4d/
dyl5pGvb4jLWJmqOa12PTEyC3xacnTH2/dHyMgZxM+bIbqSu+HR08ha7+wNo7k8FSRkNiZ/cP6X6
1I76slYA3akUCHfB6u0iNqz4hQr6ZhKM4fMacVHFTrxCQbA/ifmxdSrlrpFY8gyNc3M8FNZr8lqa
VYEMkBi1StZicc1cbHTnbD1NVwtJ4sxj+K7+hJSi5eMrAAwjMNWleCJwWcIV5QJywDvhN5O9T9eC
uuIOWVDFK5H0gzgGG38vCUUVudisZrI1+NmvBErepYU/k9afumVgmPGfWkw9NcVOiTvFcv5/zNwZ
PuIomi/CIa/GaPgIEwjL56uP1HI8GjXbHNEd8S0VOpsTqXxwNk4W5glH4QhLX2f/X9YftE2Guzoo
DlBfMkLWMbd8lFqTBenUMit01s4rF/9bPR7wZi9hvSScOKFjDMof5SJw9fa9+xnH2RAbdMiJ2ZCv
x8Nf/PQgNdO6pAhbtbqTQu7eupJ/mKoKb1DzDXGhZJnEfBcUtFWct8HlggWi/ceEi/a8L19a2TjL
J6IBl2rnsg6Q5ka+yD6rFfgWeeoV1Mqgg9UzQCxi8SuYGLCEky5u7mK4VolkfBOufQDCLDYP02Ej
QgSdINjnjgz9R6Lw1ujNxsmjfV3JUFpjlINAPsjhfC9W7m7TSljYfcAPhDYV5JrUgWeiwK2h09dC
y4BNB+Re+N7Xxc8utDOonUM6i9HvayDL1debuWcBzuR6ncWsjtn3vb7U6BpIcF96uhb5ptT6/Ffk
xCtHSg+77T3TcK6045bThPtFVTHZ4dG+4UW+KbVE8q4EN8csLcaBcUKR661Vfzo4l8Rv2yWhyJRE
/9i1bHtXX6gzj4VSI3/VoNO8G5qfNYth8QWRPpDPunCY8i7DXE2+jlLA56mKa7iXaDF/WSpuQGN3
X6olLxIjvL61b8KuCrILKoKxqm959hRfNEeVOotQzNIohnWSYeKZn4yV+S3z9+CFMZF7ycuaRyLQ
7FDwYt+fBFnHpPJD/e5fXRsuAoLtCV0Xv0l4XxygCDytA940kgdpseWfUSRpPvgOLWaAy8s0r5H8
SGiOAEMmgWV1YrJzkplNKg0hcmf71o0oHOb5j6xO2tRvQlqKGNhpAspBBUg+fhVpNVrhTk0dPWPz
uIcC6YVDHUoRTXxbf3t04BoRsL10Of8HXD8Sd9AwBhDXEjMR07qM4Zm6eQYZopwZXw32dGSokb6T
bjY0roBDBTrYTh/c4wV9pHAyC1+/ZGzZPtLFDebbRs9D7bFPNAGJp0GG7LrtBN14druWspuE1ffY
ybd5STtROza3ITljwbNrQeH+AF230mBryIWCtUIPtRpQwLkSKP6wPqKtyTG3FjULB4znDFLD7Ohe
QTAZv39xYDWKEXSpAPmpsRpdIpyRgt4aeY6QBO+OQN7pCAeoL3PHGZKBiMcNOylS8ovUI4ElMDl2
o2aCoZzbmLIKypMAtknyehvF5QUGo+yuBXMXM5G+ki9TsVrEMKK5s+OQGSekMqrW44AlUYut9SOB
4c/zyai5laxchfn4cETUNPGQiiwF1CS2lCnK+wFp2eFWc9PhdqM3dk9ouTaG2U9QUR97NIoN1mN6
16FUdrS1EddaGvt8IhpYCL3WNwqX+YMSIH4WJiFoRL1lD2VREktnbRc7+cWbREK0MMUuTl8JuuNN
Pqwd+a/0Iw6LA6qQ+/EMKzTCI9Ifj+/tssyGP3GLYD2JB7juidbewM4qf6Dfm112ZY75U1I2F7wH
05Y9ptzQl/ll8G21On3mmf2TRu4lnKBm7gTe8woXHUGl/8KkXK6DPelqcjH+47RyRz+ffS8DsHEk
AWuZz88pAp/iK+t/9KAX8VftUri/E1nW5LFzQwU072K2b+B4vy6zgYXqR9sjjgcxUpVo2OH9FUXQ
TnwWcPjrMdAhnA61h275ZLu155I4GvBapF/8hLwB1Y2wuKvqpdLlQsTX9oSacvGXcIdAKLDzSaUF
5w9lETIbMW//dchoe18vZmQ6OP+UGRmfw922txqqPvOmkxKwnrIHNQJ9HUOQMtchz2bZD8bInnuh
xcJSDUIQxtR5UfMWl6TJ5XP3ICDOpe3dWX/4ltCmm+f2FN1xM7xW845yK0IH7BEo/xNkHcaW9noB
1PqYPwbDLx5xVzZwjwFNhBDnJOtZBOqn8Lcp3u3F+VeLlyt3Odllso6ClcHr1exDJ3+NJG3C7Gzp
mXhv2xcQ4ZHO6y3ypVq0uVRec3dbMAB7eki+tKjaU7yhFr1L0E12/2Qr7aZJOCK6tbbY/nAljvzd
6tbchSAVc0b+r8ciBTu4phlq9ZHEPVXwvvDY21LPvwmND1HgrlnEjtu6MrIzmdwxhuEwMOin338H
DUDccwj5xcd3SjMBwX6hoKalXaG6J9AMEVXuBHquhNymgz9lWGYlPRbjVF+ckkKNmtBdDqjxHCXJ
hhdPnAQtnT4RJG0IsPXiLFY+1q2hDf6o/BwzRAhdTOB266HMg4ZSIc2EWSq8zqUS4utPrDFDUETc
31IbEph3a+tKNJ1j9ahyytqiGvpXGxnEJ+/VCQ0Lcy9cVch+Yau6S1EFaVXRliMWDIjsgK7Ov8A7
40xl+uYiKMoQWy1VSAs2lVglrKAMzUMf+FkRJFwhLzk6RwK6LpXQXLMOfteIpgHzRkTSL/3IOb7P
WkeNDVEwKRLrzLqHDTYJFTyGtBtA6B4cncztjwnvUP9qYVxe/rXQpIuTD3QN3eWuCqfBf054vZVo
WuzIXp6PnCp/bO/GAWse/rjiCR/xrR0hl3Hajw49QO6FRSQjO1ybtRwot+3oMsItadj7h25eICS7
2mPY5rVdUj+Hjb6cfJfacQegFCGmBoHtXdK/3JUntcIb6d5yPlX/pCmBZcJ3ghLmbE6imnQh9/HM
XlOXqrhj7eoIUPQgBBmVvpc0OEZzSDm56ZHOa3YyFT5u+q3pt/mKBZPq/Ob+Vh58rJsfGbra4uMJ
trzwCoZrs8aSNlayrOBbNQS126WVlleQt7hY+GjxLslCjtdcS0m0HUvn0HHImThFgJyGMr58j5rK
ticYGC1NRedUxiXgdu9LS0+xUEAfvcBgVAqrO/EYlVD+lgXp27l/ejRj/WWoMmpmkPzEfudydoJn
xkmCd6kvQ7rkUF8GM0CG5ZGCTQ2svr5K8Ddz3P9QGmRZq2Rm7uTdpm1rVrDb/CVnOMCVSTW8uo/y
LCHLY++Du7U/Q8G8LO62sdfXVGw1Yq/XyyfKCkBub8BwZf3Izq+zs5Nh/8h02jWAfclVNcrcYS9/
sH5P7+6ZkMv0VcQ9Hxprt2VY6Ix++ApVp9GmLoBM+q4/i1nqL+tcA6etJe7k3DJ1AhPbiXkxnbDV
TtHxpAX0yjyo5930JlXJwcXRK9LCvrV3u5dNM4XVSNosLtU6yiVVvdZhGkBTAi1c6nXYvFn/MLA1
4DOCh+wqk5kFIEptHGiPAHxzROAQ4fo5kGQt2H0lwDKhX96rN5qMbXSE7ehHuHPJcGTl17rXhaxy
PN8oljFr/+6K1cNBpKOTHBHVBPEqjJbcZHYCaMM7dngB9lzk25keRwYitSik7SHTkgdOphVPfbyA
BZ3Zndo/nxLin5pM+w/bEszIu5bJmoSuMQcdSoFhhTJoK7YfN0Zklph5A/QqVGTRNb0io1wnfYYR
4ZHSBeZJ1zopo+r0lP3Ro4PBd1uJABsObcGN/dN4fLGMhKfEGQeDjYt/P8eoopN1ABYylzubGqVH
zL8M34Gu7R/WvnjPAm2+RxqNv2AKV0ce4/2LSGQJMUB/dgEkgkAoVIZMpM3i/QFLmbmzgwo0TiY6
Pd3K9y+53m8d98jDl3byNUrdKu71bqDdy4H/Fs0EBQ8SQJ2Vn9OWa/vFyzoEI2aA2k9c9fJMUiJR
/ZJY7030hnS3Jozrpird+IwBs4P55vAGymvmm7Z5tMHq0w7GMfH0okQTDzWYynLCaBoHeiOSBbbl
CjlRavYmwwjuLDuu6tKTrER3DDmVkFAHN4kY6Jt1wH75QndZfb7ux3k1NPlmD+bqI6/iEDlAVCml
tJrCff5m/bERd0qyjEpqzZeu3PjIaoinHTgKarTsrI+MwCatT4n/Mog17hoqxXJnxlGOjYIj7AgR
kwQbG8u2VTjzRs3d8tr1wLyoSSCWL6Ftvk2rcvD0AWvTRIPdJY5LpnrDNp8F2Qw1yYOMNIN4uCg8
zTsaPSBoOHMhr58l8wgOSCcrTfMdFdGfq/bRqPuC+7fQpjvMaKt+mVatFf14jHOzjLtrwsi/5Aph
idn3B2ivKlZuKvz0yQ2QXdNtRsgPeM0R2hLIZDVwsdZlBx8ndJRyxDwRsTEveQ7UKt0rnZUwSMFA
ppD4ib/an8RBTltY6Skxl/59Y1R09cjV9rztmniD/z0YK8tzgNIebJoPlaNK7JI9wclmrhSNfuOu
5gqz+ZrwHsclvrLl+GCv9rXbPfrzqgXwwfcCFtejhjU18e81ehcytvhglIZwkPtXwme82b7PcAfQ
BOa2snWQnGMzass8SGQRZWCL+oz0/rYh02/k/jBKhiIqaDJhqoSOecm4I1GfnrLpDnf2WgNlVQZf
0mySaITJj2k0mkEGxZs1rngzawLKXs//ioACNFb3auN0jMosDYDI0yXBCVgkF6YTGutxjG/ohOyl
LRa/F4x+HJOQop8xy5HKDbf9OwrFBuTur5TKqX0PSjNbwJBkNc7rJFHEWvXLe1NeQxxXa6lhONyZ
xibVvngFH0fr2iyRvc2XPHCKnV5KI3OpKmj3QLLqtjQMPGcmAzPXB2bEaXjsu8i+33lm6TV1C3Hx
VKqozVxS3kyimzweqmHcJ4DF1uI4sx9+j4FMzjHp/hfzwrfGoYfgH5gtiNisKSlCTfjmPxCj3VD+
wjPtDSiYyQfQyYmz1NyopxHdPpS2Bl6yX2E9Teuhv+yjf44qHLK7UrRVNTZ3wsiuLIZKftHLCsAo
AqbK0vY0WbXgpmTw/vYxbHtgmjahEyEqOD5zwEd8M6rjSOk73PLj4cIxqG4ecKm2qIBPH62RVC3b
lxjowt2+b/R6OaAem4VAI7k+wPBLJhDn1pSBjLEnUJftJrKw3dQ8hxS2BHHyIgWlasPrfkyYKdGF
gZRWBN21W8WqHDtKIC/3ajL/fQMEvEKjDKjFFwh6CNRTiOS4ARelVqS0mdOwseB+gGW5Zgbec0V5
kI3/HMZQaW6HqHjuwQyrIh/zwezXJ2adrxBrUHqhepmxaLCCenumfGZJTXQzqLYefmZku8DOTxYT
FlhHBsU3EGbM2hvrntuv6DYIXZQnfxLG9uBqE4PsxO0E71oMgXVkuoIGE5kFWVune2HRs45s/n4y
sImNlJNlj6lZy4yt4HSnmIdr7+NC1l90KwyrpWNejbG6USw/elMfwnRGunOZb0893dquqCqphmlz
jk/O5tlr7vDXirVfB8wb78wyrMGefBusFbsqMNP00s55bhjn18ygVaj3JoyzEmESSS6qKKLgn+NR
rtLjGIzqp1GOnNRnD32GdXrXOHurDEV5dvQNP3gEuiGXb+uvlanN/DOBZp4t52N5Qd6+qCWpjNwG
b9P8vyM7Jy0LVZNPGBleIXF/ztoAaIB+t6FJ/t5F+vN2y/+JcsjQmME4sdYlJ1EOJRm1CsFEyily
LFZ5pnRK+lWADuevtNfRVJhWWkgEwc+VQtd7V08N8AoIV5e4jq+3tNxEG/KA4V5QD8jrXQjlly5v
/ZZi+3YBDGtP6pM96/DOIaweI85ZqZ/4TYMiIJkvAbGhLiyTk46cTUURsQYcf0YnQIvmDly6EXw8
hR6T205YuzzQuTA3AKeFzGteJnZRQXO/vUUaUeQD+2xxjCc9zSMnZ04nqYi/FU+INSnwqPaDUzfG
aI+G6zFNMAlfx4y7uIYKRz6hegHXFHJ7lekmhq/CwSCKYD2312KiljwL02hVcwsBT9RKhdYlK+tz
D1afnJvGgco8p4NjWEuTGT9aRDBmz/4zEK0PW/FI2+N8GlfV+M90pVvwi9cGcFeFpuoEOMU333gX
pU43Joj7izNYbgYB6ilWv/TggACcKYM213rBKIx11MnF9rg0fCrHHf4BKVuqq2v75rWdLP1z70/l
M91vE+AzwhS/WbLDLkg3dCNqx36s7HCJDnBJAFI3ZQVw3rkWptgs+2aTVIHc+u7Gug8UMzjb70VU
1oNWWG/mCxbMKA+f9D3OjbEnbpgHc2vZszwMEGCET7QeKoymLATCwxB2X9wpMSlWv7kIzJz2cy+f
AdiQMd4/IFKmjuo2/qd4qiusFptNzMDt6fBej1UhtybFj62VJNeQW1HpHfoYRE5GodYGIxECSw+k
7AGDypSVVMn/pHQ0Z2/rhww51o38US4oEZ92fTcrHqkcMWo4/zhmYEF1aRf1MiF6xrBbweE/tYD2
YmW0kyyv3KqKNKuFWKyR3cCx18iuvLVze4zDXMGVo3eFj2d+UPoU2P5u9J65cUHSGD3R66BGrnpg
8nDY1m+zm5zYiHCGtgM6cHrcyTIAeA0IfFilCZD93rGbZSyrhplDbrJPsHTSNmlKVJV1kqs8WtD3
8MAtxNJzbrbEIBUQ3gsX6zrCRlXRxjUDCU2rfUbdYGiXfd4UwY8iJJ/qSptXAbR1BYnXm7noYEH0
h6/a/pZOUMXVog8eJKj1Q8PZuc5bdFNp7K8PKXdvFXn8WsZuoUkcLCvVtmhFqCXofSDDciAgRUFQ
g26ulsx/UGGGjyzwGPQ+SV0t9Su1O9SqqYef37hkdgd5So8zAWSHpH5soaWbwRHnP0yeaUU8Lr82
LBrOQO/IVNjCT8jscOhmblvFWt/rgoiBxnBJ7vB0WvmaHlufpOgztMep/UzaD2BtAeFCNCmnjWjA
sPIOhSRRCMeC3kS0sJRusw+CNsOI4h5ezUrUYOE4zyE7uuv9kcWiqWmJa/NA8y19f7a66bPq/RtB
FSYfrYjZb8LgnNOgn93qAx/aY9XQolGQCpJodcP61OK06id2lePytHxiPXyh1uABoa/RgAqSm6EI
PeVv2YLsk+1nkNLwpEeYi0gUYqz+/Dafm8KPsrKyavbiAxGDwnAjHay2cH8p3WenVo2zamvmXK4C
0qLdD/tbe/PJnyWs+WWW6na0YscAqEP6H3+P5CTtSO4wt5qkjSGmf1s8okaKmea4+uTntQSkoQLq
HIsQ1KNXpr9RKePTK3r8m/6DuQ2xsR16U314ek1zbWLdPkK2HiJylyoT3cmKDSKX6EjwB0ynl1L3
BFubEY7/T/qSh8MsPpi+SwSH2W8aWh7vz0F4kL7+Kk5g2SgHe06mmQFZ4LnwdoF0PExPmsRlyfYt
GgZC/QVJyOQwCSCcvEvyrY9X3+yA55CdVp2/xBlXocjuNbnGmd3I6L4CMb5kXfNckv9HzAL3OQKu
DSsTfBsmuvnQs99QbdfXF5KaOv+XWM4GZjmYj2o01dcnOyN4aTXi2P4bVef/QriQXZR/KPFs90Y0
gXxHcfpo3HFF13KzqZDVXnw9dee3SKtgyXS1iRO0H1x6dp87fNEpw66ischEXiOcpmzW6b9UPXLd
NFZHBpyFtRbPCD5ZXclW4LlD0ycuyPnnH41Gw+/7qtUIZiEqN8IHy8Aj7ZAIpnp+BgSFX8un9fal
MpKiLo05toyv4lRAW6ovN4JfJqbG8fTTOHxczDMiKA+Ibtp2vziaF4sRUx8rt+qCMTbryhQhjxsO
lxxe7Rj4QJArzwIdY2IMRB2z7UOQPcesoSGi9ARUrZLc7VESBV0Vyx+upPhUMPdjzh3dQGhf/FFy
rl7G/VXISjxgDr34U6y0mm9R/EBG0OLqaH7ryIZHurgBkGL+sFaXVF2/JmZ81G3T5K66zlyzSkLY
iYubKd7v3BV9kxpRrgqtg6BycvJ61CfCPZk3G0F01AOzD/qK2xUgTdqi/IOhmiqHiIsEEZxHYrqI
QzES0bLGCuMht5brgf4pvat+kXVjzggn6WDp1Ld+t9LgyIZbu+tboOOuG8XECDL3npEYeoAIOv6e
Yb2Wu+lFNcBB+nsi1u23/i3VfIPS7FyVOmspQHgdzxQgnQoK+Yjy1V5ocRL1fKMrglJq+1PvmtEw
1J3DbgJ1oMx2JTDiUOBKBot4QCVQBbZjSD/VYuTOKyA2/8VF4cCw0Xqns79lzVw2isIW6I1o7oBL
YMflsnU+ge9aZ0y9Vf7bYgBuWqpyCaMUYily0E8q0uoXhSgCXhzBRodjJY1ndp9WvpSrk+VPF3Uk
T3Pys3bws9aOTD9jWKkJFT1etk1LrNX/OkY43Y8yYihtKMc6UA1OTLtc7VqwH5dNWZHCBVkC5HP7
x8tX/iggailXJC80Onep21+I6cIuSvRX9/YRdYy1RtDfDM+kh2UIDTfvPHiZU+NUMfNLPN8K5QRv
aT+S0rmSLtzdgF2xZEQAcOpX6JmKGGYS0dX1Tjzkqp9CKtR9gAA12jGzhHEne5HuWUqzOmU7AI65
DoL2unKAQboIDe99wj/DANad63XPaJgKlHmrlY3CX1or6as51fDRfXiTYc+l1WpRSbUgTrG42vJ8
KshxGOXZ5Gu21twUzFoZQiD6p939yjYjQKWEjsBo56nM1qrBh+GwoXqm3gh9Zd9+Bz77IdFyZQ/Y
THSrLabidCjTzT5CUh5iqqUpIxREqacRgJOv4yS+PMduVZGskiGVv624Hln890T9Y4Y7hb3SENvp
OsUx0om4o4E5p+xGacG2Ju62zKsY/H72KoON/B45ftThMRg49UX4aQDVOH1aP3meg4PYlx9pxN42
iPzeQdxi3ZtDd9L5ZxrfTA8Yfk9yK3ivNXX738LiTKhPckd5vmROl5muhRnpgrpe+eih0oSdHPJi
wEB1l7uy22jtzRAObrg85cd+b+sFp0olobcuRK3NdTgDJB9SiNiRjYRi3oB/KUC9qg27umdmr5de
H28daqH6m3fQ8vUVl7g/AEfIBZQ73RNe9x0XwQ7BOzYAPH7vuPh7CdW5p44Goj3yPZaEJalaoxNS
c8gDcRomU+ovTfbUOioCXTQB5t+oyHMWurjXRFEpIK0dpymNCAw4kH+adJ2EBD0CodoXJqhZFTaa
oqLQq3OD/Q9DeWcT4fTVEfwDkygOoQtyxMHyW76kfthqXDdl+3aumTXy+A1BGSZ7Iibquk+8Cin0
AengLiK11IFCqQ5QKJhChG64WEmSdRSQ+SMjqpwtGE5t9qkPNKaF5oEgVwN5xFgloLy+Bv7h5GEf
m7dOJpv1v+7Kx7KJQFy7/ZLhHnfKOspLn5pPHFWyxh/al2ymr3uot1BM+zWVZbeWSVxskwPaBt2n
zmgaw2DR2V7wcF9Kv/92pIjSDGua1X+G5JLIpo6lZEek4wColSIB3mGoBzgBm7O0BohMVHZsdt8N
zrDaAV1z2DDZqZlaTYLnRtO0bzepZAqNOJtBeeaEoz0Gt2efhmPPJABgDVI2ApqlbLu0cNmwK//T
D37EhY88wzSzdrzsC6KVzdhnAdgYikc4bFxUsHCaeS+En0/x2LNfUIUsDFNcc/ZuC9NmjxHMH/yS
eZND5WyRrnXQTgYYGtLVrB7g5vH6MwzIRcLIANwyoWW7YJ2jGSNhdCLtVKKZaRqGBQx37hwtF6KS
hi60bWRMdw6UbNWYGFhrKG8pWMZoI7ol+VmzscSShJbT9ELHsmQIx1KPfbiCLYgWZCYMk+p1UoM7
yhrcewVI1wODrEbxNbWRHHYg4mw/N6RhrL/KXNgwejulAXnnVyEv7xxiLNkHi2oYFd57uLQIBcFI
VrLJ8flktTP7tnN/I6O5rO52TwzFie4IEnLo4pchpnlBeSy/IWugxyv6zyfb61s3BKQknKAqjF8h
aOFpIaVzogsNBzpjiYzEfCYJENAE4Eo+i7nO6mLC/jOmCK0vVKPbpkbsM+QxevZypqGj+68m3K9h
hd/guQHEfyudzQ9uipPHFsNGsEDMPS8VbgTgndlkv+5/MWrcjpdedEszOuG6DtPwGNI/YiI+UlUD
FTH302+nhhTAM9zIJT+rjKXP0QywZcpD7Fqe7+gs8uRzfib4LDQNhDBoZ458n/X+4LskazdvpKZk
/0Qkonh0fpKJBferKwvcAH+/sif9HDe9YtP9rHeJqAEm+E6SgdDhLVSLIutQsRkAswjla2i0W7ov
zwE3ShHB/9ihHG/xxRcfHrEHySR8AQb/o5/7/DTQIhuufH0tnYF9JDjD/7fHStSj2q0RaMs+CsLh
+uxFOQvGaX7IfdDE9SSQHOR6aPrLT9tDS70ALxU45mjBu3fUxfY4xaMt/Tu7/o3UhTjAGwyvSvCH
ZfjPv5g4D2VDStInydZYqLhbK2j4EVuV25MPTS2PPVzd2ZxvTU6GKg4ogfzzNQP1hTvYrAubQuzu
Zr+P8Z2oW6p20lwWqYUjzKvzff/I2pd56C/gX3yx/ulNdABO9eNHUEE1K45gIjtL9cfjpq/0vlyg
4XPuzH+5kKiOPrjf/teVVDsAvRbC2gXTjUiuwEsf3RZ2/kIKpnZodBe3xIH3oQHU0HlYc5dXWHCy
VJB8nNizLfxgr/Pzu708TqHosA3lofln3BD9JcXj55us9nW3l6TAKbif3PxgbBJOupwTkdiR6NxG
5fvTJ8LHl8fuX4anntP20SIlJb/wXz9ztkQ08I0P8duJd59xoYjv4f2u8Yix9T+tnipgHVoizwvq
u6VGwELbzRwKM6VFFa66/SEShvy7uPwCCJToRR/Rpg3xoj4Z6R5iKvGwd0R2X7kqTtrSX5+8a/iL
WFOdFb8/b6Oz1/uoc8YDaS+XqsZDRNG0bETt9pKUBTmy59TIVKtHTGAfBg0n2e4FBfEeRnUm5ahZ
iMiEMZ6N1ESMyojXzR+O+T/DReMYJsej0s49dk5tUybVM496B2ePJsQjsLO7NgZxqydBoj+497Ip
nj8+BYwTNBInYe2a/4DlE0prmdfzQp5K9p9WIdpWwFfd+vyQcLMUa7kbI1NDodFi69awdG8k58t7
6EjclsSMq5OD/HTiVPK+Fl+KIc+oUPRUHi2Z2QFquyQBOolKMJf2ndrNXD5kP3y/4a0TgS6x4DO8
rCKSwZC7pm1BoA69oid+NZBCJ1qCkhFQUW/1jukJL3X0E14yeQ5TcFtI4UWyHHF0qVIiCtEzIH1i
AKERhDmeu9NJ422gedZ7tQ0A1PffwFziYReG+JxRv1pzu5D8HqG/OAGwtXAvx0QuE/6fLV3w+uTV
/Oerussjlmb4G8PzeQs62mCm+TjXwvMyIIHk/XlEbxd8gh6X4Xl5hLNEjWCtyTnAZZksOVsoGcF5
qpTCJe/LttJUA8RvOiv/A0DCDdEo3uQ6Q0Akg1VZyLNLpuPBK1VnMA0VU0sXjX7gGG0dVqMTXn6p
7Zf4y9jexvVccEhhd1VYWfdVFIXuACNUj0jp2Tq2n1JzVDbTqTtEmqCe9kWwSDM1202sTVdW9tQV
A8yksLHnYDnIbCShfuuvTT3QgzVEbai1mo2/Ju/K9lJ4O0qFIALqEhevIJYoc2GKR8hWsoM/pA2v
xb/wTQoQF5LgCWlauQzY1FrG4Zj+thOYoAzOKSSjIOMrgtq8ItOaM+8c1xCTHMeXQwLuprLiBHaD
r4WS259cqVGennkbFMVITj+rJKNizZluHA7BYAiNqebxvWxrm6qrboGl/3JpzQLMkebhLyjWxka1
hJ2392Y6opMTwX5aArGiJESHCTzq4uJfc5gseDA9iNDxbEnGxARBQvAKN41M+3EvCd9RT/MciovR
vSm6vxs/yw5JBnPM03U+FeIioC/u3j7TUXJf0UvVNC0uFFZS3YUYp6C4dMbuMJzN4Myh4I6EeFis
RP6pbvGCEjlqPSW+l8anJyVpSKy3jxcvs4VlRUiQ+8l0osVj6T7I7kcjhQrqM/XeBYi4oUKV0BF0
WP2RpfKM3jojP2fo0a1+Yc7LDBBLSrQzueoFaKbl31wbXe9H2W2MDZkLuErnqkjRiTn1G/thecqX
Jy4Ld2AuPNS6yNfTNVWvKqsxFpCOy5/7Tdzz6ISiMNcaIkK+ZDzpPgCY31RXOADVunbC/YnDh5vS
M7J2UVnxyKlR/J42NhyC/UG+p6+2QAnit+6VTs/RG4l0Mwlxi+ocXaFWTYzk8CDaunt+j25t4+BO
FTj0vXHCb8COPQ+X/2tswNqabYc5otUk+nxbX0ZvAn8oBpbRtIpHtxl5sEdGuJTnSu/mo+WibMLt
jAUhEApFL+adxt9InXmQK90tU4MvuvYpGbJVDjBdaFNU4NLTkT/HUbBFosDHAftjYgn/6qwH2tk9
cqdhvMavVl38dCNsHGQm1gSWBFOPeDvNP4Jx6HAqLOj8+HE98i8tr0vUkstwQ9Fzf7YjYviNhuEv
x1wYwhp8rbq+uY3BCVuRoe3jhvbNx0HyYty1Ksw2H00ddx5dwmruBzH9jmGyzOsZQvLpQ6QHF3Ye
rNFYbOYtdcNkMa8qa6Yx8uUedi7PtEdPDjlxra00iKezHYrA8jISqhvC6ZrgdwdH0c053IsZov0M
No42j6U4y2DxmrhiiCm1LAuCyrdl75bzGpP0B3zliz9zWxhR0IPWgJax3wCtBntevUPtsHeD0e8k
rTuWiVHnj2rqrzLNcwVwyAQJ6MtFvcoMSXOazXGOjOXKCgJ2mU8NKoZR3UeUOIaxRGaq5JeLO9nq
+YeON6zFfUxfv1tz9hooFF7oWDokJ34pu43b9G+UYYHiRpuXa/npOHAKOiuUK5xyAWyB0gztamam
9U9JXp6K36O5vSYHHurwAk0A8zNMWjoZDiMTu9XXD08coNGTpjRKocFOPEMPBhIgZIm16r6Sd7zS
9Sjy6W6DF41G+taSRC1wqM/DamXserJoOPFTyzTII0xXkGvz0btTo8r/0bGzsqC8KHx6zjq0XqT2
TJJvgXbiJdlto4mIy/nirhqL6+ANjfVPkuBwDxhQ0TrQB16RB7/MLtPyockZzoETAHRE7R9LV/P7
D8XTI1YVcZ9wCU7fIY5bhCGPse+4YnnlFtCSiRj8MZJrLO91W6iT6kK4TQkQYdC+fwFV/3N76o8R
PVLK1ELA7Sud+L9IiahNhgEYExQ8PkBOcgzkNpvs0MWBDrGKRN3bRoq5YQEyYp6Xx9i7QgWyd0Jb
OKiUEB/EsE54Ou+21/ppGbuTPJCKxhRfG68Mi3urneERajIBMSU/yF7EvYMlIloH3uxEvumIWy6n
+mD+3WvLhIPle6qkUl4aAoMfBZSsRA2Wx1ZQ0XEuXymYylrc8OqVSuZwDPVgT62dN7DmjrCJOizT
Rd3B1foVwzjnm3wyFGTQX7IKtdf+2PI4xYMTDZf2MBqj9b/Wf3qcoubdJNh9qmmAafQoCWM/2png
HP0OApdTg1+V5tS3adFz2jFN/W17wL3JIKY/3omAwFvtp3QRcBA/Tjs9FKU+RpB19DxwjMD0B3Rl
BTq4JgYNIY6Cz32i4mJdN0Km7+I0JgCdg0ZeWuzY9LqVVfQMca3qnK32a5s/d/jqrRU8236IgAa8
TQw0fHa3HOPNvpg5dlflhdPBa8zy1jL9XIqah3XOOiXQ0e0AO71p5o9g6Zu2zTI0ct6P99UrBZFb
1AeAZDcAN/lpaHtT8x7fE1DPhmsS7edeqwDMclmxNvs/5yuJXVpmcgYr8iwIcD6dDGtQrjocotWT
px+xLj47mcXBQuEZ3OF0InSHsK2ds1L9XdPVfSVgBM28/UkVS3zHz1511D6v+NgCH5uQrP3uWLoX
Os2dSC35Q3KdAZFBDeMgagU6NRk9eITPHmJou8hgW16pHXodwTvAK5LS1fkJLpzsk4oTpjiTjAQh
a1TJ0vNM2FoxQmxP/NuQ3y1Rba6oTXq29IM/YmrlsvUJrIpD77q3hO2tR5/0cLzor5lwLtD1ks5P
aOSkRzbaOqQCCkVYvTNYKb5aTHUtEd4j0VyLEpxlnsZf8DZBhZG0YyKieNXKQWsUXL8IrGxmdaUE
Hpny2ehLBveYTLmIghjUYpchtqm+QdEmmKUC20oLOyqm//GTX0/5H92hT2uyD/bd7MAaLpG2Jtoa
3Vjd6Dwjgz+PKn9xd0wkXar9BBmiH1gL+qIeqTKFhRBtCkKMtcDw4L8DlQdN69PYKjhH/aRwOSjZ
eskC5KTIqlCyY3ss7LYAUqrqAs7hlPgKufbOJPiIYuLfYk6JmCNW/vMpzI15yNbURbRvQooHtxnQ
lSsSL+cJvhyLKro3xrcZMSDMFqAxhmS9OMg40eYDkFaPWu5fsvixPGHNmakAuw7zpmw+DK1eIgCK
UtgXFdrfyT850oBsJnIbY3D6Hz3KY8mMgT/M3wxONfS6V7hMxgJYo1lzmn5P2LwXhSEEE9C+RFBq
nZXetIVcIisFOQY5zfSUmXZhdoStIqjmLyNcSm76gJ4emf0ttWm2EOHuQBND4D16IGjdMVlpfS4a
jIhVeqlnvkxN6/09ldV2MQVfbCyiIaq5a4+sYCaVcLlrh2Bq2agx3ZdlLkLJox8t4ZbSwwV0WGmd
JgrdS440FXaKbK2Nw3y7nzzYCYVRyMzYR8rrtWByEF+N90eaHzsEQkYtfKirSCuVtKuzPER0O4Dh
FiWNTTvBMw0gaK6lDyoXDh7IOs5ZDftzrz+iFBevmsMiTHXzcqKzhoFdxnjj3D55zVZi5j4icxXR
5S7XWVxoLwv8WNsasNATMd9frVV5EK9Wcwqbgrl1Stca5jCVqq2Pk//0sZ+kDAPmXQmeWC+kByI6
CPOAQY2OTjJY37ohon7F6Wr8Una7dMStNFAKQtBIz3ft2ZslgXdmNoY4SeGix+F9mBAHFhbkxmNy
RRwDkgSRVlBwMH8O4k3E/i4rbJW86ykhH5D4CtjXWW0WUQX6XrPZbfbOMRNGfNMHubJLioAsa8Rh
LV7gAZyjRgermYJWJikJNirdT4pf9FyeZ2BAwLUv83GC0VEXxhIMeC2UVUQOTB/IdNqQ3gZZnnuL
Rh4z4oAuQ73+CxGHLj75bLcPiTIdkpfxICCewgLcouce5oHdBHO6vIw/n0cjWvDLrhfQV0TyvdKL
MpHHwWoUKThII+bfxS2MUAlieIkWi8rdwcKHlYtTCKEaw+Cc3l6JcpjrFCeNElx52AJASACHXy2P
j7kwRtQ/JmVelV5lJojDlJ+udb2BD/ceUnmphOq8hIx2q56obcUPVCvTGdgfF2X9BApq2VXUp58/
MDmbPYML01o1b0VUGYDxqNGrtiYGFe5MiH22tIawCkcMMxTj0z7zP3kSRwLuWGBvu14SoGNUXqVu
Gtf5LJt89ADDvlSZf12QTjuiBF96HdYIyCVpZVLZbNKLYUQpJvzG6I7gmBRaR5cVyVvJvAU0Um+T
DVufadTdMFbc43kTWWy0C+8aPFGq2pa9cq/l4QSzrpnasQQ3NZ9F/c2X7Bs9fY9WSad4H3xJMNSc
EAEBwT2j2XTEtVJaesPnMJUdxpghiPAQP/PZLfJdZOFXsiU77igt2GUU6S0e+xVejevo0g7I4QcE
BO0M8I2qyw9uXV0cLSjJDLrTbYCkT67BGTYlIKFPRt92YHKbpGKg/xGafPv759ZqWEH3iWTvRAB/
tpDqcIECOkcjQ20CGNscITuHMo1zRtlr1MyelB60r6XlQ1nrToNyqlh/ZLccMhRfVZn9Mcqi62hg
SOfjqdEpt3+LQv7LMQrfbKbgAl1KXpVmdryxVddXRJ7WbZDQLRegbu8mwayPDI2w0nAtDca4JeDG
bJvflbWINWl8ZA8zn112UezdAL6bwNLPMNx7bGUy1zRBMvbOh2brleWGS+U3wrO5N11rm2pL7LUg
pdkhPK0/GWWCd5qCMMoINr4i+XVA5vBLY7r4umgnGTu+deyki0grfYkYhv+KZj4SEccS1pKdvyRZ
sXsOW1owYk5Plwhwr1TP5Az91OSlQLFwmOvCF6ApPRHY7mvv4CRUpYEafkHjvVsahqJ5Y37uvP0K
Xhydb+TFUZquUGBh1voeyqkkseTkuE7F6bFonuxnznQECoHowh2h1NG6QXs+/kjMwPHep5RFDqYy
hJCw2r9gNbGd6M0uiAceG5SLoIlEpNE/5dKp0ZhiuVEeaXn0eGrroZUpxpjdMaY6GKYUOqomqwkC
GSQrXG4+APihpjxVrqP9GogVE6Ts7vmG+GyJVyIV/na79E7341NIRNug/3iXTg1jLxW2BgOpWvNN
eYkXw21NLlmdcjgPljh0gAZcwpv4+6Xvh3KtIcl6fsMRJd7sZWnop+ziyTOKYdR9Pcg+z5SUc/5J
ZKESSWsVeP2vLrVrmv8yJmzGC7BQ+wGWiV71MSBmshvXo5ItuPp1hpgH4OJcyVWSJPD5IwLa6BiU
ndN/kz2+vfcuE/7jx+o3e6qhY8dEBfisp6QLd/EknYuAt4McV7HU5chyS6X6Y1aKVsfCu7ZKMK8D
bvU6FSyR81GO5giteGkyLhwKWr4yMCi+/tZ7HHbGXjYTAP+Wn4Mg4QmR29+FDaPP4Dyfh+yPScy1
HlDH3duinXDzHidXtNcRYwyARCiea4ckNEFYL9caHA+OSYClDbPT/yV+4U9AQA89ur9vd6FuIJ1s
TfFpTLaHxDDy9h++rwXfljBIfctowQl41kkVHR5dJ16wHGyAWWkQ/DGdyamzPzm/sksiYCe2b8wk
Nfx1wtcP6ypTYjID7/Os7qL27/B8i/ca5Xp7bxrnFUMj53I4esYYmEZ6Nru36NnO7fb4OXA4j41V
LloRZISK8Q8PZwCnhLNCNQXXVfig13sQgLohyqekq83vVfxSC2foV7jtxHLlgR+2S4ZhNJteBtm9
XpUGNMHb6BSgQ1FInOPVo/mJokSpe0MeSpYYYjb8KY0/lhZh9stWljUNGI/cQfpvVq0FxSfyjkKD
fwDQy1a8bIW2Qtd8VqobMhPrUSSahFcV2VE4BnB1Vm0ArxJkazzUd+jo6kzOCTwKy+u86K5bh9xT
+b55DIcbANCnz9spR4evMaohsCTihRLl9L5MH0FzryU/DmJntyxIvs3zpIN5vjLgbwew0F2Mzhep
M8YAqttoWzEjm19DR4eYb6TzebBFRSsc615Icq/BEZ2evODlpYRzAIyqsa41Yq7tzjNHMoHwrqUv
vAPT9io4zFCUR88C85th8oelOwQGGvJr5cRlMjhoFA1Vv1LwkPoX0EqSBb3p+xcv2U8MRyWs75HK
TwQxD27vGZ7XqcYiVqpl5ufhwEw5w//shDVwZWoeB1yC1Y86Z96j6XR8+bVrgeYeOUESJAReW3Y4
Yi/QIhZkVJyVpKP2A6u9hqp1mrUr0VrUpTGLzzhiiuEy5TQqEntWiiAH3szFS8DqwI6OBiwioKim
cCvBZ23LGYm0BTsTzsksT9wZ1LEHodSu0Pq5HAq0/uV0jsnFK8S3stqz+yGKgQtcuTFAFL68V7Vv
0mfuVcQI2CZOadKmZZ8BdZXgWD8S3U9B+i4xKibsTS/fMHgtDEMeYGSceiEGnoBXpH2QFycyjUdD
TS+iiX4dZi7/r6xMcDtXREv5x82wOM4cMND5Pt+OHDBJN9twYRsqo2ldmf3CdLgbpaRqUBUKd3X2
z2eB9QsNNkWgeUUTdNEUDfc1eGasmyXnniYbzidM6zkgqOVB2kM6n2TAGfabuAFQaOZI6NFn3v2c
Ffm8AOAbRpQjIPqL65Ir3g14z8a6x/b8J7fYySIe8WtZw6Yir1+J0P+PPV+LUJbLpOjOlmvdnC8g
eoU/E4mL4+al4DGIAjLp+XKV0I46+cDoqRYk5TQsOUCQhYeSpwfoGhT9AB0YHOi2GIg94lcbssok
n3cDq0jydFMT3/dW3q/dDSjv4WuWhVCv+od4YmGhaoAujVaYVYfPZ9UzWMno6RH5GM3LGaAj2sSb
KbEMmnpEk0Fso1QKs80i1acDlGKbeVjcSpIalGTT3PkWeZ6W8C1X7ic+NCbVm1fCN6z28x44nFOI
9yZeKjGhMHDm0XFsPHu9nR/3C7iNRh9jK1712Q9m1mu/AadE22ymY0/pzx6l3kvjkbqD1xBbJAXH
iArH4eP1sHlRibWsmKtWqvuCNBB+xLNE+J+8C2UAJhttJsi1Gappop1QuhzH+A7GQUQfq0w9gkWX
MtGqhemU2a9nYq54LNWzhi+UjRTf7addaG4q7dtSuLdMoxCCYaW5CvwYn+CIO7strfipBmGwTX9c
vRYisunbR5leWPM0qKT17Pk0oCcqIKAEHVZfuJCwqABm2proJk++96ID+Emu2t0sSH7IWfgHeT8q
fVWa+N25KnNrNcx4yjulK8kTZvIPAJABO4s18zdzwjPEEbnaSt98ZT7OLU2NdQL5LGvAv8iRrB8B
yiQv6hrcnNql+OaRCoPwHKPvNvlzGpKu/GOD3Zq17GMUlcZWHgpZyPIYY/lJ3Bwss9/FxHY+llNM
dtOGJOwpVW7LaFa0VN8oKaJJiRLHeK6WdiqEaBBIwg9J39H0cSSQ10ZKfBRmSdTUDBhEMjVU3qbu
Rz2BGckJgNH1+syoJ9LF2xcn2BRoY+dkpuPU0odgS0b+MUQf0EWY+PP0WGPgMO0yEohRzdhEnz8R
s/oYSQ2u5i5TdGCwMdqv+c9IbjyOD4P7lfJuapEY3phl+cnQFdk/RS8etLkmTXPIUhhyNnA94Ju3
ic6EBJjirM2CmKniEp5sPMnO9eIkQgFNStH7IAw9Tths8tyGJYwiVSTUQXk+pyXT86pwqEpzCPPB
xq2Tj/EqEcMj1XO5OCmP6cZdn2haD/aS4/gwFCRDN1D0T6JOIxW82Kq+5MsV4DTf4U4V6EoE6r+j
ADZekl2XDFKzSyroKH/uYklr490wiSSYwQlzeysZUWedFB7sh6nNiWE1+m8d4orVqeyx12J4DBs5
mF47WtA3UifxcwEsyOfU1DeJTzndiEVpW1xTcwWa8vjEY5xDfiri0mb5lsYsXpVVnY9Fzmj5mP1/
+r8bkyRxyfYxgaLDi1YDKu0oF3+ou8FhVwzl4n7jIJNOJfrdIJ0fStwaGtHRSLt9W+ob5ssEpG0L
Fo+Qx5/cMpSqYL6ohJ40i2DjXAiPwmsQL1a/gpKXehPpXjKD2DYO3oCVpU16TEm97ghRyXUF1u1+
Cscp6uappqRZKRk7qzqzmsGShVWN/d8Op2b4l1Q3r7zXZ5ssW38S4ANj/pN1FTtbOAzstqVWQmV3
vJeqcDoiLcVixda9KE9+c2m5F46e1fmezMiLRJHdPm0I6+VurmPTx2mZW2o/em1o3rhq43BEuR8i
vbI9TGMgnko1Qw7VbR7FCOnwoChOQSgq2PaI/z5q3C8ciQtSl999/dWTd7Tn3iXQ4r05lM1ULmpD
zejfQuLXt+rn9B8huDDb4Cv3K1AHLGvPL0jGOKjwYaraDagSApie8Ha7fU3HjN6G8uSb/dGEnxDj
/pzrw2aMiFn9GKcfKiW0aBOWsX/gGgLqZhEN0+qcPSZUTcKt83A+GQZnPGqKn7kX3q4bBAWyZxcn
I13sQPgU7vctP+PWk5YysaFFWJlJ8RzQRV5I5sjhhD6WdDYhXLDf0WmvaWn/jL5Ova0dc44ggrS5
XUeFJD0q9b49YchJSdCuZywsY5j5saS7RKZaDhKb0QvG12Qh9DSCqeMraxDhcSYJhwUo00h05Ria
uP5en7Lo6CjyZL0fCTn8fDAC9kD3cPOp0oNFDUoXMAsbkVsdM8wOvgMxfZKjPyflCWm+XMtBLI+B
ci3iAnGQRXgpjpPrl7dHey7LjZ7lsqEW6AVW9x1r522QP6T8RbTM4lcvk6fAbl3X5S41hmdBua8D
5LCB2JOl3BrLBLy3ZAdzDLkzmL/44aLAH5YCCHsq9OAdkoWBjZdN+m9k9ffyVIREOxQtKy2scDsH
jv/eTEoaneoldJklX+o+speBlyCC43TRdG5f+xEy6AMF4Khq5ZgI3mdwQFzU6HMAUiSoUvCLCYtC
dD3hSpMF5278q+NJkAhgAh7RBaFRacwEbxj1pRbbHRUS/ZN3UZzT51gIjUvLb0EfxmQA9HNjmG6h
z1ak+DgsxJ5t4ttl9objbOvzhQUd7AMZ51WIuUSXMKOphD7vs/uNWqm5QGNts5l4940KAv0TXgyt
iWIaP6VVnUSMZE1fs30GGux3J7m7L9g0661aLapI0biR53VV9V6dg66uP42l1ve5iOQpmBpHIU5x
q2n4YxlKjjwlX7gUDbV003LID/6YbphEA2WiSyNzWHKzGWDTlwpZJBaSe3dkc6M/rTRCktManQFj
eP/mbTpcFbHwG+exIq5fzNd3zkgSUN7wlcoEP4VNf5Dz2dGH1NUMkQNcn6MwIHRFglN1xGt6E4hF
dwnxk4+pcvXTGht/YQeIyobOPmA4JGfk0z0dmL6weU6WIkCx6KvgHckOxS5at5TxSU9Mdp5znN8V
E1awMcNlIWZUUj2v0gFJEc5FqgY1PjGvldFp5+iKAhYS/nwnHG2pMYoieVHpGgRE5TqZ0t1voRY4
Ec9hE94FAa05Nl/FY73I8lNNeyX1wab/VqTuuiZ78YtpukD5x7lldlNSHzXNSU7dtkDHVEH5P/Ol
NqpUWP+G/JSHhEDhsO1QUrDpnGcshr8NwSAso3LE0v7kGEvXW6tn9QswYXsjMwi2DRjIrJoisiHI
Ipux659NQmlMPulT+V7EKiBPjK4dr+rACgTCSZcbKiu16sa8b4pU/OtWs4dxreU34CAJzmZuxiSP
atvL8tqFXT0rfsF8vCR8jp4y41G5tK9Hm3XMKzFrbdEThgQVVx31cT+c7UlJb1ml7qChAZf+fRjV
Q870EXRlGGCLtxReY/KW+aOQDoSGM1MU9kXvlCeIlg6hBlYTJh4ABrKPF5R911aI3+JQylDDVhur
ALqaYzfWpiqHpUI6EJwXzzRKCb3XMT6j2CVcISS+3efjml9zJtU8/5aBavJl3ZF0fwGFjB9gp8jL
LOMgiXfYjcdLfyYaqjHX/1YoDhfhOVWjvw10Jzgrt82svwNTUWnOpHWXTAja9XYhPFSvD3gvZM/Q
S77KG+wxv/R+gWEVeJCIxZvmCmMi+fxOkpuIVgOCPHzejwUYfEBYB1AMlVvvAjtEIabrNQEJHu7u
GlI4krcDrJ393FOw/N0y13w+6byKqEIxCdEGHiVe8oEUL4ZEU9TI//GV0kZiBuTLLO81mT+GR+3Q
lHc+aA32zBfYmtK+Cm3TnUjt0Tzm+Z4glUkTR1LYEUMhpdd5R+5WvHvRF+tZfuVfEipSYSRRuQvs
D1w54YoFTyJL5Z4rwDdcLgmzchLWbzEYFzsskGFpWkg7Julj7xJCKF3odrdXnV7JdTyCQdmPprvp
ofktYJ75vqwDghLBTOhSdZbdM/ylE52BBvMwussVMkqENhMxI3faGY/q/Z3pD6f6K94G/bNC+8gi
P7fANpX8S21WQOba/9Zb1/DdbiEGgN953SRJ0IKX83vsI+z7JK0aF/f+su9JXh1HZD3JANEvz0A3
v1whk/MPomCAf4QiJtGqzcgOIUqenz/hw29/3x/9BTDiAJo6/A6FjNa2mcOHXxY+3sXqDoDNFaUm
AExV1eZNiBRV+yIGOI3jd85K949Os78TqgeC1lD5T08fhGFbqx9t9wp+H98RXKd+Mx6o0zciacli
D/N+tznMVaRIpwGu7iQFZc4LAnq3VBgG55APCDLKgoAhtyBaUde8WF+UsHpZxR4rl6jrkpaBbqEg
X36QTx2u9fcDu37+oniF2HWylDXx8XmxPkfb/fNN7snXdb0akom+RGJgq9pDsBgGVlsQXmH/NxDc
h2F3qui3zTEVQVUlRA5lTGA/6kssCyR7k/AmMXFNWpvCb1pcQIy8XWiBhDVjg1x8l0Y+QKX6rc5f
j17JHnTGy7Pp1nqwcdlNbm1wFQkqu2A7/rFQ7v3a+1jlYMhj3fkIdzUenvTeBhtGwFzwY8DQ2MOu
XONll+6ZIApstgCGAuJ1C4VTMFH34I8g2QZBCGuwijENyNxlPsyU6t9O3onuHxry9nu/hMPYr6JC
WGs7GfnX6O2XXLvVwwBjE9Rhx8KSsvP925rybY01RETWy1tM4C+fksgFtrdSu0qT13W+j9oqgxmP
0fkO4rIjjOgVc6Dt8Qn8nC0l1XF/bDU2p0FmwAMA8YJiFZPTxoVP31Yw2GGuArJml4Nio23PZWsW
6rjtGYLeyfaIecUdc998N5/9QyfBKAff/f+MhNfQlue9GuMozkG5g6tuvQBUoW9vj42ogXO/wdL3
Z69zUcWVxt4SnrGzo7Qun5JNsz1uHyFrWDe6zUX4VaxB1GEMixfWz1a7ccfkL+G4I4TWA/7Y0sPs
e/JV3YOtkxeWUApJ+hKD3JdP30WSi0DFWk9eKg4nTZeq3eUg6hRDCUILlr+9RaFpC/JfcmLTkfKQ
OJ58LKbC/O5EG8D/kpGSV+KBo6h4Y1LSWA4XuDNgB2JkqcEjQZxfAfPEJHmi32CUoEHGjZTILeDj
lNo2KlriqnG9fqyLPY8EQ+mWfF3vzBE0VdV08LBPX3kzrmjrN1W8aNZlfgKtV31Jid/5/0InrShe
I3oBujDaLXqOsXEPgLwrsHxdhmuZID5tivhMfm/Dn0fhuJNedUxMG+ib9w7BLqvgOykcdmpkX6vR
PILgK68gooGZHx9g5AUd4cqyWwrVlaZlHLvN1uALb0lzBP36z7asD2L5hwMv3gQ5MRExvZD9ynmR
q1DPR1fGJqv1TF4cmJHytMMjIsfutX4oAyV+4amRr1v5GexM/4zkVgIue+MaHd906dCSa7lLAUDD
Rz8+ETSDRTYmrSAZ7GT7Lawg9bZIsY25julSzAD34mV2DT6/IEFEQIbpXgR2C85BTSQA+TjHKRzL
m1lxQXjLhLRaVOLU2/3lqkxULnNkaEKM4yYMSz6UmaZlq1d7bzndiOiyJyW/HI9fb5SjDA07GmTv
3X1b76PhQ9FNeaicNT0+gYaf+drOhKRYTHewubpUEfR0VqilC5hw+F1ePmwKP80Dh0TVHs8eipjg
HAEUuukkMP7E7pUS3rPyDWvqRV8koBdh95LHqNcawrm4wdc6H5thDIvSugqK0FPTnO2cwk0grb6z
KldvAaTrgj6mMe0K3stkHcxf4HIoVU2OoCwl91JDhJxFfwb91ddT41yRX6vGllpOGyR9nceG2W68
XgT/QeY3TqvjCCtPkhuhfij/coQ+ehxp/IXkkLsh7yFa1rWcKZfz2dVHxT0RkAT5+OwRAoUSSB7T
p3JFw9TYL7vq8bYCQSQxPJHQh2wKge8t8bw9sDAKr7iP0ClsvRFpioue6SYbEdjg4DWeIsPzLaMY
N/Tlj/RCgvXTIMHUx3HT4YPYURLMOzDx7GXt5QnT0hjlB7puiVVvJREhptIjt37iz/pUIjLxhlXU
0lgTuvE5QQ1X04FCocncmGPeYw0rp3y+VNh3AZtwaP7AtHJTBoydhwjyMWpNeZS5bjDdmsWiEjF8
+pay+oe/g+Q6336HNiuIEZJsCCzWxPowM+bPreR2wJR54FjElpFNSkjOGgeU5ObJ1KDLTGE/rDLT
7oHDCSUDx8SA6DtrQ0EQ+mdkZ5CNP7O9s8uccRsnJX0Opum3vDTAQ7gCgVcjOB9EuWRe5e0GBS6A
eA1N2fG1Jo6OGjAGPpWlcse2Rk1M9Ok9AUDGXc3+zBNS2i1ogB6LguTruZSShVFA8hiq87KO/GCT
8PDgQhLPJJclUYs7b7cCVm9IT3umzC4UvGdYeSlUa8Fv6EGM/ZmJKg9MPCvFlVlL9zm07hO1llyb
HxoLPpqrfaaih5kBzNVtiOr1vT/B2ao9eTO8NaJZxwFw7EiItLPeaRaAK3MT1VChqPvzEiRHSx+v
MFFyNW5W3pcBIXpuwMVfM8Rywn7fOkxsX3PdgpHbjyjKvUXIJwMxVc+fjl9uAmFlY9/EFKbju1bj
dgBgKrtBm1j7cm/QErHz91DB9JCj9I/CnMNWeQXbuenYNEjrDcrhRdD+QhIy7TaINx8E/Pvh7PIK
8HZMU1yQeGLyzYdkV7ncZHwuI9N5AaPL8/Fz8HWUcvGZttyTWUtYe7KNRl+ruF0dLYEtk+YOM4XE
fiRC07BfdfGFosOxhCpGXGrlFgcvMHGcCpglZHEanTy+smaU2YcmEMvCg8jy4E+lEwU031VIW3VO
ZQnQEJkO3Tl+p1KOHHOPaO+l+hxdU3rBkwbhOV1S+nDV6AhZ/ZztiXwL2knaxyDj2BfDO8XGkGv5
KxbOktHvvEWpKnfYkGCTANKdA/6PbRbX04UY0tpBgl1hXEAGIDB+7l9aKnZTAAAm6OgPvizCwdlO
jb1W5X30s+yH5hNfqtunLvZgdQGaShjdl5VZIlN+e6x3T6mg2sg+PPFFLvE+idbqvlnafSga/6Oi
VUE0NIHCc3v9lpyKmwZi+7nP9fNsCKgRmd9QBAXwpu6tpViaDn/h3W5R0P5cxNPJTUGZIL/TOaSH
sAmB8hJzqDGuTegurm/MJ2nz3wJCiGiGAQMp+1l7DbDVHq3ovqqMN/nIyqypY0nrBgTZ36kdQClP
pfa9rvlsh1V/L5E7i8qmhCJ+5jRF41kZOy3NTAq4UZNqjmRo3V4SbPcn5aV6W2Wfx25AmQhXAIep
kPuzbeAJI35e2CwQqf/6AYEeg5mkVCW0qDV071j+BGoMfmfP30H/PeHzNRx4yeOHRig4R6cHL8yR
U2Vxpohs+zO80HnV3VWqdH329dcxE8B464pNt62UM8PvEgqeptPV/52nGtky4z0mAyh+hILBjIrs
RmnZ80gCvtJgYhgkxiK7H2uiDSumkA0hFYOd5adZ0xXX4W2GzBmMSAPF+WsnxtjrzlMv7hKdDgQI
VsGHi08P/M+EqFxiEyPzWu0A/5namjs/WLJuskpdX+4MYFEpUGbrEsvBTWVtcsVV6kuRnR8qHWF9
Vpk0WnRlp1BGyxhDsQbb5COA1mLLvvwcHSYGUq9kcLIIYFZPOagAQ7ABYovdQ2hthWaVX+90sOx4
ELO/4uMf3l8KIcgUHqybgPojbgCM8goJ43VVkmH28d+pRbMVgW2EKw5p6ayQ/L8KB3b7IWUFK8WN
ho1lmYwpcxbjt8Bk5E5/u7a/HQK9S60QP7LsbEHhVJmqfGv3MDd2jlhCIBcqjzKqw9T68eNZt/K3
j709mObJ5CGDNfBqAB1qnR1po0b1usR+UwUnD3fkwhxcJ2nFxbThXzcwzktXfLXWYcEENjKisQbd
iKnKfiJ+8HdTcQN8UwxZlzHVHTf3zQP+2wGTD4vWP4/GLoPN+PICksVezc5vXbayf4HSX394WYnR
K6qZWhgn5PTulbD/qHdpWO8CRpSfIqS/LHoMCzihDpzdDroDB0INGzr2z1LwrS9KqOFwsqEuKpS+
mcGsUbOk0rFi/FSnRrI4BDWgOt0EJ8lcGRWGzyFAeO4ar5X6bxr5/uw7vYFBMrsbHU+2MI3uELC2
JA12Wak2zgBrNob/nLgHjqBwjmHwJEo+PD6xYoaAUfjBBI0x0It6bm8qI+al3sMnmuxt4BP9CbuF
ID9Iav3UPLEUvXT5Mrxr6TLLcNcghpQnWAUg6opvtAEPJvqYs7QYRqG8n6hAZU/48/5+kYZCrTdu
829s+B9S4JB1tqZUxFA1q+UufOrvkOmw40M0k6v6V3BVlhyYjpbfVSk+BSiPzKPsfIRnk/PquveO
tzbMNlO4rI2jpJPGBygjCjnquKgdzKkolbiURmo/d1udELV1BalNUT7cs+0RsvfKTxJZY9SY6Pza
xyZ6ApKOxc/aNSPal6PKyw4pYnU60ClkeLasmDjrSQF7+bt5bRKnsQd4LqvO5Dj5iv0zWe/rQF0V
vPzD5Kt7wT52T6OcDTW+Qi7qcAvzkOq2jt+uUOGAafz0vQiXcFhEa5s+0H6daUl++eyAQmWjYGQl
1Clr+NjjFjH3M1U80CRI6WRYhomBuVrXWCCC1b0l6P51SFhvn0mgi9yHZkyO1+jzxjcgL22cvF7d
rzx5GPc0XPxDFOF27xkgqCW9P3snKQke6nnemZBkPwkDjhmPN6zW5uhS1gg4/vzWKknc9E4SY66a
lSX5PXh2Rxmv/rWxxdw69qfR88W+Y8rfCmWeUbfbUZHigIw8egKXatF3tebVqi3HUiVchOFsSWtC
agCMvY8RAJvfS8zAtaIetX1Z1zdqAH+wf5wEFw72qkPaiFu/oznOPA4QeORkdWZSBt7y3z09J72H
mS+F9mS7O5mqr6Pd2UGvA0VgquRE0y1lgTVnN0rwkcLv872nnk22UUoBr8QFOkuym4bAhy4UDMw2
MQkhsh048R36w2hw+oMBl47PKX+xylbaj/KteTTJeAbf5LY/6RLsVPhJd+pPduywih38GiTa2eAp
fereHl9Bghx3imZSwXhxP0hLjBZw0VXOgajtrkH72wiVEQhU9QE8WiyU06yLHmoC+BC/bZc+BWEk
omX90Bne5Zyz5hWoLkF/eO0081yKg7p/HCQQhuyCrRRqiZmGAm//4sDjXzTrs3b8LUAxRNYyZ1YT
5fz2tkscoq+R6M6hR/LHwUDOWsgkxl0MEbabsmb8xdZfLWdywibW52fuZaAivPt6Giazq/zVscxz
ac/fy/5fTyhLzCTrNzY4S10r9P/vnk+1EjlBT9RfjS7Adc0RyIQHTs8dlkqZhWwQAMPR3+7wAPpL
nOp8k/1/b36fzb3mvIU65FGl7J24Ft2kXFS0pPBpXSx46Qak8hP5uEHmlDI5AvrN5bEk++W+foz1
GfFmS3vOHQC5UX/skHQ2L5IG2ipbucOHyB7NN2qJuvR619d38Yha2/Pj3agg+kQ66v2FN7YPc2I9
hKJvXRETSR2fPSo+ifATm7c4tDVJU5+OEztmuD3ukhITGuEx12ZEealK9vSaCX8/H0Lrrhz09o5j
22bRYlYOq/P6yER1ZvuNV64COeHtRCo6lYcgQGUCdBXKq7HEEOY2wLNEk9EIbt3ZJtIWnmoYjomS
LEo9twoCKdMKcjryDByyth8AvSNnXXvNWBuWHWKV1srooorc9ck/GxV5BGGaLXl8Fp3vzM6csdxu
mzYcyn1+n2TTtX/OyP23ZfMH7H4Y39JeCqnW1lZrxvGOpZgp6KM8/OkDa1m4zvTTgvbdvEBw8IEg
2NINap84aViS8izuQ4D+HUzCfOROLvMMgDSzFAYtlzJerbSXWPqhpUw4SNK+NKILl+5a8OSpSy1x
hhLfNQhoUHMD8l1hMW33NbihT3cA5c06vNjBho0JuhW7HgGrK0HLraaaba1UVIvnLatv3t3bQA+l
TpBwTURN3qdlrCIC+Bpx4smq4t4MxECo8fuUpXjbaecbqS02GSwdpYoEWSyFpCTLAWSkslgP3siY
ilVEEhtGQyoDTXVPRpUmmZFhVbELS01PHr1fqR5BQRxqVSIwxNtvgkk/vWx20J47bu4sBNUWIS5K
mweSb5yP/qUJWUPkIzX1/1F6Hegql+cFySl18nZDrGgGNaBz3pyO0TlP0z8FHKE1uWlcfsCJ6c9W
MIsvzZYZgy1IwxrAghbemWq8uQvUCnePkz1ymUv0Fy81ewoX2Us13bhHy2H9fGj+8f+kYmcbd7A6
hkBVaf4UpJWACEnDrlDAU4j6hy41hnUXPaGfftzwyvkoGJoJUe0jN+QyIOmS503mFrKVBbuesCyY
wSIZDAq+z5BXbigZHR4QrFjmDyOEsZuDndUEGuOjImWdXyCs7+7GJO6nz8iB7HFLZP0nBaYY6GAn
Y8UBnweKltVG3PWKKp8gGhZDypdDDMry5lau2VXtfGlkc4YadAFPRRcOHYRrYHeSXNhCKhZEE/Z8
6RgiePKtmU+SSB7NdqS/quXcKOZ7CYO5910Pu3SglXQopOdZnAPaS1HcKiBp3xGbstGI4oJ3DqiH
XGtwv65utV5vZOf8oeIVHDxGuW6kaf9Wsr9W48FI9R7o8h0rkQUBge9NisrAY8oYRZ62ZImPWSfu
wEdQ8PE8mK6MUy484EuYS7Hhasu4ngsGjK+LMLT965jCWP8UDFpDs3FDX02eeMddDAvnj971B8jm
3ZqaXEyC07bB82Natvtvs/8/3Lf9rYjl1oSH76Rt95Beu13MqET+p/D2ipeOLPZu+U8qEoOLjbyT
T8EB2dAXNglKBWxQv6JDBkhGxEdYOjSioPhnfC9uxfU/COaOeYtmwJ2nEjl0V5JBL7bVBM/hCKiw
zFwYUPEjQ32WPi12t42xvfxzg4F5vKIjR/xi8DUOR1IbE8zU+5gHmndAwAutXCuUzx5t+PyemS0i
dzsWsgPbBzp/1ndEdZ/FSZbfFDHd/oQb6a43JVVYJy6XmCpFv01TL7F5wPrz0xJU+wP0xOOPNM/B
n2W3ekqTjwlYJYNuFb7irXT4JtZILrqTe5JKmCla1+AlsDWF4oDD3PzeBy7qNC6SzBYTI+XWPcwV
ofIk5i0NLqhrHQvSFYWx3HymhFjske9Xp9h+eFtN1UrU8QozjmRVpEXk2PmX3XUw6zd0wF9aSfZm
DEI++Qvvj3CH/M1plSO6vPYeZmPhkEIsKl/NVnJl4/6iufDe+tPdaxj0Q2/pJgMAeN2rRFZ80xeX
FT6bgCMo08Ej+df3wpbiVurJc8NF9LKelMLMuhw6tksMk1eGNNT5UR8b2/L2PtZAa5QQvE6muR1H
T1Dfo3PiUapolii5d7ijjq0wcdyxH96N59p5gfC2YurfOGjC3Yxx6sjf/Im4GscspnK8ylWkvl+w
rV/sfVYpLRvQ2oGm1kgbLi7y+LAz91fFT2siBNW56y6LmD4Dup5nBn9u/0ANeMtrn2VHfQ4AXCAu
gq9fG136extvdh8dk5uro3zns41QurD4lNbfQ4av8E+bYvQzeWztTPjNre5JgxlI5fhtaY720N14
aOLi8uAMNo4LhzsQGify5yzTJ1kUuPVFP4yoFU3jBVr53QSByTyRpsjuUFViQyQ1TDLF3WCHSkLJ
5sL0TjJzpXwip7c6vO46uVzaNojfXTXp/1nvQPSbYKWnmvCHM17NGpconc3KIe8O8BDdwcApKnTs
CuxX3xtmqf2ZNWX4elO/mp+zqeM+kMZKQytcddXzURTtwB7de64nMV/d+Ir5CF2UcnacM3MOQUM+
hDhypM8uDJh/RWT31Y6sizoKeSLa8cRfe1KksXveIMhvsxPxCe9UG5oz7Nas3kDFnZf2PSZnYp5f
1XhMR/iJgaCh11+4A1jvBpkYoLV0GuVgTPaLIzzTLyZDEE0n8cvhI3oSDO8ER47hhtJATxcQrK1V
K7VqJv1CiW+oCtF5fiTX4JZTx/pKPGdWTc7Lb/Wa+b3Zd3lwA1lkvGyGtSsUResFrg8cRTBD26zn
jjOs2ZSp3nHfIJGd393rAHa5+ntZ4Fk0L5i+LZ/c55HnlOh7mudD3+/tPkPH8sEjHbXlNQLaYr4q
U0QXYjOtJij4lkZ785/6zdz18FLJeQwWO0WyfgcXmqVhqem30kZdF9XH9jq/M7Y96CgeCJAbL5pt
a5jT/okwixn+KIsk3Y0qUYHRZ2zath0ZSYVlkgWQzVYlm+GdN+UUka5xBX4LLfUQs/U1WzNxJUMF
7LY63tSxbE10sDlAiQBaacizciqF050UbWg4MiilXTsFv/I85zf6ItUUlxsdAWzLDxD6g2NuGAu8
IkLPsKgd1+E8zs+1KKK4kNVakgiS5eebj9dZ7D3LbDnr/1ivwVS99wr9sHcFkb1z+OGGUXlshTKv
tfwTJX0qV2YKwmAL0k9VbEersnAKZCCS4pjKikSL5+VVF+VAmBEjFalvinejJQ/TNvFSfN6hVS41
Ge0TOZ26AQiywt3En8/ckSqZz5riIGJnqrVKEVtzcoVb86MJV6/N+0f6GHsiUnZVcHSSSU+wKxif
BPFWbDIbMANANNOC6daIrVM55bCw+oB1omZgI0uBIT064d0kfYaH60bB/PNSiZy8cgnq1yNrqF/9
3lGkJPULCeFHEll2SO2/8ubLUQO5GicIAAVv9BICEYddJYCD30Brn3eX09KFgPZHYqgTXKxIYFuG
JRqRBW2QvXqplkoKXGGSwYdqNaRWfFOxnvxDCZg70Ehisx9wqDciMG6/jscBGpLAMmrVpSJNX1th
EueJRVpHhHipQLrufXoxsOzRx3S7eMj8b3x9eDiDbM8DUYhX0p38/SwpKeRDUpF1lAw2B4l0p8wD
hdH5nItcj/jH0rmYIvDkMkZXNs78q+wYRxPC1M8L5HEj/svQ4wEsh5uveLU7DpquXOlfPh1HBea9
Z5uZB/KoOHFJbrfbhuimuSkxox/ipeflAPjxErJuBg7xVcwNQiSosN+j8eMA2deTCJ85QssZ5XXt
JzBH+Zvw+OMPrS88gs0rvhtwfhGXf7frIEKbpwH8MyLTxtp14/JqZm1BIrofblRn1xdBqNQdWxcw
2rsvBvjONA3XnDHeeUBNsrdsr3dIhlPHPXsQqV3JJyesXEearktNcb4t7P83XKFmpJdmxYMSMa1K
I3Ff0Hb5KLhabGEpneidNrOI8ClnuvgRMq1ez5Iy76O8ROOPt9Cz42sXm87RNmVy7ydlSmNBEKdO
nIxux90sHQ+NhkE8yiPpsPcAONiwPS1KWUhvh0m6ybqooUT/KEj26TaKiK/hyDWTupbvsjQ12Pey
BtPVNWGArdc2+tUdzY3bBuPrme2WENv0EgNeyWTaexm25P1gkQuCV1GBHSDEKAayl7Iw9w8z2bTg
attjShqmqi/agOHTn4UcBxBYLK92+EPTJObOgEuulwVGZc85T3dP6T65DZ85exNvLTv7u8Pbsf9z
ZM11fWWn/oaj4IKL5z3teob44swziXnCh8BHGHi9agzRCV1thDMqgHWiBdoaUQx4Y8RfgZulVI6M
eDGqtChvfPqjhpKyAS75ZqfbRmgZt3FpImy4a/CMxv0QVWznoJCCH8WSER3vbskMLkNgfNvjaFdM
RDL5r4PEjJ13Auro5BGQWOEgXulr4cdJFuMqMFFkRwbAVHXefzf3mVlMpn6tOOt6L09v6IzH3IvP
ka6brH2t3e4PO9XjL81Vx5MEN97O3DP9Lb4So+06dayEje6Wn0QQPAgpYun4aDMLTMXiVjmjj/bv
eSBGf8u6r/N9eg5Qp0MT5gf+msPzTOVAYy1IYe3MUmg31wcl4E9sCln/2hO5aPp+l3Y4F8yW6TI/
Y8UkMKcsaQrHmjACpquLhgve6GxPKJP5pk/3DU/IovvPgVERe2DIJjqTxpL2k2wilWjlYBTTEvbb
HaN1kN7S7mC3fw3qEAalcSfdVMr4qRfQNK+W6b/u7lWHhNe1yZ3SEAo+stdRNO+sjpNUXkL5d3TL
P5vuNz3rjKKOxylU107HP8paGWWDbWnm0f5/LfJh18BLT4S0Lha1K6bTAr/ZSHTlqHR+aG5u4ybE
4rSMN+LE9U6/OQJN2rJ+lG/JDeiE6fgSPXnzAM033VOjmOmQLEEMJ048X8DQoM1dfNfw60+W2HdA
9FlD+GzsVqdL3v8KWATRJ+8DwDRMEDwWi7SvqUnuBaQGKoz3e1V5BHrUJreAKb8bLbBT8fas4Rb8
mT8W5oT2gNSglqdFxY8JVlzomd7RvYEnoOB0PpEcbfBMBNbu3bsR8aQ++ljnwo05N4U3Wd8Dzo0L
Y0dnyls8TJnKGpj8e06xYXqJ1bQR3PLjVo7UEDBRPRrrjlqQldNcxUhJOzyllwpOaaa1cLiQ5rm5
ryL8JZNOan0zNwxPiOOsF1/Yf2gghhKS/tqb8frJ9lSdPsRaZdhlJN1bAM/B5r7MiEvksbz9orz5
nZpw78s3DOhz37Y0ux1/aUIzjIWYrB3xlyANohFRRZoQGEBtnIjiD6OzXuAxOTqZ4Tm/r9MiNfwO
y270uo3AnQWI2JrGvQU+s9tFLY7yzZH7VAUnUHdapPitseAfopbqJm2w8Brww9C4IYe7sp/YLq+k
GX1dmUqBMAmKG8qTh+/wTteoJTDByKVug+CSgOgieAgq7lfVjf5/gRfhvCBrmpNXcuHiMPEcqRyv
JZ3cCBcApd6kqrdrfLRTtDgBxu2M+JxdH3Yf9lbuOu8wm1SghLtzxWab7eQv+RFUaVAPAhR5MwE8
ngMfWDM5UKQpNfR9gJa4feGN3a8luNqojM21oYr9ZUyUEc9Kzw8OJcm0MPgKtCgDZhlpse1csrbh
qI/cf4gDwsMPVXLsmGkCqbJ8WCU+/3iv1B5sPYPo22jlmRUFc06cntdFLBI7qkrT1Cn+E8WqTqQ9
nnsRF1f1/54//FtrLhrBzSdqxpQTdvqx5gv/5qkVKte/ctnZhhI0WuntVwOjOQCeF7R1MddrWWcn
jd9wUdhcnXQ9pteFnuLr4fh+C0PbliiLvwjOSfh6oY/wT9n19O8QtdHg0BLntJks8pgSUxcKZ7k2
pYjqFKI1wF/dfm/nVv8BuIbYjoepWvOWUWP8sFpiyqiIB/n+qm8dBFHRchwVL1zOPUzECdJUkdUn
Kyocao1OzNyNFwILUtWVicSzL11SsiaY8Pp6nytR2BEl4d9VQfhO1gLv5pTenVoxBWsJZjtSRE70
S1sfEHb8hi8YKKuVXMQYmjphrcIB1Wqbd3kekcTIsQIoln45nI9iz0HC1OK88tIwaT4eEIDNt/zr
kt5IJSbMlQSfeRY1tqSVWHcr3PEuG8muLmFRJV4vk7vnfjSjhEBfe5UotNkJ75Bv+7TPsJ7Hz2zE
S61/5PILb7vtlR4aGTP2HLaRxTiadHoAf2AwFPnurTTOh+qwuY7ThrMwz52fchZCky1l9L2XYMbO
vKCKGIo1WFt+/b9xNTLcSnd6WaLstTVEn7fI9M0smWhpOBk0BVEKLXZYlZQ0LEkeiH0d7V+jnHUk
+tMGsPIDCd/6p/ytLBO9BfsmJ7RhV+OaPIyy1eA1dA+4Q1fNq3FRB4BsRC62zxPOdNDh0a2cPAX+
gTzb03Y9EPY9uV7NwqvoGTDByzGfvrJQpA10WWLwM5DjHncYItJosgsEXMp3CMi9eTXo8QJreMqB
BgMO3/GxoRc6TUtmdkOhUV3ZG9peyXT1p+aqt0J46408xRz3phlMw1Uj9sy2DlOsdSigF9BB2jpL
6usQsvlOPzY+2dSHHCgj/iaIkGVjdgyd5RWQU6x2v8Wola1o9xpUT88UUIauYC6wI96BJR5scjUp
hV+baiMajCgEJnXcsQYOSeqSaz+tG9DY7Xq8+4SkSF2dkdetl8gBGcjJkgUya2FS0DVZenj5jcRb
UMcosM4E0Rq9VLprTSeDtEG/pyPxf9iIyJnXHckbx4v3NnwkNH8hdLPgFfN52bsGadCC5iybYJCf
9c94a5SeFlgZEuYHrfuyE/1ZagTOMwkrw2+a/+oKuDXttUORZ6b9m8/GByU4pg6DpZX1DL/jmkYQ
S1BajVNkOVbGtr9XnaGYKjRq3Ivc5kzaTNzIpLS8ZGKjL1tmhAocPoqZLvHx1DBj5kiCZowsodKL
Vhm+Zkm0V9AZYMmPiSsfbzhvWzop5WcMRg5cYNkMYKHlFWwvNxe9VgjQn8j5noGbfLyg0td8Z/IC
ABNLNbzkXabEZV9sJ4viZ8VsacVYyLGwOyNcWgmNE+fzopo1cD2UHBEacgzuz3MLlCKxj7vgCQ94
y4R6EZ2ZIID+SS/CPhChl4bTW3GTAivj4LRjJHTczrHI1BrPvhxrU0vQkthmNDFpTiwRI/w6q4Hx
4p7ox9GKgxyOoTlS6v+9mAzibaJ0VumbqC4ciKoUwlfBVHmTRxFDeWi7dyaM/ZCsbzuggTrMJmH3
8UhYGC1a3P3otxlWgClHiVZbQz47qeyzaEc0AM8q8C7qLm1bWtu8ZI5lSi/CwgCVRT4Atwa895wd
KmtA1zh09rmA/kz4REJ3lM0cvtdDAMjq00nZB32mK2EqW/WYHdwuH8MSKO+qXuh/QH1kQi8R5xmj
qEpeQJJTAK+3XqI2gK8bpLsEZLb1X/96Z9OYXkYEdg/FLKKe046yVWnhFSITSwyxPIcW3SL+aPp4
vGOBl7BCwynESsL0JDhp+RkKiKYlyDCAbnthEp7nAFjDyMIBHt8HsFq5MG0lGQPyfTP4wuwXvb4h
BBro0zBVyXlzeGidzK6dCoujX3B77WaNOCdHX6N51JzMNjsjdUadlmCiBYCx9gETF7tV/+w51DRT
ct7i8vIofNzObk6xwobHT7Do3Jsqvf71d/rUPcVOFtVceerEkDbf+pL0b2wcya2s+S5i69qs9se2
+TSzC8Rui4h7cDC0zeyWYObKm2qyt7OQyOR0XO3TF0XOPqf/m8ZoFP8YHc6pBaY7DuMUrz87+SY7
gF5YaLMiL4yo4kbTZ9zKz0XS7Lb8SsYu/pGnBf7q6I+iB6ZgaKEyk3DAHdNrP1zrFMzcqYcPkmHl
WgBMtSgWREqo7fLxICAllg5LoBycjmiEst3Z5c7eNwS338gYay8+kqds9bSVW40KEaImmgEPrn0C
zd7l+1El548iRbVsQAO1E9ornzsEzooCzrxwq6ROllBgmN3cieJsenciEj89nE+RaWFmRNz7Kap1
qdTCj9m3cLQijmnS8hhaOqOj0lwtUAW0/u+XVand6hZf8sqkM6wmxH29y4BqlVf7bZEaVJucODWw
IQuusPnM4M2uFBrRESJTA6wBgu7EEDqAnRxG+F1hiULln31eNw4RreVszBXpIo0k3C9YPkcwXTWg
FIdQlZIp3P/COwTAeSwLKofe5ROeA3F8eMtyKK8wQOMmIEfX/O39QqibiB73nSiSvjOodnrBKepv
8upw4O+hr2H5jnKnZWVuuHwlSFv1QIQ2e6aLMxOxWFLOadCgmMrQpwhfPZAysAZAKZD2gwfRz8ax
2ckKSoWqne2Z9l1NWEDzKtDdPFlDOGWkfqNdxSUbNPFmVdq8ZMF/OPmVW06gjMmsak+Ex7DDDc/o
iQvNJBdSQLgJAR1mn6/URtXg+NqyYZWx7OicNolT/ic96zjcwV5MWZU2YlX5hGbF6zCP32HJZF1x
kQBuW8MUa68iM6m+Yf+nmXb6jwa2TuYouZHpQS58nnaF2sAFqb9p4BxMZ+szBAMwa8b1BXA8IzdR
ppDPt+k88rinc6692iKMuEbbsCUZo9uuLz7wpeupR4j0nFm2lk3gLZEtaz74uzpGo9Nk5SOX/hyY
rTtXnGuRgtkWUWk9uTqaPvKDyeo8ruSdI0UMKHTaf+WadGPYyg4Fj2Is8G0xLOeo1YdOz2alZQT6
4wW4dqdxoUii/R2QQ91p6B1mZC/O5zkTTkJVorLweZ8CZEaMxHRUrNEvgnUbVlHpF07BBqCmFARQ
KijwKs5aC+Tjdys4eNUP4nsRt+POr8p3zBrN36sXckBLV7G1TdIkliYveSBW+wVce+zZEYZuqU8L
Sv2pRTfc2LhxLxuYj8xaIGT03USDXz91dwLvhRjVmlW2IIgu2wfKK8bb5cOrzTfizUm6/Z/CZeac
Fo6jOq3H0XIKcJovBV62y9USTglul9/srIhYkUJiFqXpo3l5N51duEXZczmPIqKxsoH9XVImjB9n
KUOJlV9sNwugl0OWyMpdzg/qFY4p3qnBwCr1CuJZWPW5FPWGBZqOemsFwjsnByWso726pMO2AxQW
aJLL/P1FqSXxfC5ZJ949p+TD6GRYfmUjJb0Rq3iRfb6mkQRX+C+2UxifuosK30HUx0BHoy3AmlDZ
tMaLKiS73sgC07CEIb+sgK8RhcIE+Xr+/acBbOSiJPPtRJfCbEC8tUdvvkxhKUhtj9oTAeZD/r5q
PhjE5FmDpdvU/PuNC02COH/X9xJr6m0A4dccJw37E9btgFJ571zJzDpaSHEc0e+8vSl81vOwndOO
S1jF+t3io4BzSMbRNTDGrHgxszksnGwgzFRcZ5EMxxPjaza1sSBicwwv3vEr24smoSw7v/GMkPAj
ISWO6mVLQKVZenNh0s/WLGV5/ocRcyN391WXn1ggGx5gYdJ7R/2nfLz47oZZAfuoJRM7QybGsEUp
90BdbAsPqmkmlMiNZguHA84gfWP3zIblHtcfHq/hXvucmV76qCYIfL+aPEwRwoeennD55RG6qg3v
dOrUqwfgrY7eOxCTjn4FKSZ1XzwFqe86JxcLQ3Qbrm3g8vovrjLN++CG5dBHDiBUeJFeou0bXxpX
b97PXs/2/aTjqN/OfAorJI7aeP9jvG6a2yc/hW+sGAMWmyrvcZ9EeJU4JzTHlRoYg0odmllTC8OT
fowZL4oaJh7TVyCyehA2w9ZHKO40a7pYowDgG3zM2XqjewXA63l4a6mIVYHxI92dE5cd/vc94xwS
9rYOvKJH2iyGNaEdByXA8/iSIaYNuVtDGcKnfZi69pjoQsdoo1whKPbvCHSYFKZvAMGM6AOzuiqz
x9nizV3H9zGIWh6PFYy+8vf9u+CWm8Vl5T/VVEyRRsEmAe5u8+x3BpYILQQ6lYXOmAA5w1Z/KBTt
Zmi2pxHsGQd4Zc13M5mtd5jO94SeqcvqPOIIDBDjS3Fxilm7WawQxhlMcg5yoskGWUu21t7EeOpi
XrzyDRZo/r03B2svA/sKv0OFZdMzZK+t0OdYgxW88trIlUaFjT0fBMjtF4PzkjFhVlKZSAChsb+Q
uCnN5Eyr+dLoaKFhz9bYve3BnjK6XF2goNaicXon1i0baNljbPh0kih7rrup6FJKwjYE2b9sC48W
Yb5PvoecCCwK5MwH9mO9MtnRlOLYkQkg0Lv0ie9RuONG5p8lGz5/KSZVf2Nk/bJEP06sc6zdll4r
wciPTi5dcswQXqJ1Chsh/4mbeugXM91OxsCZtK3U/mA6VPFArxzc22MnA2zPkwCSpfibggoGjbm5
gRf/s9x53k1Z+Fxsx0b/jSY3RTDMQ0OCRphioXDQIa1YvElA79BjUWYIFBWJ5zf0AlOXVLtBb6rA
lM4GwzdzrNPH5xIB2ib/8B1eQO7qzRHl0upxulUyamA6CeD5IJf7kcyti+tZdJhi1UWV4FfQSyaG
JlVjzp1k3ZSpZqoLUac19MfUXT+8Cfys7fP0nGRqygEcXFX69M7ZglS1ITQ4deQ0Rqx8f+86DccI
26F1QP5NHsBv1ub+m2EDEzqIhHY0ltyIeTCefCPUS6jpq5aNAVa1rXKI8PWgwlVdbkCBzRPpFsOr
1OQ5X8CSnmjGs5/pU+V1QTJZJi8myDNaNyFzDK32ebm/SPzlxrSIIjzR41ledyalFvGFjaqzSM1Q
vJZkQEiIi6h8tg/Dh+Nan/OQ+nQK+bx7MCUgQvMLz6TUPRv6l36OBKqeixEc7WgJwiZupHbxriyE
pjrSgkKX9kHmhdI1/9WEaP5B8O9//whNGCA/lQSBotNHbu5EV3MsJYtkgR7qiBC9Vt2cSceMbggY
LPf0C2Ws4HPllu6pU0EijQe8/A8zFNZn0bOVqF61UJP1kfMqaS6ZF23tUCaxU9/BGMoyaodm429e
aI0CX8groqrzqtTy7pNW1tRXDfoNvx0zvaSP0OXwUCv2b0bdwW+shubNa9ZtyIv84z4NV28xwpml
7AgJeK+RcbzhVmXj50Rs9nZqe1HxuF1jSteZgygUDPNXDHr4Gxz6ww29AgpqifY1IRazZm3MLfya
T2oMfHTRE0bc4wh1fnEt5ZGkCVYfmsqB6z0eV5UvwEKEs1+HR448ciHkpSWer3ThKDiO5ask2YZF
zT8Ttwx1fKAxBe7V+PDcdJRqPXPvxQ/un2UkeptsU2KVsUPfxSRDE9EjXbPsg6RL/n40JSVkKjIt
3smzJInIvuG1zEaj6Rvq3XoD4EjjY1ldWVtOQZg+W37cKODzxG90IeoJWfOSrSWbPhg51LzOWdQW
HRlA+4mSKnKewzJxIHiUO/JUGrl2fFJvnpI+pAB+3TDAP+mwYtieV183Dp0gVNYIAL3+6x4qAv2D
NNqixbQizXglKe9by0UOVFtgkdKBQ6uKW7U6V3VSuT5mbUfvFT2K1Gzu5hrBY0SHtk4b7UwU3KtC
xOtbtkS5Hl+MhvGkGYOJHYZ+R97gmVsl9JocAo2JjyH1TfGXdtJto/Js0THT1L7ThmYpAxxUZoY5
zuqV3FCrT8KL8DJgb0xvCwu8tlJiT4uwodMmQFyCnXrIe4lsfuBI0I7L9jYW44sOTGvxFcWa3WPL
drBE3onaxM9+vI5Cm1n1cfAm2qDktjwUgDFIA6VmwuHMyckVpLjd1L+oh3QTU0dpFTJawTE7TVS0
dY+VPEjhoItt1Cjqow12dz+e5Nekb5+DpxXY7ZQKV9ClRRQNHczDQ2m9Gd6+uYBnHRd+4Mn9b43u
2OrUlzwLGHNSlQKSbLJ+Yx5JSj+C3wWFXYDkvgeKTYVQ3V3TthV/xF2WyopqD7ZNmuA5INsdZSEN
RR/MtHuhk2xpdL766hM12NAY6xZMZ+wmgV3qGGPyqxkJeXiMffAsMuO7h8hy+GVlWfYHK8YyTpC3
cj2dnNzokK+4PArNCQjfbtnywfoPhilfwkxQDJMiKa5UY+lHmixWnk7i83lDfy31R0sdkn0r14NI
4ml2FgqUC2ZZJJ7jjjO2kDxpslfWhD6EHgbz6IZeVizBnR2EaoSwvmMn+cB+rcFkfw+LMvg27Cvm
NC5pseBTC7tzLoGCTI8bip2o36rT4gw0oY8++7VVBdkk+U73nOjRTwp6OYt24SQEln81/Vd/6kX4
fB7ZpoVtonvotcZr3oW+C3iMrQHsBgaLDeTZT6LWIhZUaQD/9yXGPhwjqt4tuAWVWqBHpnsTX7NI
UggEw6g0qkF2ekM02MYqidmP9GFemEc+a2iqs9ud5c2sslidbIb7uB3SmjupeUD/DpfCcfs3eF/7
OIRXFCjRJoKWJKXZaQ1E/OooXteElGou2gEfbJ/RDyR7NiaOQ18fdrJz7qYnyoAj8ex02KjUseKP
SrA9dkgpCWtOME0lRkQI/PoBwNoDYmQ3ltrKZrRLPLTgb4WBAMQB/QyEpYJOEY+hJMfOjzpKVUAy
aVa99qTv54PnTtx0XfTkhbpywimfgkGC/usj6HspEJP9iTSfa8uLOM4ltHwwWnhN8zeDBvu7QnKb
fzOhg5Ao7s7KJlm8NZ2CmW6g7kz0Nk5hQ94HqhVjochiJ3yll3Gc+B69xoZO3Rai7UjD3xQUq/2k
MOhfh9xNjP7m5da35grrXsTo8MPNIVMC9A+EyyXO4KYLhNKW19feSpTzsuxix/44L9XRJKdy+lU3
eO6ZEyfl8TILdjsAwGPbbGLx+pZXrZGTnlXHPh21PEuXrGHMKjr0eytmngYbynvo2Qch/RDB7yDi
BFuPQHVfOs8duyPFxbm1ARvbcuz6gnqx60f2rGRfovHvUo3tIHh+jMAo1aqaASRNjvNqRjWXQDCS
PLrtaXBMf8W2ejkxqzwplNUVHZ9OGL7LMyWU6DqvDV+eV1uVqIytRQNFfCSIL49O+1F2m02bhQze
iZTQ7Qpjs9zqSnwi0lCtFCvqJW41cYoHs+ijfg+KvFphRgRGou175s0MbI/SS4CZbLbefwoQXUOU
ZYE7Eu++p6Uc89wg8jfMeLR532Pd8dQqpdEXRvmvKf91jpoTC5Ftx9KLqeLmUUedugGsIBtqqmN/
bfEcoCAgM3BBryhti3wFfS2SKmpQXnQB21bKzS/WUQbbaWjXjAwMEt8bFSk8T7iyI987F9+F+Its
MswQzTMJcQZG4FzCTkppuWUMah1T/3M6yQs782klUN4PHJty94ROYZrZnjIm86syPkDZPmOf4dYY
LcZBfxOKv6kpCMY8ATILIPmof23AsxwAFq1FTnc7fzsn1JZC/J6AOXKf+AM/F6LpOtrVu+dzjayw
bDaWXaAAV034A+OHD6uovTFDghxO9V/0Jkwc/UqOhIgXfzCsHQKBARbdkkfYJ6BI3xBWCTtMzxAr
GPjIyQSmzXIpO10qi9HNPwLTv6XoMU6g2c9Qv2V58OgzLoNNFHjnAemy5Zvs3cL7AuqnSOKNHmUg
WplYy2e29ZcABk8fS1+nw5WJGK90Qqs9zPXCy7lfzt59gf8ZdFPKGL4kmbgPqz8skpBHD/4b8Ie4
eOW+QyN/GNFdpjt10gHRlq5wsN5yjIn1cLqP1EgdSI77mDcKEX8jfOtlL4wfjidaIDJjF1keBB9P
69eGOAs5fUSHZQtU68iDSpqZFC5Rr/58WSe1SFaT6wpdenTll2THVAZ7DM/pmUETMMrBVzF51q/n
e+Ib4SSx1gcBaB1DjXIaRPA5+9vPJJwM/g+fHWvPH/k25fC7m63nKZez4VkH1PqhSYJvEVllkIUR
Jf8gWwS0VyfNDHEv2QB10NkrFPX4VzMeUcNt3oA1pxO9NB6qW04h+qgXdeMFR39qoRx6uFbB1jTE
er/f6Ono+FRKjoLJ5G/ExRByUki3WxUPEeyvqNmdZ/VoC3i5fsFuZhmAuXG024WwwKPmzrVx+i7m
L+6RXBtXQfGhpFZHgqvbvnBNuYVGZFNJ8nz+9r7yVFW99B0Gcd/YQvUetijpIKeebRQMC5NudOBh
EXuc3eQYqw1kEGhcM250ZIe/niRyw/gDz3PolkyXYIbHwT0rVwZbfVTJoZjT54m1hKn/neaihIgS
Qt02eU5puPOh/bwG5YDPtVLeYM8kwt1Cjq+oeU/VkcXcAu9wkhXKXfy17AdGvbgICZye59juLglP
BBKT5j50jGJMEAtHb9hUWVdMjkqca0UPY9fHcv0jXMZ1Qqe42fr+/IYm0OjMRv4XuCi40fMOGNOe
pDaGuLOnbYlHpqfNJn2CeG3Ifi5Mo21/6F5d3m5V2AzrTlH4YuUqTocYPZB97uzFvHJd9uqWMJsi
QxLKN9yelyYPIqNm8J8DOTyBNKPmv/qNMQzP2nLBhW9KVNKMYG4aS88lsm/HdxxjbCjjglKW8fhU
c6pmhYPYORf4FPMvN28BJw4jIAtnfy3ReUrpVWuR66MGKw/OvC/P0fXi2/tUOCF4OHVCv0dB1WIo
qrMz0k1IFSjFLfN4VkHutfJO+wjweYeeewa7zcU+qPZX7RrADv9o2PtjV20B7DJbgP6xTMM4//ME
bGh/YkdrWWVPIHJJ8J8CAq9gFC4whnsYfWaGRs04Tgrk8KaBaANd+qB1xujuY3Su9Gw3cNxyB3OV
Pom/MWjAogJB4XVRu7kpqtvdVYubEycWvTsGBtYwGUUHjGl9F1uqtpYUtHQNGElIlNdhh466W1Em
b/KIh9HF/cuno2fIcSNOq8ux6X7PnhH3A47YMI1bSRhrRZTLkULSFKeMFzsrss36YBCCD8SuIVfX
XYiCAAV5Mc06NRtstHe5mjg2ofj4t7oYzViK1jl/DspgwApF0MHO3IS3fpZm16tJP2Foa7IBLc4P
Ukmr5GpFdCWXTV4ZSPwqKyPqZIb1el11Zx+fe64Z6W/dKZyRzJloPZutjUYg6on5r3lEjrO8aR/+
iRgzMsvQcslrJ8CuIkxk8PjGDQ2p4jP3SMvQtVoFy6qxIe9AnZAgP3U9eWHAE0SLAviFXHHjOfU/
vQ++nb9vRt7FJNTMNhADZ5MUZAm8Un5UT0YiYgjUyiA5EX/Nigyl7vzPUSMy2j4ZT13Sa7L3ZIr6
KAjxFSXdCalkjcFiHjlwn+oVqZg2B1cL/vbdYNVNV+N7VKCcrRviO+p+A6glu0p4VxKKYa0sJ0JO
oUoHZ3kYQRd7StoahE5k/AvQJzsby/ID/whMMIvJjEnCGjcYPkKSjbL/ht6GbVFdZv+qk7kyh/T6
qOC/35CkW1BPhgd/gITpPVWUcFg7SvkKESLuH5yjxhmlOeV1EsNPHauBWvQW9DyvOA8nCXlu+8I7
Y/6iBtBACLJKiCynO6a94QawGZw2F9aSes5PM8nThsfHe3ADYeVj9NT35xHVMUnsi2A6aLBVQg09
J9H5kcOsbxEPwlRWfZ3QPjGkDuUhT9F8hlvcOdk+reheEDKWrfisBexYR/S0N7U1wJMqyLGlgUTt
xSfTaIf12CZocf3g2SnQ2Ii9dlVOXpoXs10LytcpCD5W31mqjJOBGQdIBFkd6v9hRuPN1f9KylnV
ChCQ3Np/U/imlbfoJEBsG1vnhVgl/q1bSwWmnCwibqFMhHwPQ91e1OFzsJx0VVBdYxsrcBDG/bIS
M52U7HXKgs21t+hDV+HDFgXwnyTaz4aJf2jilPbTrNqZDtH3N2agO1XkHnCtZsVHT2k5w5yuQDfw
ITKp/h6qVqYJP/i+QY0dGtvrHKFL2bEkjkTeOepgAcwpReBmEDvJTvL2bztpJMHG00IjH18nP+kA
Ol/gOjV2MD2m1/Aq7+N2hSLqyXBJ7FY+9jkEQ97qgG+DRPpuML/F5+DAbIZSraN2CojaS45T1ctL
NlRzWA6ML1juHhEk/GbC7UTHeA64TZaxQhYa56cOvddanrgubU8K8iwZBLqjkfHx9NK0GYd23PKE
AEajV4cV8QG4zcOOVCTiSN+ej20aE/XIy4G9WFILwUMEPJYk7oMoCPoExVj9S+FkdkAuIJlcdyrO
18dd72lQJ2zl4liuzOPXDug2++JA/plKN51YFz2jKKcEbQ28vEf+oSAbcX8DW4rOiqxVsmyc/rkd
eel7RIHknKFuPES/9E6PeqR25jgC+eRRin1NBYxSwkuLxsLa4X712ZnOLXDrsLJ4MN+OOFHgsNxc
Lc92rXG6RYY91U4vOlGOWYlRo+E5NI8H1Se3oVREzbVN8oAaTsHPlLrf0hF4URCsoKf3N76GYew+
w2FHgubPRwgcUVWa/SKUZD9a2uRT9z6k5GPsl19Mc+380BGZ/yXnQfUFm7w61QWHL/XH+bX1I5NL
hf5fQ1mT7j8H7rHvuaJtySCYm8kGrlhIvpe3d3MMM3ezx0lNogdv0HxJrf/FznPwd+TZOLUYjprM
N7L0Ziq5kA2w2yyRfGPHTuBnNYqGGBHXTiJnIyiHYdggo3XZPILq8OiAj6dfbtpMLLFl9p3T4Ns4
rZaT9Q0MEd2ajUYuJJihUJu564yfnxgWjcuP/G6kkyB8zJNYYKqsQqztHE5zRewJZJ+59irOl7DJ
1KHBdBE1d5kCpkw+XrqGUo390g50kQnVZ65K3+4bqxNBR44wxqW322FzGtl2Wsq+yasN/gb80iW5
e1AMVNXmT5VHc+of5gi3fLfOTqK/4GJ9deRNyhBP9wvoldyQvEOSEKb/6hHFLpJ02mX5NfwYCfTg
42xslJ1odDucPQ2MR48gDyeFRRzceU3X8FinSs2Wj4H8s7GeLNwj9+UrPyWdJCqlDMXQA+o97aLR
M8lzw3NTuoLtvonbwJUvXCcuJSDqfsjuTfiaKTU6G7qiJsnN5f5k/UR6cUHOtCnJ2xt77ye5FRwY
PTkyBEQceDq+lkFXX0GnnBRZXDDas/nXlPjQb51RIpVIVFA6joqeLtrUbt0yai5hcxDdRt58SWJ1
JFKs3zfNYneIdh/T/7eycWcD/7crklYPWvqLwIrAX3XkZwhAge7nl7gZ/47XoAmjxj0QmS77mT7k
aYs/PmpXpehq5dX74NzjNBN3shG6GZ7QF9RdgTSYFflDDb4F4k3xPZ48hidF4HreEsSGZ+TjlRyv
MC0RdI32zUcyONbRNk6nNc5IKHhHUjgs4QuK6EEeUUL9Vxr3LBI5QTiQ5WwoSwZLCwIi/fHtGX2U
vN6UI9xe8OcLrfE3KHngRthNKn7Xu4fA6jqHnOEflW5XPHas84XGlMT/6SYHGphhaBIkfPGcJS7G
Oi0Q21WuA3MMnMw1KwUedH4TdC4XE78kWnG1PV2VYtBCQC5M7a1fNmnlG1vSIiqTWHX8VUHqET4H
S+HbFSwF8MweuaXbTjM/C03PIw76v1L6PDrdo1eqngrhxLs4Nsqui8Pz2Turh/LDkLyqaiLkAsHC
i22X/ExLEOHHWyrcQY8gzBasiHbFU61g11aRhq/hDWzUL0lju9V21/gIfAinpE9roZUilboakcE2
78I+usA3GPueMS5HKGJdKQBjMWKQ4DJExQBZVTEST9BYuP1IzrX0Dok4I4lguAeE0cG6dGIvMIeO
vKgVsGqU34Bx9NoYxBF2uPXueoV7BsDvSz7guGIh8XZK3lnoJiYla/sJFkDk7P4t+5MCUIRSpU/p
FM4BNIo22MJ+onoKty+Br4ldzMx6kknVorILdmT7AD/SDybJausKYLG5yHnKMEjsyKsnjwavlNLF
bqNwFy5Fx/Xy4MshVMyx9fqUCFWJZk3uHZIiAzCv0mIfgAp7ah8Um9speEVbFYiejVbtAvXQqx+3
I/mfA7Z5IUSKRFqi7y9Fd3yj/KwBe/HM6lE/IziOCSaEUZA4LIcHdd57uxwRB0aMnnm/MyHdC19+
stiClJaXZoFIDFpduEMPaxhLRHMY6e+98jZta/OBsTXvuaWq7q6T9EAJz3dX8coHypSn/8D719Ln
nAZcs6IyZ9STfOrs2WqbhRvvkmSb8t0ntFH4SE7yvjnljBrQjyaak/ZHGCKpzV02H0DpDFAHBmC0
/D2JktTJEDnQyRWWk02Ql9guY+qtpen0yym0Kmkd2yZ+q7tiUgHnf12uWNYqi7ZLmU9U1e7ljf3B
yeb5QEt2yEtBtErWVuGPlQDYcIhYLBJq8bIganAhszus0Ffi/nM7ez0lPIJWXs1SJ0/yENFX9E/t
g/ZE8HBHEcpEiX0plryh9T/X80iT+AS/qvXxb60JcKdTF4HZrJzkDDcMoFuY6cEuRcQeFlh6xvrS
kb7eglyxUz0ZY5djFZw8ZhfrywVeU9+vWR8zIssWAKbQFW6aEs13fAXC8O4rNYvj/h+skDOsQgMT
PcuxHMGKb2NzJwoWah2kHF/fU2KDjRGnSLDUvY5xttG6STX/e5Oety/yhImmsPVfcIGTLY1A6GYE
ATFBXw+MairoTTYnDS8Giz63zQCY4oZqyJFXIukzQYKRqX3qrE+vjaAxKiofJXOJtP3Yf29W5nmc
IqBdG65phdKm5kLnLnss2isdKvzv54QSN/s4ouhDLn3YgK1sdhNYZq3XvsEj6xKtL0oqwM9sbQXs
XfDZrCa+gLDRLJ2e0X6TRdQo30qZkuKOSkjvWpUMtfw2b395rR32pRHClZWs7WkLlNse1dYCW7Z6
mJgwo2zdYwWFM+c2OZDhiIVcFG0VHS54ZaYp/zPisKteIbetT3du5wDCdV4t6P9WIApUNT2rHQ/R
E8/P+eCRKytIO8Ts18JGPPEQvom3DCrXn14eCIyWzf//1eokmZrWe1VQPAn3lORDv4VKDq4R3S3t
8UMvtTJZCMawcv5EMddaaj1fHNR2dnAq4IznIAi5+Q4edFwDj4+bnUegA0F5Ggd593Y+XcjMkvif
UROoTBbjF+QhfEZMJRcEDOQpUNAsgMBecQIpHrHAUUFwlIRjoHTsnGtzPaMxALJj9fjtiq5Z90WI
OexK+kxtZocZuIXjHeVI+yjl00YDDD8ps2RKEohIzAKHDPjS+GMZ83Jw+WJoIDR0aMOdzorjIYWz
GhEIff/UoOmfNsVBAkK4E9ZnCKYrKjjTP73UrS+o+Za72frNb4cXWTWnnk0p/rK2+lajrqH0S1Ea
YGmqjOHciXWD2SdkQEQoJ2qlDJ6VyiEYjPfA7GY1Akf+0n0WdLLrkH0mOjnqCIHuiG+UKLYI+SIU
EcXRqr0CI4/Es4ay5qO93TgeLJL1zMtM0i9OfDmCjzq7x7/KXUxFdrDA5LZwskiviuPnvirrFZ/Q
NA01qELoj5BLfJ6wU4v11XtmBIoaE/QPIrywtNdpAXQeWAsT+Q/9sBI9mD4Xe3Ere0rFn3gv8lkE
E4ySDm+OO8fXPP6LYKRwejFwhOYMot82IrF4IYxsu+FUaZjbUIZ8RSlaKsRd/Y9JEdMX36SK9ZFx
F4njDTqTSieRK2aDMEWpciF7ByEzGSiKLXiONfuZzswcXmDkIL+9bQLJZ0UHyR/fAPfdZzF3jxP5
RpbqhNufh2Kw3yC2vBiPkCCTMbCPtVJHogc9YHb/cfwdhM6fSJyQe0sOrpXzEe7YH9XI0/TtCe25
9Te8cAADe3hm8m5mUe9y3N4H8Zv241mGWu7YIuQytx6+hOhmpa8o/zNfEeHkvkgv9FV6JLu6v0LR
lBIfZvDOeUQ+zlt/y12bdSg5hvtJpSclt6Pbfv5mZRPie7MN1SzE1AYwSXFbUjzOj4wi4iiRsxKW
JH2AuHwe5si8cW7lCHllUi9yci9El/CGTWN83SAlM7DDGuXw1598RNM3TPWg0UHjV642sRbwvciH
pONyORfhebFj8IsSGwh0IrCMPmlJJ+pnz3NeCmYi9VvEw0GtpOgIRtIKMfDd6gSRacSJrnpbltyv
rDo+ojDcKpzlYUAf5DIyLMAWlwqg6aZzpE11xp0IxoEgvD/GNPLEmb7wmFtBZOT7pgqPKXnU1Lf6
B2nOoCPN+Ag9TX9mehNEy2pNR4t1s+gNUrzxQLzVkSQFAgyTbQ5VPZPWcs8uNLOWX9M14uhnbcpD
wqVso1QkfkKwyfsyO9zKPMWbQzbWlJKpwDZISspx3cYvQBqEVjP7Ahx8y/3xiCOqvtV/tgf/7lRZ
FaFOtGY3kyV8UQMJvns0U+O4h802pFP3eM53OH8/fmQWpLan5QBInvJNuyK/II0d+hDXuh2/7XTt
lPHDFuhjQSOGnHcSSDqO8+egBvLKJpSRzwxGZ2pUihOHnXjwybKL9HVj20C1IrTlRiemTuX/JXDc
U7a0FyZtQMf1PRNlYvVT6VzSHrGTSISERs1iDKpk6OIyJ9sA+s84n8TgqzJTxxOADUQnRsL2hYrg
QFpzoeXOoNfRq1yeGTUJaDLqWCSGmjtXcft9jKrukLLrh03c5J5jX8U9J2SyQHEKur8lnbHM4Iab
STYu8KRWsKywfXf1FrfDz1L4EB08IIYP75RJI1z4SJLxk0RPJT7hie1WCgZ2jOD2Ew1e7bJBbCcv
IB9lngpGOXfq7T7mrTwVlPHCYdEKeUCbTKr8r1pQ/cgydA99/pV5XagI97lR2+EyilMgKXwL6BRB
cDO1wA/SJphrCWOdaBhR9qA1fY2iBRZJAoDnLuADv7Hq5/2xiqaBADToSAioK4K1OXAADytTOb/n
pK5lmmTrazeqB/ErzPwVKTxBWPUNhuj62fqDfA4nwB3CQ/3J8oZPZb2VMxHSasgYbEg0A0FEdZ75
lERsRfejfIOCwgvkxdaXlXPf0UTXU838ynhlHN36UMwqUWcDNPkMT2H8atvdlPCznhpqd85v98Ny
k13zBfMYzY41vaLobZcparZo6neTSnNB9JavXyPF4Hv+hpPMhprAII5mbWKH64u0VmOmbF+OQr2q
NsAV2p11U4n4TUI+YJ90Y00+wM8uXGZqrVgJkZN9W630OhEBqLX/bBbFggWKbc5leSAPmMy9Wtcq
jI0UecxcYdJOIRxsOqEMPgmwxHWx2qJF4B4nTJt5emBq73TP4rRKpWm5q9ykFI9ICBBQ/jsOuKvH
8XGrENna3LoI9ScZulNEDQhXN+es8tXt+A/E+HqGaBYU7QhH0IToPC5odreb2M2E2nKLW2o2ZBac
JPvseF3ZQHbO0nBAWMhHeCLrUqSuCjD0yQrfCjsLXiwVGr3saUlwvVecisOf4m7T3ApXOJ9TtEy3
9P2yXok5lgARjGZ9ec9QV16AR4MdA/9QDfxMcbOp/QMcwU5kvLGwAX1fkVQPpoyiMR715Ue+wnqN
CCQ9EIQIMW6/PeoEZBpv368A24cfHgPU8lbO51slEcD5KvurYdMG/oS0TGXHklJw/XwSJ1SoOvP/
I8Ez5DxEiXySoNYFe8H04wd+Ba2GJqFPegGDIePVQSyraOR2X8EobLANVJpKYH+PINAQGecHVwt9
YSCwRM+sRrUx4dkbSvowcfvJ7kwOd0lvB0MnNWwLvgO5PvWyj6zfRXS/6+tUfXaCRBoY4FzTG9E0
Fiavp8S1lBnLkLhsAXhswiDJ1UoSa5rADl+ma4T8AJUzHhd6Ey+h8DXGAnmyCEZ/UvnwKCpnKmZ2
hy4N9WlD8cCMIfnJlTq2qsTRBgDb83Vg8LKEITJ2LRyRJ0bWkqozUic762fVZr4IPOWhQlpMFK2X
pEd8MbxuFKPyJI/YXA2GxEeWFggNgxUx6K6FyR5KexJO/QcwyvBdSSvUd/rI7DWLN0Eiocjbcnr4
IJad/FIHKtxMVKk8gqY6hopiqsvmCVBScDUHrJK0NBLlv+5vcw1qwIGTe778kEF6PdDlVTUZUZzg
vyYd7QM/SYbIKb+WWrfkwasswicoau++6C4bWnlx9m0YJ+3RYqB4chLkUp9+TuopReozaW52Nnzv
Rf9n8tAoOH6gZ4nG81ackx29wgiB0IhPxtFb5gLVf/fQKSZdKvNAXwPARyaa6r0/ZFF4EZ83E50U
Q3ouHK3W5l6/Z9Etj5sYIftzBWNeokap6yQ5MEZKK4KEqZHa5LZVOcFMVqBCjYGBsZUUoigXMCfm
ry3CaQvlmPjfhpq3EnqkLkZF2KgkVZNBjenSQQwnxJRLH+rcwCLVa85+qHZWKOCtP3hxsy4fsi4L
AKSSbA2ggJqwLUDtHOouc4Y4E3SbCewIZo+O4d8OTpDle94b+FUYR1ZIw1DVaYwxNmKJhmQNAH+j
UEqEmN1g07PVVVM3wpRxBooosNALZtLTjT5nZ3OGwOccaPzc+FdGSlc66e9t2Pa6CtqTTvBJ2m6+
5usEzblx+SmJ7rxT6S428HvQBK+TjA3/gXrlFTHlidu6viQYnRitathH3wP7EdEdBov/qPaXnIx8
qNhsjkbZADHhuXqGoNv13RNOM9Nm5s4pIm4YC/sMoUg3f6OgkV0QYUcAKShqCrbBWbam4tTvV/hs
K99GMpoO3iA+8k+F8Bs4lsrRpzgMJKanYP/S/arI0xgzFAfoMorXtbmMCkJIC89d3r3jYJFrLe6r
E1hg97KI2vuPhxUP/aVLHfX0C93z4ZP8PfHGBFZ/kkfwaKSLyfaSEDuVvwW63iHPpcA7aFHb+CAu
xPIqKFgxB3pXXWWMlSRKXynO4i9jzF/DzixlTDVOp3P1ojk3qfPuiQem3idIlQJFQhO1WKoykVbd
O4/+Mus8E8DykgY1f+BsfG2sWGlnn+z3CyhFiIIs7YEU4xCg6JTDkvbygX+63pkFwGvZK1hgKRzB
iH/T/Lpo9qGBgYLSTM5z7dG2fptxP6dZTIBcKaGzodPzYa6QgwGwwHZF6ce0WIaBgQcMaH4MnbkG
02zZBCX7f9XK25DeccxcP0gmnigDO25RNyJVY4WA00NXbI0J9GisWoGlBKP4vRDPqT757zIobHnx
GYch4odu5so+jHf97y7HTQA1WnzBoLeVyOpcH0pSlNhQV/xT/jFk8xbfnbPImZ9rSjLklB2vpZpB
HEs9F3vk+SknRopurX8YdfkiJNq9bOYiWGqCP5dpTNH/VKlACxWSt6Iji4bjVO+iA0d0VDYTw9pY
uy0zHelRupMYr/PVNDClb4U3+umgKq8KjlLfhE91GfS3zCF16grc5V3Ms5I5DKalkT6OZe4Oumz9
iFY7S7cXzKsXtbC2d+qZKmzRp8E/sJwyY3oSsX4DJmHFKhz5w2s/Kp5yKLV5nIV2WiI7gNKL89EV
Cs2rFmUrvTPePmsw/dIEINUhBSWRRwpo9R7gXm9LrxrSCWxiVivBv7ePCurCMxQex0UMQnyLBNBe
f8QuLY5FKy5l3ganB1g1JIKAxKyJn3tQ87QyXY/A/cy9FnlwiS0VRdJVz2UuuM5wBdyZwsewixj8
ghEnf4AVpTc2+7ymfPSmPgOQ4kMvToM07Zt9yay1owFv2wNKO5XNkeq5rfKRb8DaiHIsIgcuYp6J
SWHS5vXluBx3aMoxPK+699QejbjwRm/7wp919/VBv/AXbzJkrYQ/n7FZfmqYVZZklzbRChRqxfEd
rHsKusr/qXOKWmhlyy0TWFCHB2t7MueXcAC3SNe65QOIO1GVHYDUOtwKezr6dbZOnR28qkH7fgeM
mHmjUduLjLG8Q0egW9SKpNuuoP3bebgVG+8yUEM25Wn3mlibvggJ8G/BiBjY3JCanPbC8SyMU6vC
MzY9txP7IHQU8BVBgU7c/AIxF0chHsWm35ph54hSUxPXsNmrz1jqBGTrIDB9HluTgDWGyxi+h9xp
Xb+t+kcNVQFjN4FQ8HmNRaw5DjPKr0jbzYps7tTZ6LAS23G5NHJw4i1ZxYDjaGz4fNOj9mo9mnIB
qE7IcpD/9QGv5LpdTVo/sp1P38OohizJAJuCxdjy2NoahiUIq/re3FnDZ6kzJ46Y3TLlfknQ3m9U
skWG8uJaIVN5zGa49K77bzSshgnPztvSOziFYKUSueOqUUW6wPvZfGLyJkRV00qXvXLfmRxOHbUy
cqqdkuKHV34Wx8H3zwepk2dTgDaz+qYukC6a5qSXWunOyVCuyIZfaZWuWHugSP26zQrV9uyVET5R
qawaCS8Ina3qF4+VhE3aSGNqTorsIC/Psz/fGYluKr+ULMia/EoNf34Ar3QoxFMqTvru//+AXhxA
UJmJ7SLx9tJwpSRJ9DQqOzSaLQsljyJbXAnuL51Phm8x75m0g5VjSpJleBvkHk01vpXAO8GRqw04
DJyTWjXzPrNKcF5oHzVhoyGZhZynNYeEJqRP7EyyrGfVSZjj3T7URiqMP/SQLzF5f7EQxBYAxv++
Xk/L1NJlZS2cLyFbRSrniY+odOQZm5h6xkF1xPxn4Lz3th8C5Onz12ng/w3k7AVAWRGFKGOnovdf
IZUKCqH79egTPu39t4B3tkYA04w2SWrbzlX7gslGNmxxXd/aVr2fby0cwEQcb38jtyylXmr4XMPK
0pC9j/0yRZbBL6TWoAMbzM3DQ9CxJ0iEHNWSYb+pCi1D34aQAdKSwkV55XlR89XAiPp3jpD3l8ay
Svvly6YmtpF+mY4mRRN+serNc4RDQ77d6KyWC2/+oFmLVgiYaMt55aLl/3Owe2AI5T1DTefgesQY
dGdWJRo0k9dCjjVFscEbtVF/BUlky14ufWLfjp7PPVjzvbYzZDOa9qQlAHH5TauvefVy/p0c6NcG
tNg4zOEUkCKSGSt/RQ2A9LCxxip1x7m2m9nlP2jrde8zwLI+ppQXnK/8NB8zhXrCp1UYzCZV2s5J
jU+qInczfxDu6Alk6jmGDn5cMSMsZ58uEVgnW19govgGoaimV0Kbl/i3rcUlVvLaYricwnhDrBbV
x0CoRM1uN/kMhugJNeHX4xOjHup3QvPFsFee4OI7haLeRrnbXYFMwX8cMKslkXFzexC9TbabNw0u
S/zAwqUVDIIr62eLqi//lNj/hIMl+0ZSGJ4Ssea1BNCE/A0fyL3VI0ON5rja4vKEl1qXL+ehuFUR
bWxhyn8EgS9vlbZAbFB+LRzp6tUPJXPaFZpW5D/N50X1E56ivoevvAULUbl6D0nq07/eSKH833oF
S9rzfjbJ0fRdW+y1Mtfs0XvBp0+tKsAXPDUwJyTl054venjIvkKfWV4ahoYRw7iX1Jg5AtLiHx4K
MtDlsswZxM+SSj+gPTdcCFhF5vWridOjd9dte8Oy9A+upSK1gt1dSJsZwOji7c7aRBe2u4wnmJV/
AFCRr+HTQTjP/5Fpi5dPKkO51bINgZA1gWqzvo+uGpTshaF7kiQXmC9XG2Ys+FHNV9IyO9PJG/AG
WUtk3/WLudakJtieZh4pIrP0DhIKf86a1jThqd+wSeIl0kG/vHeq/tyc7Rpj6Kt0ArnPzvHDeRj6
Ul1Kzku1vrup96Ub7HpONzWrNtzC/3KO4f1r4WwgWd9fhA5aQmWqQkCjTERKQrtjPA4yZDS8pg3J
k9DzWtynJPAAYkN9pYA+9HR0EITJV5pavcR4U8zqPFUB1nKXDye+Ruw+5vt5VoV6JTuuA+9rO6KQ
nVI0jFlW5zkpLpbybvYgkSw4bFjy6IeV1kNZuPbOMolod6hxWx3C20Cpzg8gMLPcJGXCLebyW/6l
6EQf4o7tLPRywlWxJWqv/EA5+rxgBzt5zC4ik+3ctvV83NxUS+VXVmiqul1L6ky/E3dfRIZWyy7B
iuHOzBox9sUe0Yxo8HIugZ5rg5UMIH563a5J+wR2e2b/QbdjOB0eaN5qLhfjjfFFgM18BBtL79ED
5s7rSnPCMn0bXP94lMy1+1N3U+oc9TBf8XEJbjArqjzXNhBizVPw4vY4c2/yBcvPGhYi5Rj8dGhv
ccYxwtJerqlJGx4Sv4A4A2v1WPzSH3poiZ7riogTyZm3nnY47hlZXRxmTLON+jwj7WUoA2RQTPgW
NQ9/FscY/wtq2viK9Ied7oEuWQwfWg5IFeM7cO+N5GEX7ngmU8S+/LqDA9ccaQrBHc765MHsnBOC
Vk2srHSr/QeQqpQwx0ixJTM7qbLOkO8kMDZPkAdWews22eNn5SpOXGWKKmM1C6spim1XVNj0gKhv
aqjuqLczeVNhLjbmd6ii76Psu1buk0qEl8B9ocXtHnPRm28TtIXtwcVO6QO39g15Y+Bmtkg49dIw
Qn+TdubQlB/DYhljDLLTiJmnAXzMWWkyxsLuMzQvl1xCOL7xSXd05ohsoFmcZ0gMtkki/zHQvDgR
1NMZ/AQtl3IQNlWLQ4uD+Cx83YGS83QjaL+7sNkWraLrtXMBvNdY3v+545lOZKkEo1t4tKHL3Qj0
ukE9uV6SSAV74YxrHGHPjrEKbVt86HzG8+bDfAmM1vqnBOotdbaLWHabRgsoHHfbmtexz8GJB/bu
Rf7KUCXPvtNXfe00t2B5JdJjpAZJxOyH2qbuqtaCCc2gj/DViidJwNWroofS8sJUVx4VSQHQDADX
1nLVxm84aK9Rtj7Agq18SMY5DvZOpS9+jNrg38BeNwd1PUE+OIGmbnqtig5Z97iLD8plmThUMzgK
gX79Egw5nu8iBu1kEL5O1NzVxuU4/9zptKjjFKt5JaDCgW7p5e7PGl/xOz8eNUuHePTFiSHIuQeK
DN1P7XkqrvYwzk6VSM1i0cbIeqT8Kr9PlYL7Xde7RoHkipTIsD6b2DoNGJYHh9g4MnsXMG3+kp/G
dqUjUeHLA7vsKOx5l0vZ9oNWdfuMLCEc+uv/VLyOluqKFygTnBuRxTgEFGDVF9SH+GJVA3wR51Lx
onhhHbLRNbcyeRJp1NjufXJbAiGAmuIkLHMsymViqisPeChBW5GBiI8IeczFBmG9pjF8J+gmCpom
oyLH7Y7tTNB2FAEKvs4troNAVBTzqoNpaei0rWJy/HjM/1X1izFsUQX8ymqZjCr8mhlPRH/qESev
CLVRAWHjOuRlzRcY9OwILdOwvNl4y3az4Pq4R3KFp64lEahvmpqyZ9ot+U/cq7z4jmC7VcrO0dTa
urLU/d06dr+33JPdPr9MeQ6yhqR8Um2ibpgHwesa7j44P7jVKKB6kheYKuaamyFDCET7L4Qtx/wG
fWIZuwfKGYaZc2MMmkaeb412kEXDUKYIVT2OUWD+Jb8qZNSf8GFzHYbRE8e16IDNJlo6SI7lsSu6
2BoYdSh+J6J3mjyK5Avc98+F66IKxHYCa/KPuzbz7BLADqkgZjp1rOQNk0XFh6GrYp3NvZEe+OaR
JE+2SmJkAfvzzWzmufyhGaAqeibKPgf3TfnZvrbm8IgS9iyxVM4FORdyNHqeGukwn7Y7jQuV6R5T
Ueqynp/lnn0/tLbGYtK6RW0+L1PQVtL6EoA0uO8e3ftSle8z4PPY2BBcL6F9CamY3N+E6pmoUwDy
tOMnnbHjJwEv/49hzlfLsGMwy3MWzeqeiH4w2EyPzV/BtNfWgfm1xRbILLYaC2TIFxY0utAG+L+G
J6I0unEQf5v/+3xRM0N4HCcvhPFnPISzXERnNw7SSu/BNQ/FmVZwdwU5beyQz5UmRhQKp2r7BKyY
9MPO0M/B9LgWqqcjxsKMrXoREDjLzJJOgvbMwSF663w7n/mlFE/400tfIjj9RMh4+x2N26snPjCI
q8F/VT30dGKqduOZWxfFLWtGR/13EdTWZuJiE/ugLE97kVX+YHINWrcDV2YvsiAr80wWHWZOKDm+
fNRDrJn7yiDRd9zZE7ZqWMCvrRTvquAlbMXLDbjhNjBKV3v8yRxGNlPAOyAulTS43c4+bIwo4N9R
/YGBmoyjg+QfpPejmASpmxjlEsbXCxxU3Nh1iN4MD55+rwJnXvSjrm5F4d54necy2H9q+qvzQ1L6
7E+/u1YIVBOsc/U4G0aiQ6sMVZmFiu4XoFI8jUkR9gM3Y4Oa4bqU5pFOc+y6bX2TNt4ZfHP4zj5j
B7wH9nCL7AP1zeJid1bQV2szCldy/QOIf+tvpIZ8THCLr3w4IAKCbWkWxs3ZtzEbSnkqyx0lIjW+
QmQ+daEQbFLTvDeqffmZYoqLQ2NBM+DulEG9fqXTl6PYceFV3dZOy0e5xaWWKbyXiFIbyN9RtP5D
ImO0PkXx8IONtanczii4Gc0ta7hP+t8zZ8U2RvUyxl9QzCGIEbZn52RC0I5OEy9p63FDYET0XZAo
Z5pvGNzvnPMFROwHR1WYKoDBb5uOnj/keAruVT5HdLkuTDfoML+K8X87yDkbjg6o6qnypQwDiZpI
ObZtOx3lrtcfoqTJ1EZ8RNE03CqPWeMs3QzUGYRxzWzj8bgcMFK8qhvkeraWWYPu+UUUELImz4Ms
3MfUf7KMelvWmau/HgaVRCPKJC+uaf0IqNERUYpTxTXXhjXhCElUNDekgHYkjAS3wro+y/lQMu25
QKFLcl8+hKcSuyMEg69R8jw9CarM7jgC6q0gnqjV8SL9PJSmd+DyigWbv5bTziYCDTz+e4lltA4s
HYWS1fLEiDOBoF4VCAV5lwyRlUL5JKz1H8RwZDEV30SSMPgzHbXkLqwqhQQLZ6qJYtDrVurTtB79
xWdhDex+Np3ia2tGIyVH9U+Vx/z5RzEt7coyeUj6PE6NnNcswXSbqa4ShbZQ1TiaT05QVm9P20to
B9DOT0R/J39a2KJPOYSoPofIBJw1+pLCXxpqoREheEPNxENz8GZ/BwY3uyX+ADIwvQKMgNsSx0Ra
wVk+D1yHbrh8T4DLd4OiWpx01GW90gGvKLGivSX//y5XdRZcb6ORZxQETDJgSQtVv0yCIt7OD/We
NyV1RbsBC/URGACrsm7GR9u245DKZ1MsqvQwAppCtNhl1+VNye1WDkDUU7zumgwxqF+YdXvnePP2
mxF3kGJolvFQs2rF/dDezUy9EiToPax3cOwpAEcVBHAhAOPV+eSF/IooLhxf6QtKKdxNKDjcR11r
rnEbruuFc6Q8WiDtIrkcxc4U/S/m3+iBrRNjU3OtagBTY5KAnR2T6A2wKuGCAoWTeHQQC5Hkz8Lt
zhwA89AsbyVl+PeU6KjDU0SO6KnKeczLsJgNich42+icYI8tRX4tbS7vav7nL+/9iTJzHTyOxYIO
ZmNschFevapXU8B0kkEbFi7mBg/R51FGgmsYGx5eL8u/Xz9A+lpmL/lvYChCyQeotW8F979mwTix
LCuOUfnh1Dj18i0endTCzRABpSKmsg3+YHqO4msdW+UhifR+Zr1PjJBoGuP1vatvO9CpFyXHRfhB
Iy+P+VxjtB3afBs2pgK1hhBCq3P6bTztCQ73yKLp9i65jw1rMq6JL2OTR+dfkbDo9J3pyRd9/cXx
pa5L0oGXZCiq5KfWm2+ov39vM6rKTBJWLvc5DHEOMjoZtVN2nj1xUrsmrKpcGZxld7c4NRFuNqvH
DJl/Uplc8Jr41rnxc87EEF39TBwD9Fi1F8b54WMyQ5ZXbBLpy+3OmcMn5SJ8p3Men87vjlcdtd99
UzKhvRDAEJSglTT3FGp3zenhoo+QsG4ZGr0dwArErZt+ToBy2KgcNWyFBd1OG2cCa3A4tlAUbfp8
lxRr2PDmScZLtJZBmlBpL6u05iTfIACNeN+vY3X78HC2cvKnQ6Pvwwyu+yn1gU+/VH25YMCBTX+H
45LTD4Af8gF65M+tp/KGEdhLc2VaKPg+EH8II1QqunC0cUHDyzWZx+A3mK6P1OXOWHvzKbEL3WQF
qFrMRA6ff+KJ1yQXl/7fL5g/jPxt1luIiR+CcVlFlDgquywLwlK7iJh6UA3dqyLjoG1QoL8KHZY9
rPlUbCavqGRRYTLI2PjjG40A2rUlh46Z+qjEs2YzRWag7F9FsLX+V9wBc+K9i6YhLL7yDBtWqUk7
AhB0bLgtHl3bHa7Mz6ub6k2XgSazQfcmJdR1Fek4cGXrdXOfxpDIutnjUIFiriONMt5RsB+fs6HK
RKwbI1XU6UTFyZUrnGQlpIE3DgIzzhANN/6D+Z/VMpMZs9DxgmuQoyyQL819T2D8I49cqm7Cr6UY
p+Mt2LIjSwFoX5rKQ3vB+2BXTLOaQ6o1bTZz4JQbdNn1cOiKWKdh4XUUvexD64rycxcniQwuwd1B
sSTeKfhoZDhC1KH1jTb0StAjycEIC+6qIxkUaiOtZp3u2FKStNFrYexnIvgRhJGRMbF9TO0S/oKh
KtT88k1plSFQFWtjx7+SAVxGrnv9uCnwkNwBImo1LlrvKZJeJyaixyM0MaKwbvIo4vfuuvOma0WS
NT4SyWqmR195y7oDWnBcwSJjXYniC9YlJaWi4LpWDWtx5xSWq7CX0y0Rj7wCox8n6J9Kcql4UBmO
X/h2JVAwnI7ktyD1CZ3ouvgftEme09eyDEoVkNr5sS9PhLpzfd4EQ8Cf4gRUadcftCRyYZ20RAUO
No5UmixK08X+AJJtqHjBFgSnycZXlcub1S8komRnV7++Ci7B3ljnQNqljhucuvDiYR8dI4etTOkq
Kl6qdw8h0US6dq1I1vd7rmA1+YdQ4cHqOAn5zD/SaKVLKpHYe8di/n6ZdhVKU38tbvXvbV4Q6Fcg
3RmSMjO4Ste2VlJ4kSx2jgIxCb18JmaUyR2jua+5mG8BgTQFzt+whiXHJjXMZSwdKYV+dnO/3Qhw
b8mLNgzw+ZDv72Xpe3J4mdy8Ra8mITMvHVlf1rd2CCWSiWWTqHQTpRUPpCDfZdzMqxgYOwVUXFSx
3wfvcJ5xWhq2/oiJ8d73TxRcUqw9SOa2XA0hMLOB9gUMTcr5sxccmGiqrYNRgtXCMGmogsdkH0ID
P1avy+4yskOvOJXS8Oh2RWaivPaVyywRgg8HayQSqj654+Je/CvOWigUswtb+Z6oVUYtyBtwPhz+
T8h5l+DCAdYy4ed//hK3U5xPzSWj4qXchRwDBaX3Vw5z/9xr4yPj7bsKapLiPA5DgMu3hTQG+n3V
eK5Xo/hV3Ujy16vQxPsgZSncHuqw9+dz8nmEqllfTKZIrBIyNRAdSH0Jz+jhi5F22fquNHUdaiw2
2jg8bbaBw6/1W+94+K93fWmo+wQ8sAwXpsiFI6dgohjqFhd2nlYw/eaPDprqPd54i+9cfoBkAO99
IlsQF2DXzWG9waahAA1xs0dTdZ54YRN4xLM/Qxg8OxYHwG+/S2ntuBJWp3NGI+W8DGJUHK6NgkS1
HfFURYWlQDxnwhbEGxn3smQUgh1SMrFEUDvhvoGikP6LjoFhX3AFRmO32+L/yuHTMlApN6Qsh+M7
VojxZJFxm3AGdZBoEx8OL92uzP+jZDYmnd5KyRadzcnS/Lv0bpvUdsXUL7NdLJ0oRv9tN6bmdgCz
U7QzavESyvgggbkWKTMVzkWo3PQBowVfHrXZHlQTlLa+ydSqme+j4xYEM9P4NWRUbAWdMnjb0JXG
usMbT9jPuo9p1utX6mWr9fEVjRChmRKLq42rZ3jCQuvDpNwfWGfIrm/FTuPwoP3ZWjesnNhy5PHh
PwoEV34kY/jJnZPyFz0uLpTmYzUZ5Cb1mEG9Yh2fXXA+haE/+XI6SCb+jiG+ZwMbZYa+KjRQ5uwk
t7UzDAqz8+ugeo9wwiHbxiFu/L4GdBVk9IE8KPLbYf22y2+Ta86arOHnfQ0kk146VqbSLPrs6VNB
w6Ssgq39cZ0WX6ij2Lmjwx4wCKL27Z4dc8nOsAn7kDba9EhvYh8uMcTF97949vHo7cZqW4TOxGh0
/gyzCsHgE3QxtJ0tre8lLx8YoD5m15zFZltBKrrbERnusuOCdNsoRtJqnio+N1L9rmK0TljkJFPP
32Dw+PHMRbEddCzRnFYDAvhPZjmSi+SDTogaylzRJa+VDqG4be7whe4Hs2zVEA7WpRULWWOWE1BF
Z8ULN47Eyono9vlT4a0D6+L5s/zbKi1UyoLCgqBTtrIPKLX2tou+Kqf4h5ZgX+nZ0eWCcQnafoQR
gEOxDZLlfVOSj+1u2xx23E4Pd6V6txxqDe44RqMBK4Q26bwE35TtTHxAwDbbKAycqpMKgxgcWB94
4yRjjBltMkelTpPq4BWexPONXVn6DncwqFeInm/Oy3RsZNJnpuqgrN+3/fCmGAYQoFmOXOYfTPZm
NRMBS4VsnFK71F5dcGomYkYRKgp7sgCIOJu8roh+djwVmZIJKcBTbZ8HS62/rJqAN7A2v254Foij
j6iS/4l9QYE1EdORab54IHr+I59frvQyIAc4fqm/ZkryKYb2ZjAW5fWqKTY/MubkRvEm8u1ncp1Y
TG+ieWgKGehVu84BtEC3npyuqQA63Ud6R3+ofdvGWC8PckDsTii2qcRZbbwzKIz8lcsmAL5Hy3To
k0PscLIX/sE5fDMi7gL1vMXUQGQ+cse0DdXXoG0WVpp/l9ERS3UDhE6kq2ZKfKGTwIdoUdc0L7zR
9Y3d3mvVO3c//IDwEdYNd7o6dH36DC1x4tnvTZQ1HFd1m70d5p7OZGyw5V5Pn+On4PiA/BQsM9DO
hwNdzDrHWbs2cd7ph6oMWC7zBBJfN+D1gteDFStnHZi2CEddMQ9e6WJNPcLbAV0CD6c2NLScLrrR
ZjU53MDNSoSzpmtXKXUX5hzQ4fiyb3DTpMxdVJfYdMEP1vY06qM7hAYNYWu15NocOLiv5yYFZF8e
38PCpIQT2I1kRJMXTLs492f5xydKmHnZT8zRNN8FGLVdnyDR5/PnKAK/asJp0x9nQomFVYImYjS4
YkPH/5jNPWcdMiRBYoscQixbsy9jzdv2RV0gMhYJ/WRachyAY+MinFfV+UtMIfU5xazcfDyzriKD
IEnhMQuYpnX+pqDddqiD2uFpyEhd9YGww7Hf2o6xNWzfdvgd/1mkYTVLY5zvatfnsHFWyp324Rvq
1Kas3uzUvYHoMRmFhEbf6wJTVDIdJVIXVDSDjmpLpJy9yX4s3e7beisFmDUCAi8TsO2VF/yVBIpa
3QVh0M7V/WGr+vlufzEiA/oraABqtFOjg/Ck7IU9KwVZhnoDoCVDRMfuR+kpFtOijNKH5Z+su6gs
NNAUSTiDRbd9n9BLpX/g37Dkg8GpanoRgvFnHHp83kFuDkFZmXF2+NJdV+1dCQND9A6mNZ64s6NX
6ALS1BAYHuMdqF6HVKw1NS9qXK1JYUljhL9b7N5Oxo5VNKMM0ySpcV1R8aPiFYWsLMJ1vQwj52qc
XpwjIO7nzemOdzCNzcPBnGOSKGfEVg9tpAT+dHASeyffa+bT4FFxjdkrKwdfhxtVBHoeIPTb5497
JDnb1znxV4HXv2WFU+mfJw9kQx/PMcfTnKc+iuF0jpm9lTuRBbp+6NfErVmGE0oTFiEaRQ6t2Ey5
7vkoKLsI8RXrLK+hCY6EkA400ex14fvVHwT+se4852QlxmVKotJW/bmqdHZSqObGZJuJVMkAfjzO
RGbRKWwlq2qnJ/ZkdU+KdZGA8y2xTqyXTk0RhFjVIehEsN2iNNAC4CljLSPhkX3KwW6ZioltjDPt
G2VxFWtW+nlHugGSJUbvCSuNMZOhzjB2X3PlE55UG8Ye+VTJE8DsJHE+4HTLMHu8pg3OizS4M6Ei
PuMLpy2ttBUTvqlIp1IM1yMwOV80T8DgN0eX075Ra1wV6GdFnaEGsQjJg/uudzbTiehP1H+VMJ5d
hSe1nqS9vEboFfRJORez81SXzL+iCM++n4pJbXRuRFPo1w5ITu1u9qWAlomCO1nxuQL8qp6K+snO
wJP57upaMuf+qDlQGnyEPQMegSDNIV7QLNKYideAMzyQ+VpkKMXMP5yo7NixN3sDcwGYOIsbUDds
rOS4yy6ivDaCVSIBTMWe6Qf1hw+v8F3pZlvINEk5ztVwrKxrRiI5FLGKrYuA4TdEHaa72ar6LSIf
+gudvhLgvcvWcULjtK7jJuuAQC/axHQN+Grnu6qK66TADJ96ADXnHDmCbbw4jLchQtGT99EZvJaq
p53/S+rgghwF6GLP66W8obc8B2rXWMOtITPPfIHY6c+V2JGzJoxMKUuBH1hE1Yevp46ggrbSKVLo
ft6gOfDP1/y/YlJEZ1e1kni/HYt18XJv7aQwpPSYlvjhwB0/0yRTCMU712bNdM2lpxbNNLT3ev6m
6ou2EfV9bTbPy0l2n6yG/fvlOkWG+51A8NJ1bltQ2GZnW8S02XaCguW7Y5sbCMm+zb8PMo4Zt72k
xbY7xS+40FAEKNEsW3jGdmcdjYBiNlEheeZ2qup3O+JnExVZ99Ddol5AVQYIaMrsoHkDC+ahhBNp
QlrHi4U9/+tlaXblNZ4hgHnAerlztT7gf8DD7FhffnqSgsUqTarXNhuQ58fxb/gYqToGdfQ34O3A
lGR1ONfm/Pwl8levu3zKsCGsisGqH3Mdl25gR0gEmEisk15wHasWqkaFcLi5SkELZd/sOIw48z9T
x+qt6fgWEnzyRUKpnwm7V1iSle5I+8uWtCeN1w93TFJ7NLZxeJ1mI1AHtzQhpaChbqNqf9tnPT6w
4za9r1nxBJRitQOaEH5ugP0oxuchgX0IxCaw9tAgg9uJwJ+gFa9vfUWyz8rEvkD1XUvafmdSdJg+
zUbxoMCRkn1yP2DIz7wCIvIgiFunhjL95wHA/Su7iSpk3YsTNHjbbg1DbSALsC9y7FQZyZkV/5LF
KUkNhimwkZwx8y+B/Um3CuC6dvKnTlZeiGXrCxxHJAHKnRnJRakgiwIOY0lGTKyaheMlfaCKeddi
3HakCDtB1r30aJ8rne3aSrXSCdK4gt/OHUx0HczlepMUN1aC7eKY3WG/MxgC0SX3bJXlAv/RJCYx
TCYd/fnyihYAjHzggVnjD+NFlLpT9a0y4Z7EZQwCFMSIiq55Ejoap0pgNu/+YfTrnX9ZJl6jDuNt
vHH7OpdlaPe5UvclM46s+h89C9IcUV844NqIyP/1aH3p0lYt8xIpp5u9d1ntLXmtJ8K/YnrQ8DRl
fhEqjYZaTeBsKhItNwNc+5sSf6z9ISz2eOjTWrmTkpORChBeMEJkXmMesZ/pvfr5bJBvonrFXXlF
YvXDgLIPI9kwmokHYk8nekk21DMie8hjMYZLnVzp9ojO4zf6iUTGuSImmFeUzCZDY/VIa7WZOByW
IjUnipF5kvIw/aoQs3mq6R8FO8rzbxn3hUndSCfdAQbBiw2m4qauNwmuoDf94aziTbEDrsGu84Vc
rJnEfTaSZ8C+00EkryPOkWEn+b7yW4aLr9OEsFw3k3C0IwG7JySlbKFPo00/1JvSaNQYcRsoIYNL
I/dwnplmael0GxurdVyGvD4TiueQrP/Jnel2O4nV5PFAI86vvG2O+yPF1wRCgzIjJegA6EPMoUEx
egIR6xl0mVDV6Z+2/16ihlvLm2Q4IsgxWF/RK9baCoguVaFT52SRFRdhFDmRJ9HTtXhau6q+wBbn
zMKJjhDm2BvBHswm3ulnrVjQG9vpD/n9zJaCa8+ozuEpZOHvj4kAz88LFHn8HT0/mhGtUvs5tBSi
rPS+CQz297aNZtYQSE+wYQhMWQ54mfcIVrk8Q/3XmlYuCpxqODV+YrkdX0qtzJotuBAyXgrvYGHN
+wRJuRFJxr0ERSx8QdDeL8p0mvGd+MDnPAJhxonfg2uJ6WOkSSAcCyacurmuTAzexAag5Kwt5mBn
3j+LTyphK7XX+MHqNQ9kyvFmhwP5sNkb7zjOLBFlDz9uiWj43mKrD53kfQT7NfiDeG2JnQ6VusOd
4ZjEm/fzJayXV+b+AbwVHG6oeWWRSYlJTpS08cSLZBmnjtNWaH/BOAAtsboFzLSlfxyFt9+U0yAf
zlWk8mpLRLr6LwmYbI+4zoHy51Gwrlm4/6jUPg1OvbgrpRxCgwldI+Z8A2bwpeagGBiRdFf81y4w
r5plpYuMYFufPKHJb5sB/YTZbmUYeLZ3utiC45k+4dRmuRZe6LdyXo03nmb/hOOzPn2NO9RV07ed
tspOnyv0beBJWpwKrdMiXthI7K0Lqijx2H4GXTVw8VLkwbzSIGBdiZLBAemw/3OMOa6CU+Aq8JVY
rExf7/SQ3cduho/UZMQRW9wQZW2PdARbHZiYbiicBwVvKfCI5sNPtByt4ihwBkD8xdDmJlP0Jm1Q
WPkgddDMBjWH5kZUtnf95ZyTGPnvfLSe4tA3r/pvk/3eOdi/ju8e1ANjYbMoG8Kb1HgiQ2t/AiVc
U3ELy0vjPWXBHZ3yNzdOwiZMwAtfBQ4aWZtteFZiPFDPVxUr5Q/PZYRhDCnodevvbnnQxx8dgm+E
pt5plQtuuCJ6NkpVQfcXHsCu1dNO76xqSCGG9KKnpj+ByZK8C7Ijk4xAH7D5P2a/cEJil5sIu5NB
N+nBM/TCBtUvwDOiLbJUy1p2mPHSzsblkUYTfW6TBJXW7Mm7a4gEJKUc5dsc4KwyXXM/ENsRA/I4
bESemBX5MP3Gymkmnj0o1vYciBUs96pYoQZpcC3OGNjpxygP/4WR9cxJaElYtoefi2h8v4E4pHpA
J7XtryoVSajxBbOd+rS/DAqqy8lpjMCka3geo0IyTz1J6gptqkIeJYy94aS+tNBd2FPvvG6e+l93
CFuOXpOdoySkkFvD9qkT3P8bDVSMm9Ww9Tve5RxXaOylVq0joJwL7KNdyEpbaHqHo/8hn3om88bE
6WqTsHkRWQdNGHIUpU/VQf+iyKthCsZYAD+iChS1no+vwaFu7sxc8n0IJXmQrR0gW8SyWzDijUBF
8uAZzyADlz3kp3Oh92D7mRlfy7FBATrgfodt13wc/4JFMNHk2oIk2TG7U1QLciXtPWOu3VHgU4QT
O4AJ7eVMxTBnEOZbQlgSTKo57m4Yu+n79Dcqv2u9vIfxIv6FraoHCuO/XnbmvlZAtkJ8t7SgPHYf
eA8hPuMY7lRCkliKvYsjy+QhdLPI/OQlvZjqVgvrKvAeyf76OJuUWLZiYAchYxhzA3avNaOeoTGc
7fopwBHH5vo9Li0NWKQZ49hWcS0ucXORMO8K7tNLvvcBKfY8uWQwyoRyf/1L4c50zE+jHfMSaP0C
ip8MPD9Cn5NXbXThOHsVVSCwCieBELitrzRRwPxGDJyHoj90GdQHeG+NH1V3wSLeWAsF5kTf8n9t
h8cnF0lkEF/+25Bj7c4Ktalo49E+0kv75gfOZiG3M5e9Hxzf2/FNirT+iXOcESFUJWoKmjYI5P5M
sjBRLUuKcn4P27uHw5mLGbSYY2f3te3tf9RtcVT4liasXGgucteEl7q676SdUC8VVT/A/m/PatQs
t2UwvwbJ95UTj5Ecu6eTUlzOf1bs3qErpGzHeuxW1jrpHtBZ0pi9WWR1qy3c3KwDBC75ZopsYbq6
Loh0xr/RqVAqcxMw0wnycACt3ujlgVKwtbpKU6P6IT/U92GJ6i1vGq+XwZNTN6hduBQKjgEJYggb
D++86ib+V1slKD/EWMHqhQk2FaSB2x+kLUV3XUuxGLlPABB7PB1AM05XK3ykhDJLM8kgT8sKXjri
fgrJemga90Utx061d5cD8C9wbP+ExFr4xVwI2+0XGtVTDGHoIsPizhQdg7KkejSoSkIhCMdp9eNY
uOlJSmmq5AgksptC3lTKT7MP+21jce7Mw9R1e/zH8PaVB+t4qJNpAscPBUpIGFaLWnIphYTDI8VX
rgv6YsCm5eEvi3npkwvAcsO6utpOAfYmCQwCdLPqBn2VRKwu28IXvwbPWUpNFT90bzw+RYrjSksu
KhuCNez89cALaNVHNuSCeGoY4jI61eMxogKoYl00t1lPfbru7/9wmIfilK76wb0hWQD8BEhlrusa
9Qnp2nDzIYnHVeCgdWpjEh+Lhk7gC5AateMTDCaFJ35yS4PlwOt4r80Kfu9BUVRc9Sl6V8jtHThN
QUErM7GYBJbSMz9CvHkumKdSWLQmAUyX1CGxpXcbSthR80bYjYsE4ZwZmwkm3/ZMOtJF9DhOhJz6
aZIX0mRj7qgAo4EPsaBzI5P32zhCNB5Y1DVlAne4UET/5q9oGnUVSI3cfz586B/w7mHOOZTrrjg4
KqKYGy59Jc8k4EPwFke351kmtVXCDGRB6+2GBJLKAI9vZlBMuoVnKPdR3xlg3niNie2YVIZhaWeE
ERAx8nsGYccAxWf8Je5Oz+rd0cPSF5EOyzqPWOMacWacNocwEPf8RR399VuBCR5/UDjHucX37yo7
wUl7R6RK/1qKSfe8HFr4oHwyELtCKYcDX/BK+o+c0b17uLKb2g1+P9u6CdzKQEG36xb/wipUfbcn
eRTjYwGg/sGcp7VKHuBP8NdU/Elxxp1JXsIBb9OLHRYrCQuD7O7sLR8DYJwsHew7wT+5EmtK4ulo
pAS/i3aRjtYn+KI72vJiG2q8sJQDYCK6CVZY7aWcwTibhWTJDQC863zt56kyMsu1CtP5I4HR/xMn
fOvztH03Z4s1mWcymDtZuxBcVy2vj71w/BYVdh4Ox+zOXDyU4Z/sXhMb2A+XrBUcCSGmFqa2I4LJ
CLh7BvuSl3P0rEJMyDZao9/Ai/A9mFUYMcA6e2KwiW1PBeo//vJ7FA2znLTbojcr3U6CDYgjBuDI
akQ/czvvqeZvzpNl5Hq8eGjKodj8ZVGo2rdyJ4OHbS/2Br3+AxDw3GHdAQMuuAEHsdXwPxc0sPdZ
Q0TZ3zH/ThQ/EI65iVHB6QbJYQhObTb0MuVg5DebrbdbjXXhXlG0GslR4Bbu5J/OK3Iovl0p/U62
0gF2YD4WvhRdEaAonWIrKn6TRSPp9dAMhxtwx9YWHIHbD2oIyWcaiiuOxJJo8kvL6lHANTF1W3PL
LY4Albod9M2jONUrndtrKJCL1W3h1g0+umcUVnmxaHba5+AgU8AZ+UKwDHyEx/YO1p96gMGjKHb9
v5hw/So6SeMb9HtPjUDN/o1SbAqXMXQE0B+zCR4sS6SC2Q/SW6EW9uMyXv9rbHm5H1vIoVHVVKMv
KMBBifmiJ8yQNsoPEuei59KtIQAtju+VD3w4YxCMEfodWm/JtCWru2toValzZzsiNNtJd0Og23DU
xWzafPQ5jAvWa0bcEgpWke5s5jP+TCNiqqJ67yWc26edClaRCAghxCTVFM5jzsg/MH02OAAYuf/I
doKciCJu9FncEitq9gHqM41Mok5LU0qm1egEsIGcC8dSZtuTf9zSdTA/gJf0vD9X218rdkE4KZTh
H9RqbqpF5l9sRYnMyaMdulJc3ECqaDfYg6MmkPHRMwGA66d87j8bYpGWxJTuRakigwt42GOF0T90
Lxk6z0XnI1x0P/aPIt+1gDrMTHjeD+71n2us5ifnrTKzV5CDbFtWm2+Jx5tp79WqpXOt3vNCYnLx
LlpfgZA1JVC1omc6fPzlZRcLcvIDx2EtFqu2iea/qwVOPw/HwCZTidBFF9t9MJqlJDcQANXweVUI
9nQxm5sMuMCqd7GdbKDTlO872V1lLXjMLk7C7yytuKNDVEIU6m4qdEifHgFGnRggRsCxcTaJLGbs
PhmZJqfPSi3jKkknxyFOu+4LUXMRrYxMr0qmJFzFRmva/AJAg9qoS4KrOWUBpKv6Tq1WLw46ruLw
Ep1FFh4hk1pnQFncnj+J/K+4r3rfCeVOa3LgsznYnMSiSW//6DNQa869JCymebggXmo1QZF9byl+
4jWDOPePjLgGYTAn1O5+OvqLwKo9mlWG9g0Ze7HamJ0g3bJouPqp9iuMOmn7VVWXCMBW5fWz6+oq
/s8Ww5Ewu9JlPcw9g4cUCfBjj59YvMuYAnDwuOITYFgqbnwt2JZimIcK4XOzF+R5KzMlak8EkmSa
wLStoAAW6UWG2tr8OmYFpD4ARXEOmnt8/yF+zyPxt4g+z8Fvjc5XRtknNDys+nGOa4RyNMIgkGVm
rZCFjZuqFg0lAs0tVrYMuT3B7ZoEyvVtATNPmc6EzqGXuEuutNLQ3dqDCc1gnNYugkkOrYFz6Izd
ypyPSX83bVdwzUwGr+b0QnCMGv7svGkFjoxp9fL+PyNTBRYQ2mrpX9rCe/Rl25+WvONAiPdWdt8V
aS01d5Q0HqKi+/AhDUpATj+3Ikbd7ig8k7OGdBzg1q/3YfTjsVsT0Hc0CcZJpvD5sS1neYZad+VE
44GXtHaKlzFfOBc28FO4BNEQxnxlNKPXEHZ9oXZB0pi0mw/u/5RliDxv8sUjfh0iVDI/CeUYc8js
gRqmlO1SttARjkgbMKs7hCTocCG74ki+9iC8RrWlQ08K7Vafe9Dc1NLjSesDfy8rea3SIkuZ3n+s
Kj9VWei7MXLWNZlxovouGlGrdkTgNnVZihR+dyjD8qG+b4qNq2CDa8mZQhnLVrgj6vloVg/eNnOm
RH5T4uD/TXEyjQ4ix1Z/0RQf3ev80/f7gdy0LSvBt2Orci6Z55HiM3sWbneC+skZ3YaEWM42edC5
kFFJUnXPkPH/w1iiabYzB2o+qIg4VBQfoN9avJ/h6Ds8RGAWO0DuFI0qDE1Qr2vntRQYYTwK38u5
IzzXSIdgzW3zoO91X2Oa+g9ApqenLZBws54th/W1GjCJnd+6sAQD4YWcI0d4OnVZmQtlKHs+5HyB
2nvNKmEfFZMdrN5qfif1edEdE97hVRS9JjJf81hl0pSqbEOFwvmdRLM+vJ0+rsyZI7C5aadlXos5
NaUbXF9v7hKBQeD33sDkv4PtRHSwBmJ6KW0ZKLkTEKEQdHoDP6gXvceCzCF60i6D5c7IcuHhu90o
bI9SWH1fcjeZSxL5ek4lG2lXHEdhx1YOqLOuaxJE+rDs5GosGOj31gkAiSb1yy39t+stgNpesK18
fccMqiRV3LUYCRPYoAprNe1PtTXsRMm2r+j6x+zTXsf6DhhZnI/jC+kNVpOzlfEzF6+fEcd0HAEP
dUQ3L2YILDztcinFLdAEBPLVa5LPiEmd2muG/YpgeQq89/aztVvRY4nT9zzZ1lSI3dGv0BOzldFe
URJAw7JmOMfIs9vicoCWBrjL5tMDVoaAzk2J6OwpLM+b10HBE6SMcQjGOybijSpyBKOjLNXo2s99
qGnmGYRZBf6zz7TSJGrP7LSuZ26Gr4ZiN2X791Wu0OKTRbruQtIFebs1CWCfVkGgvVSTyO3RYXu5
yFXFH8T2Y3VB0MIqX2VChlhSPkEHZmx26fOpNvdtlGFUNK6XQUFvw1YnNTJ2RbozYBf0dtQWkMna
e9a3s4wfv+kcn86a/SSahelkZGasd9C2KleY2+Q3m2eQTMgABlIGZaaEZ/GXtPc0s9GgWHk7jC1R
Im1hQfTzNQjSov7LnF6zNX5Y6yTGRQtsoW52wduj/fWHN2BoBBancMgPgUXCNeoun5kDlQZUuuL2
cDnnfMN5p5El6CQCZMroVmHAIS+s7InRLblnV5WjM8xot6+uiBc4LYVb5rFYJuf+T8Q01K0sK+1L
+fi5Bq2WDXlu8ohGTRqTjtnLaVTYB8k4uD2e9lqdLLsJYgWn7whU90T+RZJtVCIZOrFMi6l1saCA
e5t9w1p1ADRpK31xf9a7vbv/8+OI25JeMziHB3BScZ2udDwegzVSmqCJcL5qub6/0yHrOcH4GaFZ
+prpO2sawyDJu8zWm/ysbWUJgbz0492J92rcw0wP1FNis6Mh+EA6ssh9rUtzRVfigv7W/vd9aNtS
v9wgeMooREIKCNdjjUo5JBUBHGi9jXaHID3A2RlpNK51IB2KaIQzqR+f5h1QTqB9rNVHRf1eIUnx
11nmZlSfUh0xnKdoKY3f5mrIqCfocZ9qUmBXPz3C7N2MmauUrwXp/duNibKumHL/OApswANdL6lJ
7sHfvyIq/38wo1xBGsBaUQ3b1/zUSdxCsZxAtX6DbM4AebEvVXWLSJG5b9Cc4b4wZXE6vviRDP67
ai6bgIJOGc5tDuTYaiKcfg4chddcaqkYppQXnY4jMKf8eRxsfPDdPluVSXdzEIzhOxLkfSmMN635
AeSyeEdUJyFM88HkKlcP7qPtc97ZM2nK8FTlcDXe9JzIIZh3NpvE9UcB/uX4rBvIZzRXLqXgTuU1
kayqdgUpH3TJaYjbX2sKv6M2lIEtBUlb2MqSqIQJe2WY4XTjyU7pJNgpsToGaqS+tMs2If5Zj88g
XgkJD3n1BCc6s4tAFujdLd0gyxisDQHdt+R1Lz+fnjU9u9j2NQLrPx1VCrQaz+ZOltpb9IAqL/8+
VYRT6QRhiZGW719khiWgpqzxgT3odfdGGZskfDVXPpY5me40JmocmJTTP6oCKZ5w4NUnq9mKb3vg
TA7ZhXs5hPmxsaV3Q12IZdyXzkQDTCh33YQQzllK3FqL9F2OSfGgiQlK3IDBOYOIyX8v3zR8Lo0G
ZZP54HwSXKv5+4gKxUh7SbZGNucLhUog9W8PhFu4Mi7g7PXq/+7hUbSZAAjPsNta4FMjG33mNTEW
xQtgHZSUb+9V+ljm5o1VnqY2laZmI9/64CYFM8VdbH+dcbv/pc99axDiK6vjXfc/VS5Aqq0MP1e2
7uqgmvISKcDKFZ/jLr22WYzEtlcMygR9fhunPzx9QRSQKLW/X6XbWufi/oaCH1woJ58FSvSXWVZ1
ywQr9RwYJrnj9OBMfOCWdux2Bx/IB5TVTb/QgILD/cZEO2WHJjY75jkJIOgCYeGxqjY07MesaBau
v4g/HCzqhJLH4Ii1x4G+1BB1UlI4OBXddqGdtw5+s83OhERmZFXa545xuNYG95GIPr6Cqp3FCm7t
UvjvfrtQLrEIhPzwmouH8AribLG91w4UsDhvViTLwEv7PnAoV7FUKva6Ve2tVG66nCdXKoOcLhkR
x2jtsP8eZ+Vrrue2Z6gAfX4TuXP8BjeB8luCJqj7gN3r9p8/tBagAasD7ehVQC7SD2jfIid/3qB2
A46ao7prF+qpUa6TtNRP6ww8XI+/ytWc1rfmHQ1DWW6ugYmI5nqqzedokolKnxo1DL3qRD+UN1oo
PQXzHWZBGm93CvlibCA/lTOC8Piy8DPTsdq4lkdO/64GCVT0WLXRLPhqIaMFYUDqGZRrCfZ5t9Bk
DTThG7Hx7VPXkXFrKsVRcsLJeaa7HHaaxipz/EXjwIt5pXgRaeJAher6wKB+kNcfr+mU/O+NdS+l
xRJPpT2o0iwwg62+tk3W2nC0CLiPreAWHaXlGvQD7RyWmzj36PB3fq4mQSg09nklSzRAKEelWyDE
Hij6PjMFBl5auoTDCjdosbKywjO7A+DSrjW0at83sPsWYl2Do6l28Cf7nmcrk/u+te/EN/2nj50i
QXZGfJ8IQg6nxziP33+5yel41QEq2rJcWR47bzCLg9auGOPKCPB7UqevxIXh/Hv4rSMvBfBNp7sX
wYWWIEM8RXhhhk7QRXHWMDONAcMsDnqrvcG7PXPU0y1URfj0LddtaoPVDTMBP59PxeRsT3xnAdA8
a25Aw+xcFtzZbMX/Tgd3eBWPnu5JNv6+aG+qlhF9SlTm0iJB28wafIE/dpEQhpzTJj6bp6eGAxt3
eewNtNykP7dF7z4e4+3EFvbiPdT5oZ3glr3CBucC5RMUysEEZodlK3141W/vZJMeVY0Lxj8Tf8Sd
pJWfv3AjjGnayVkTuJdRROkNV0PmNS8UQfBFg4DFagj0z0rOG4wrIkIURwhPrSeqHN5uOttvSvQD
mhhCsZT8RBrzIDZufgoquNsCyd5eHa/548OGBlrC+nNrgVoojFeGqR9EDWk3mhCJ48TmW12XBSEg
3ExFqoPJ6t8kUQA0WcEHP/TB3BkUqZte9T2XbMPCEAMLmbANMQfNF8k+eQtSXpRNuGii9vJsGGTr
2iM2Dm2hLaiPgoAFoH4bafcI8fbw0f9wCgTBD5ZuKjdCFhvP6wGgfK3Zl3brANe529sf/Vbm2qtq
eIJNaI40WAmGybJRya/9TMG51BkiJOJxhCMS9M+/DNAM4w6gP8DrAoE/2+7Bp0PUiufqJRz+av0J
sqGjHfbwpeLRU1EKqrfR4C++JWCe7+UJWcGcrkb1KhXJ4Pwg1j+XSS6r6APC3kBXBHH2Zv2OmeUB
FxYX4deIaLQxwne32mcmoEWE4lc/Dz7vvNMC0CKmAiHQvDrh3cY18kSZ0FwTP8lMDjK+P11s1CKa
PfXmQGQ+YsRrUe6nx/DHyZWWHMTqoCjG/EpU2oZfZ886rgPjY2uhwjR0FCkhoLPNnmbubb4Qei/2
gDZvXa5KpTcYbfoyrtR5LrFJ3+RjXbtjl3D87Nkd/U/OvFtbAOm9MvVNHxYbqiNMXTljZqpEyToU
OFb52/SYM+b877XV63BbNjOdElIfvIxv5R5HQyLK66nNO2+kNQZoLrBiIQ3EwsA+FBTefD+T4sGn
MTqCbf0NJCTwf4gbL+Ui0lpk8a67fDQqsILu36XPdwgxUvaxP69T31DYeq9l1M3ZnqMrvpcfv4LM
G/cYtFS9UWnEor7CpLxdbLK+sfwBrm9B9b1fwFwFlBZCWOVbEpQTRa0fkn7GE+LxCDpEQEr9sT7v
txoOpOwujfEuoNwj0BQAFUdlSVcj6BcWeKNlH1kbxa97csklcrTA7bIQhMYs7clu2ovBtKkSRssn
rGNTdu8ea+JHfD4pjvcR6spkFwX/9wrJuz9dfu4UNF7cBXFtmScYJ471g6GgOuC2eSzkS2dZiXV+
Wz/cGqhxAduHMIiEmkwqvKquS8VWYOE47o7xanQHC7V+KyvwV/+JeAnpHUsG9rw0ioB0LUSE4ERb
i5l7glmbPxEoTW2HWZADgOcGVGHs+vhFuGb9N3GzKaxPj2LEGa0t11niOpsfcPe1ikDx7KPE54Ai
iPecca5bD9XNsnKbxLqq/1WgyVo82h0/plGpczmHOpDJadjpHjVxR97S7caa6UWb1LAfZmqyEGVb
Fl2ETcv4ZMz6XT29gv4Z+Qqk7EUldcFH0yyfdS/j1LmIwnDEnWdH1vUU40rPFW4B9mYcw7TihRV4
1MqJ3WHZoMM0PXq1yrhNhk4aPrzRZ3BI2vlxVcmpyZlIRjNqZyeAlHVQKlcXHVGsGExIx2e0qEiD
hdup7A6svk7QXronoK0oWD0mmSr0h6qcfxTFHgTJSE5sOjGZ/43uRRdKKpX+E8uF2f0IG35y2B8/
l5cAIYhAaro9g4agyP1DXD7kTKIMOSclD2LK4ET7Oos8yYzg6EcLEjS+kgP9cKnEPHEXaSjzH8fu
/9rUgxqnmtEop4EIXDWoIPCvXuNVkyIU6edndLV0iBHTXfbzuCAck3/LtcUBEJDOu37hWUdizh33
VOSANGK7ZVqAHDBLIe1kkFv4+YyLl3KPYeZUFbRnFnSFTSW+EIOTC3T6+VQjBs46ioPafVU0kkPK
gnSRbi3hR1b2+0b8FyvqL4mtOtrB+yRHqnuA1yLtMx9sy2jXM/iJykysZPO4ie0ufuKDrbMTWnj8
M+38bmplcoJs0/UTzzfIxo0pv+owKXWzLZRRRIKql/j3MOoVbgqVTcalsmXjoo1uoLjKbwUml9mo
u45BPHh1y9ZqZUCz1TIlK/82rLfSq2UXFyxWy2/J7ujQ4o8693IbOtlrVXhUgRtDccqGFgK6H9mS
XkQCOnCwcQrLC3CQRfYI/p4KatJS+8CmZwx5AkhOOQavZtXj+tms28YMFbcEqRkwPhhQ3mOoUJMp
sED54YQk57d9ejMCPrZpxohvYQXuIrZfGXKR89chEF4XIe6cXyvz9WDxhC9YU5UBC+VN3NbrgoT3
XAzCLiqDRrduh24AGuS57QoulgVjfXKVQFTlzMLIEew5nE3abUfT81cS7jbFhaKJfKCtO4UjAInf
TVHqB58sYQBR0LXEl1ngSqPKlGb1pPos7z5GVT2yYf6ShYrSpwyLBnNmKxu87i1SDkXc/dItn6OU
MciXw+8OJEKZOkgGLUqiU/PRaA48E71WLJFDKqDzRWtArjv5+Q2Sf8RIt3EukttUgYTyl4Y8aabW
CoFOv77vO/ZlN5PZPfJKcIFU+5mn9TfE/TehDEk6SbrV0Nglc5zhOYjyQbDRN6S2kwxx/YK18Wza
oCemPi8Ir4WpQkleQPjs7YFQunFnHOVqDzxsOS0sNq6wbmfk61EM9orPPyqzmRpTakRvE8JWwUW4
GSlxEFNHr+z48E5Dwbjk7ZWHrCWsr9A0WNkOsYXTQnD8UrLGacgQxEd5OP3NQoUYE1CAvssKste9
EkbUCkNyfSbRzX80dMHEMlaI/2LHh0U4lv3JvrlhDlv+ZrP3YtjnOVQ5vBIqqhiWXQ+rKW3+7Jkg
QZrKRNJfZNgdoXTqOwdxJ/RZvlbZol56GQjXkFRe4NfcDfxWVqMvqxTNC1TS0OW+HDfElFm0AmIr
84dV/4/5ar7IS59d6K8w+6ek2+8WUqaKOXhXBCu4gD/LzzhjDSX/IJh2Ds7aqrfp510rsGw9qKGQ
ME5zNiQ4DnUVp8fUazkp8XZgvR9hW+MqFvcwBj2wV9obSYIkXrXKGy6uapvbecHwtbGcOJS/oDuF
tJG69UrmraLSxJzX7YbklySeZtOxeRpftUvZ18hReVXDbbJGAgb07JqCb7j800zdzpSFbOIPiWVg
spAvaipzZq9Qi0jiRQ3/odYDMUafDta7TV5s9riDps0/Btcw0Nur57TZ/K00HAklodohNyJvIw9X
Pv6HRP4h6IWpR9Uvwmo97Tuse57t6uzW+4NbzyIUNJcyQHbClerPD8FuwFrhD+EGLTPoi2UX6CFJ
2vusbDP7rbt/LZAB/G2okQWXpAkl93wUzsZqtgT9O1qJIX/vXBjjLE/UNK74eGydxUYmZw4T1Dp0
4/O6GR91sqppVW2oWz8wsgsu5WRyVFGL9M0meJcHOrhgcGFBVDhbzEhwyH2lz2TUuyMJzcQuO3vn
iQjfcu3prPP1KZ6ijVbd8xOUosO2RXCHgE11axkw6+1Uv0iGj05dkuw//vHIjQ5IwcIpLansZQnW
CFJJ0FRonJDeFJerK1UnujkOsce3EyMB8t74KaW9CtxHgUsfwH/JoRNFzze9TavXMEJoFaadDHxB
vaP7weOy5aQ0E+Xbl+i9ozP8pzYqDUfFcKWqCxIu7cRRbLX9yKSnLL/tAAkufzYYa5LsxyD0MJQl
eHlTplPEiY3kPb1XfyWL48cUUW3rcv3vxxRv1Se1dQjbT5oC5Mt4KS+ECYTAQCW7dlF8UGwL0Mwc
ZiR/qpN9IU53lXS6Gq1py+V5DwutSefmf4zVXTtGyiY89uiqhwIiDRGvAfy+DP1fwiPt+Zm9fSqJ
LnNXsFrVEvEmzEkMDmwrdKHFp2ozviecaiI/AVWfZ53Q5AQP6ek71GT2t+Sb/fdK1895xKiwmZ2s
NLsF+RNvQjsuEqErbgbuYnGSVUhthL+cMOm9g0Z00R7QHK/t5Z3SABSm6P0RHzf383Zk6h11+yvx
Osy/oIQWke9HEQPdP4zAw67agEMcdNg/RvyFKnIurjteziIhsnf2v0vxaKVatkoj3lrj+6Hy9ORh
6a9Eru6keT66E1aYxUxkF5fqf3P0XePSQlX+TSqopq5voQqLu8Hnfphzc1lucIWIG17URTgthrhc
h9Cq5e6kVbzBSHTn0j3phkIxZc6tqcvco9LnGbigR+Y6+FFr2B4ghK8PfuOpHJGoRlf2obL/kOsH
LSCjmqCChX0RcOazx87ua/hnI1A570aC2nF3w4fR+p4Gl1sNpg1F+1QsVHmkghTgje284j2LiHbQ
PRO/m1GR/o0WhvBhE1pkL7siqxZMUj73qJRl7HLfX5F8jCeRF3ul4Ouei9PBP7NvWISyOpmHhQoX
VkRgLFXWdQXogmtZcyH0CIK0NOhGIMEBZ3Ta2o6KHiVhMGAxTOLzTx9qcDDb3JdRSVCW9uYeZ3pG
B6pJ3qRT8VKVkwRlsP9vjBoG/mvJ0knYGh9L5nIt0b8Wu0CN+Ngv2KSgjN6Wq8zOgLpSCITw1B8V
ShQR5idXp+1uAL6tIL/C6BP/E40v7Bxk+3XyXdmecM3Jl0Su7HDaOPl94DPRQNr2QS4R+oL29ULZ
4MXnzMXqfolKR9VoUPzMxA3HyY7ScoE/ifNQs3sezJ3JXWOdafSMr0vPU4M1GtiXhns9bxB6FxCG
YnT30Reso0iDcnwBNJEl9PqLvCs9YhRc/yGSpzY5Np/auvh/h3IxkmGjD6b7SGLTMxXkGhBd/ZYY
D/OsiraHzjXAgGsddMFPi7X9ix6AVSerHTbmgshSJCNm5wfjTH/3VfjeaeNkA2vbIj94zLExaFTI
3IkwpjDgXaQELqy4eq6Dk8FgNlJVUXQjhQl4rE8ErJJIhVk5WhH1zMiGeYyO9Tx0WrRVHrGyVUjf
QA+4OS8wWCrM9XhEestVO7/F/KaeFJwkSh4FfRruxvoluertbjVmPE3eLtVAd8WRqA6hnImlLl2r
1JhNu8OETmOq0/Ir9RbJqVhPNtJX4BbeiL4XAp1Ilr3YwofTVc1ULyB/CuZC+E2UkAyzakREgtMA
qXlTR9bCcrd4fbDJkYCPJftVe0rGJVKZp5Irn7wcWBNKCygn1Ig4qyiQYE87YZZMgrjbAsyLoQBn
r8zIv0mB9CdZ7LvtxEglaOiBmALBQruraVezr/LNgRUBwoVx0d8cU3c6Lhjj7lM0+oiRZHyUDTjC
ubmjKX/FGvtmo4s7dHibjsLjU+EjjqXH1FaNW0KBNGFlUwCyT3+e5aAeUHezvo2Vs3oWN4aHvzu8
YgiD/3OUmV+M8poSpeGeNjQRFfqPyHBPvYck774XrJd14g30jwlkfcsCpD2ggZmsqa3qpZQ33deB
+v2x8J2Be8hiF90vgLEcmzKRWP+1Xi8mUvELInCjWx7zQX1eIB41EFxhuXXP/ibwTXWjk063tyaY
Y0245Ow2lpuyhDbDNqulC5//vteOv0v6A4Amstvx4HYJD4ZYEmLKxyfhSZ7CIaTT26BcluIfBYi2
JumCRXGWZ9yjaxdyAT1MD/zT0pntTvRvYRwYcisTX7SKtF1DJwt8TLuNe1nq85yoabz0xoWOWLUN
lSYVQHIUFrw+JKDlkElCKe7yCOlF+6r1JCXoYyoqie4YKAf1KIb5JDdkhYZ2Uu7Drw2LTH7pjTr/
fowxEv+lByJhz5SXwEir3wjA/jD9Rp9euEc7YJEfajYAJrCttXrfwT9wk9WMBToGTWL5HOxO24xf
TuiZIaS1LLd53GpIoFuX1nQOzRD+BQTUH0dwLxRrx71UeTL1ep7qHVKcmI/ekjDFZ154hqsZRGBE
Vfa3I/t+6W5HFN2xV369MVbINShaimkvSuvfxmzSjE9EelJHxLvGpzPbLuaZ3v3Wz1b99LUOgooF
Tcjt4mytS2SSH/tlMX5BrSgHFE5cI3GSY0ZHLW9m9tCENigRsjPqHj+prJ456rwkDhOXErQQ+aN1
hHtwbPJhJ9Ytw3dhMFmWRDpIoOlZT8Xf845SAI6Ag1grtwgTiivEqKJ++IOGdfNlBMcvtODBTIiW
qT/TaYq3Ru00ZFvO9z310Qy/X9+deha8kzvwig6MDi4kF6F1QhlW8234hRjW+wc/XKCrFqZ2k5Fi
YopjZlmoH4nGNeFrhRBZrnHfBVbqvTAuPDSTN0GC5ajBwuD/O6JVp1QK3VL5w8GE3JAAl75El0E/
w2w+NX1HuXhEyZFkmnNRvcXznwX48N+2lPM0U0awkrDO2nGRMYfbnKqrZnslhqKGZ5nmJkOEs2b8
4kcAmOKkk9xAlzRovaiJyuxs+t4vcDy25bo6ulL/PN0kP/AmdRAt5dz5gH2wPXTLdkfkX6sP0AVS
7P1qtmRckPC9gy3cvHxqeHVbgvyTvaXE9g0VMTN5XBhtTJbPeYle6gIplRVzhkeVCFpaCyZkzHcd
5c+1m0qjfflCjaHYp1gtVB7b+ThGqYO3i9osSL9s0KGB8MwX79DyoG2+vwAfxg6Ats97b5WgeEv2
uPjQizs/fGNHVn7KtSGyikTsfpoJuzxB+zjLBvBDowSoeQkkkz+4VU++RSE4O3dSEVoB9phNYJX1
EtEt8RxRV44mYFih9biNC7YbUvRxNKwp+iQSeIxFI1yest2wu50ESVYyUOq5wV7NJ85CxFBQVnnJ
j5HJGgY3GCVSjtG1q7cWorLkPRSaTVt2C7UOMYdfwRrfPcpkcC7iIH/tkvk/DBnbjY2hNCGYtVFs
K2kGmXpCNBtJpNHz6q3EdN4XFFJ9FMtlvxHOX78RkVJ5mz5tHwJk1TyEnbOml4U3fjIrivPziZhm
LvXmQnVa04078pt1+/YaWvg3FHl1uUtXmxEFZgMUMPw/lWlRQigDVMOGbhkYomKVIBpQTtDCyDnB
frmBA4Q6c4ZmXeTFy94LucEG5uAAfoyc+bha+6uR9w1mmu7zUnAITumrusbKE1MAhOhP3Ts7dPvQ
xPzHy7rO23c3kl2i95IhFnM5JLm/ksddLTMA3oHulnfv67s+MzkkOGKHWFaDZ3VY/uqkRRcgVKwz
3AgweQaAK24OoHCiBYifwwlcQEywHBweg2u3+CkU0dbv8GMaolz9SByUdSrA1XgMnGiuZL8Ty70c
sRShQaBBsdJuritcM/WMSDrPaNIg1eFathTpNDGGVt0h5WtmbQzfrGyK436yPmwccEnIcXThawXB
4ZiZNKoOiqoIEUag2mUbTcW7bWDr4Q134iynoaDelzh2HQ4i4dNGjd6NNuc/qHJor3fXpiOrA83s
i2b2HM/71nJ2F1eOAvMVzJbaXJfGFady00zUbSTU6ahsfHbAz8kiZjXAf5zUV9wI7IDUR/2JIbBD
Uo7Ixj1ECMZJEsgjjolpnRhBzWO8pElEGsH860jSz1GqOmraRNINECxQZVqRKCa68tJhA+RlDdIn
D4HVvG7t8ckuL6SfaFZMhdhaMAPX43FwgHCsACnWdRgyt/2wZcQesPFHpPgg4NRt0zO9hWz40fQu
LZm2l7H7NW7RjFUkyy5gm8Oxao2tTsS3/xGLaGAh4Et1K9fySyo4ZeqoL1EBgL7xtgAwzp310nsf
WpfARwXqwrHcvfVH997bPqo3WXRqZ42anMGQKeEOPFPcclNvxcvwS1fSLMQjhbumCzz1Kk7HqwuZ
fZdqwB9PwgdWD7PLn4mOhwb82uVpPPOAw7fb5fxlnlOv+uypZwn+IS0xFdauXt+AvN1WCPEvHYPT
b5rvRagDB6Zf9yRJ7+KCwXlR8Y984j0yPL0mPz6rlcULqas3G+wz1Gf3T5fTXmHqlFllxCHFljAS
rkir0Fa8lg/saWO0zQdp/by0E5YTUkpLNCnBJxMMWDTn84hf5qRKt+8Py7pWqxQF+fU4HdtcnI3c
oY2a4pnLd5m/vmR0nHxLcXmfzsioFULEUFROL+pgd+a0TLy+H5r6t5uI0XHyxVEn8+hKgA7PpuAx
XB2LFNhAqH39eNX6NqKqWrruRrGTc3BoqGVxbgKYzkq96bBqG3i1hwj8lQQwKxuGHPnQtlp+R4fP
fWh6Gf4TDIPKcPXiyHLNg2lgOSiYW8F74jt0lhQg8Y67KPl20gU4uZdgAnMXlMhDk+nfwZROJE07
lL9g6DzmY/zTVgCRmRn2ZDBgH09/q6Qz6Egvx4Z34zEq9v+jV8e3ZgcgR96Npv4NcQSddNFxXnW8
HPwp+acvRguk/RM1ET1Q6UuXDAKuf2A79y8vNSmMYsZWkKcM0uc696CRM0FsUa4nhM34V2RBMa/0
Ep3ntm4LM/+IS/4xN3XcA+MwNbsHP1T6MGJJ3xElQ5P7pTSoV1WlHNosgamLhxU1SNl4rEaOiqbB
dhnsAFKWwbWKz6Qxbm5pNOn5G0XTOSN6ecRmE6/drF/io9zwrtIm35OJpVLaDK3d5N5rs8AhMhDF
xkUrdFdrbVLvpY7vxOKzRMYwwhD3qJb8J3RmSghvg7oKg9dGYo1u87oYsJK+yPS0Utc/w+qrls+5
pHoOVU1bBZmuhC1IegsS+avrgMW+BIoVpnkTiB9YZVrQqDZKI6jiuP5iA2m2vwIl22TFdpXvS46Y
1OeXwtSwq86I/rxfAlhHsw8ekfeK1r+3JbuvyytYEuCa0sej5bg/fUWEO55N7XDqL2BF7fgm8ygK
1entOv0Vu5PaJtgJSCzE2PMqHCKKF+bg6XnHOvhqY4pcvuE5RqVWgy3zx5KqDAoW4dfFo4S3AzOU
nF7ljrSMzu/DQsdSb9Wb89hKnrIpVk8hCOKEEr6iyOm8taLzGRY1G6Ui8FCaP3iUTaIrjVrbmtdf
qJjgr1ANX25RlAbuiL0dq8p2dvaThhKifmjIZW+L39u97knbC3MEdXA4UX3kBGNC7rhSIljJJKCC
o4vZRnbtgismNUNL3deaBdf3q/RWlh+ivDwRQ+h59ZnRNor91ZjmFhyW2X7C2f3AuwUk6VOF1ER+
aA+o4OjCGS6chljQZj46IL/972yAVfz3QMsmqcB7orWq5jQldXcaNdRIF6pTiocH/rh6gNuluZT+
e+XA4/hbR+ePc2/HYDiscxizr49rSDtuB4km1rvqB7HX4ppsPClSDMtC5eLWb+AwT/oeKfLKEkjs
2rzW3Z2sW5+8hRTdhbf7aJlXl/gXps8UOZTfw0sRiqPSc3iLU2GAjddGdYWCSxctqDg1ii024FhW
NfrHqsFV7uQvD0gOAnr0bpJy4+OGEQJk0S2gGRlOLmwTXF8IuIcL5qD6oxt9C9hhnhc19wJN83oN
RZR98bavf0nvuoroL6IU/kCP29BE9fes5H286fZr9Nn2L6cJvkiu+7ZQCMBxX2Zbyu57X6J5k6K/
Yob4ueeoKpSiw430o8rKyqzIHRQqqDUpAjSRtEnlH0lMI4JkQPdzFVeARzSfyj9OE4mXKzq2zLce
3OGY9okEH9Qy6vZvDAoLgx2zu8XEYg1V5Qwnf5B6csQnXjMazH+oUifgJrgozGgDBg3XZcwZ5wi+
/17X4+ZLeHtfQYVDLMrDuS/in32jeAVyDllP45CA3lIhVyw3qmuDE1dgVxDg3jDFSjQ0FnWnbnOS
5S/1CtXtg096AWtsUPA+zcQEt5ggntq94JadGZxyRXMFCnPvFsal8MbjflnsDZOG46a/awPoRdjF
DwxWF0Ol9Wk3fO3rooPLSpOlyhQtZm5f4sdYSVqZtOMWcsp4U+RCiIQ05Tig0/BtVAbj4WvUTTyl
ddYdQa8l81I2yQ89CKnBn/nDffWdWq377pk4WPDbFdzmGkgQw3Rd6OtVCJuYniqZhH2m2gLMyhmN
aEBq4YF3YF2S+ui2Dd++wA0HKjn6LhWI8nR3bCHgY2QDpcrVjXUbfKeOsmBunUaFUHWBUuZGupOD
EtJsgVRPl4LG3Y4vMbrf6+r9DzOhv3+Ede0IQijsZGgDqrzqLC/T7YXy5dzFNmWcXrsvD5FwwmI+
3gon3liALGJBcAxFBM6EhVbpGRd5ftGUN5DfauJ5ccz8/oMQzEDuc1OaGBJ5XrGgIuyCyo5/2Eww
yMVmnf6L95POYBQILA1LeQQQeRToXIwQG8IM9GySp/u9bLWbQrfrKHCWC1dgW449VT1NTBmlwtKs
UX1lUVvwziARgUsuixjlzkUbDzrOznGFMFMZ9s4YdEZrjLyNOXanOEG6PwlG7VV/23MxnVS/PY6A
X6evabKqexeBEntJhudGqig3o10uOwRMum2DweUQPptPSecFALXlpn1QEXFd+N+OxQC1QzOjA0N+
HKpDQPjD8r1K820OM59LacFkDIApuahhAxZqsxvCEP/Gl8Z6eca5R43Sk/vAE+KMZ2O8DgYTpnE3
gDofJtXh3r5beMF1p/C1Vm/aF/9ofsBtgtsIlXgmS9YzZ4VTnj3rqk9DSkhOEYMBHw2DPWfKCL5F
vxqLy2QkKFcuarvaiEtbV1RcJzP1lHsaiJ3jDUXvPjkDAHQT4Gj9n8wtZQktXMbKn263f2xrmvmr
TtGsZSlN965s8jH/nuP1r95ibt70TKHhJLIzihHXF6FiQYlR2JKBFmanGrKU2tufB/QNdHB2pXp2
f/MebXmrVzyFfnxrvrqe97OVENfHSG8yFU+N7663VApll3z69n6IiGfdSiGMCvuqxNH1YvRkP4aM
GVdPGusF8FpVLoH/qV/JeGK/iVtuiA8ePzF3jWt5IXsesuNU9jA9MOzRvmC3CCoijnjBVp02Jcc4
3+Yp7Oo9SKXAexEaQY9GhONHk9tZyo/s94DvQ+wvHLtbCrmvBpn23H4Qg1c/0ImOhuTxQ6x3455c
okmnDKnvVbNfy9qF7zGFBmdTQXJ6NuwC97Lj6YvooJZqYu1cGY0F7eFfs75WXn48uh7S/82Gxq6J
odCZjoPt+TK2Z3usn4JP876Xmp+F7kmAHKujFwSLh0KH2xmawZcnrysoh8rMJoKp9LeCEU+2pr0r
hw0NnUMjfXPFhmXv6yDJm3PmJz7AOcDWHqoBi4gz3zWImo0sMJsr5qlY0t6qJNQbZS9LD75Okgyj
++VX3FkkTa6yI4lIEHBoetE6pf3A5H0dZhBfVnjW5y+nEbCkGBzMQ2guMXd6hqCqWIF8igXm1lHc
FiyIUY0BVNiq6VeNw/FrADAz2QzZ3UwVb4dZFHqaq/yxBm3/9oHa/Z9b9Ox9XglQky/L+WiQNwnk
bAWo0w1Xi3TqUx+qTEaNFj9RKRHM2HVcKyYcoLoD5eTDD/GboP4lOz+NEg7JVXC5fak8kaZdXXjz
EL5SsWVLVf3LXMPzcuV9yZHq0m51lLQbI3ZNyeK18D5HZVwUBWPJpwpdCNBPxkCTNFED9KNTfe0H
rumK+ZuzHnzlc4SZZEvZ2Vy5P7OeE+LkCfHeD3tth/sTDj6ya7LI5P8Io0KlqIY8J8M0LTfg32x3
hJ41M49oNZP+XjLESFv3KVgWoDk39GxogfTdFZyTBDDy1qDcHxlzVCX50J+nF73kEzHvODvlNtNV
IOwchVz5OAAN8ui8paJYu/9bdJiD3GDiLe1aMiVcYrqTF9WcjvNSZvsQrFKawjBov9LvXALPx38I
RZiFOZg9TY6KDdewuut8SrSRWIk2DBCscGJzebK8p+BKcilOzbsVh+kbToHpP55oBdzEiNdLvs5K
uj7I9Uf835oa+llv5cdQ1eQe6gLe3/gbqjVEAgU+7IeGDWAFklqwNQnrAt0hyIqorKD974ihw5sB
ER7pe/IxMZnArHpQjlSbBRymCzoCfihdiT5EcXP8Ztf9KuOejDEfgw10+aUnGwKnQ4ZEJH35nyQW
RoDO1YY61GtJOMIgIp8l/raKsjh3YT4kKNpLOjW28mKq555io49Rk+xMNEOPrFQPhwRdwtCTsPwK
LayE+H26vClUc7TK9OHcTU/8FtTebUslidbHeSyLxylIy6DmIZ+OV8g31kw4NnKQyDTxh9hVy/uT
q8yc/pLqBqOUYgSrop9Oa6E2viCCHkG3lpzD0A75HJ4oyURS6ywIxduVxYKmQsqCnch9haLZtQlJ
6y/LPDWqYGprU7RIfPGz8MnJRqTvWsoetZ1L+hR3XSNr0QrRJgWY2gEvPv8hCNl7tBM//tvCNez4
vTMnlWliINRXCdORXjyXke7enjRpnOgDJiCdKPS0PVj9NoAuCTfc1XGqrboxA6anBuI6ROFd4poh
MVCqBD3N2vN43Eg2a80L//bjuMH/loCbABks5ENfJzaL2WAfcWYbbJ8ftHu1YvY0TPYNGLuTijZi
1ZzMw8YK4IgV1BOPPItFN+IhSt7+UYV+bL7gtRpbTPunorYwr5Iu1DHzP7n9H/rVq+Us96UcstnL
QvLi8e/8RFrvAeqJMmshfNA+kDoUvwQoXL9SFoFS2Cl49X3MA5fJ2EAZlu+y42tctspjWH4fVr3p
ae1Jyz46u127fJOKGt7JTUQlwKKuVE13SF2PBkcJP65N58AswKs50bKS8R+0ocQV8CnJP48Ilwla
nTe4lRXBIV5sCKBCP2FAnnzjj6u10arbEpYW/Op9W4lIoxxPQucL8z7lxuvA4Ggx9k78tbvE6DWo
7iFH+0evEwjDNF9eTXkMNRNSi6hN6tmr29ClPv8unvG8qPWYANorgGKiw9aA7GnrCDG03G8xZn2h
xZ3jVVOFAJEKkVMZ4gZuiXUPbE0dqpQgo1gVR+iQdhYrIuhkslQxJESNcVLKSZVnoRcF/1u7tI4B
EG5DpBRLpndEvIxjQCyHt4hZ9IQL2bd3nosPPOYJHsA7uSub+PMJIb+s5+Ldw3/2+wsj2iOq0cN4
ys9SzN27ZtAH+1zFEH9CXLyiUAa5bx77hZwbV/+wy8G8bn0RQ/u3CniJkOMxwKna/fZz9saywdZE
ZzFRcdeqmAOXZFIwijSlDGnA42uJXweyjnkzerP977NUZeQk0TjKKjFDXV9XGowrVyaHXHJZf+KD
LcmTk9K6fyigOQbKI1on56Mo7e7adVywcMnWwXKFCUTq5CJdYb70loXIO5g4wyWuwtqAbowGMu+W
aGnNxRQAaezIFxkrxopFNa8a3hGM20m+0JsD/lUHGXlHigJvV9MCSBps9teOjTCbX5LLz34Dc741
A2uaOFDT76hWTO7w5OEbGlpLMH5ZavTbCLt6NOGsz2eIQZPz6nPjbIXN4MseQwZsEQrQ0bqKaUW9
yoP9Wkd1JOKHH8X75k64vS2+nBXv9Mj4DebycAXF4/u6WWa6bHjxKDI9F1EOb4vNmocABHqMXjSm
MztpjFXcPrnk8BQs+uzqJ33zSYSwKiRFQ3H+BYKoici8gjdW7t/bifFbk4nofbH1VqTTOX6BgcL0
QOyJuM6/m30G4uljut7gCTUZJIvArbJla5TgDeXKhcgfwytWLUBS4CLUlAkMb0hpOtsA4ByK2xt2
nfpPXXeKri4HG6yPYlCmSxHjUDL6Mrr7XHUv1bPSl9Hbzlis0P1hYzNo+bk0GFrfB5UKFvI2NqVh
99Q0jdhSXV4RdUWcIIVxDT42c9+edsVZJTMyfrnCclfnAsMKyWFwFmt7klLpT3tbXIgJvyDPSKOO
ZPdCC/QkhxsSDGR5yQypMoS+awoawS36MQwhjsXICtJ7rwUTfhm7cTnnS1SiBYQbSc1Qt8mMkXPE
HX21Ljf7vm7hoaG9yyv+1GTrQWYYxG24XV1EPOr6yac05JihqqOK7/HemgDbMasYDKe7B+Tg5QxD
jzVOABqHXKApr5LSi3e2GwLkVBDztZWx7l+Du8GAOm7nf6d0rtvy+3FsmJ1UAkNMxMPsOYAQf1g7
Mv6M3tSDqXmPZb/ih4xUqLFcEYs6cDqkw5N17xVZVootBfjzaBJeMAzlhMFeNc+FvEYe1x8Rr3i3
WhbzOTF0R3OPfbIAf04A3ZF1dzKYkFlFevIUiHm3MVKaIYG+BcqTGeCankgic8rYoRdJDBWxMWVj
OPaeakD+VPk82ZgFuao+ecgEmDW2Wpx/HSCi76Lyl7HKd24KuXvPLYgYl9MXQ81JVt/mtKJx/oqP
3HS85uVJ5wOw8pmd08bEZ7PTk1uu2UbwGp78MHAygpNAI4yWLKQEAVaRd9KALLSePGUM9/gj1Ogd
r8PSfiYil9IGnJkWKrY5gtCuS43y1mB3Vy32Ri/qXKpoAH4IaTdqaL90s2SKaSbirjbDnjNf9LFr
UU2lIiXFtL+x2ReUtjjV5hiGrcKb812ynlGol/DA/is2TigVpPfmA/cs3+QGI5wizhwNS81nb4QS
ws8EJkmzoZ78sLeM8yfo6aVbn+2zDDuteiEnXYspK89fQ3b7NbgE29qEy0crs/oB/10o62WvjkXz
mocjeS0+BzTZDHcdFh4ZfWdCzEgOE5ImtK9NmpmFPSj1s6hBB4qgBYaFFTZ6ogPO7d2djxWlBCQC
Nzqvn0RYMDjPCH8yjnoMOGYGBZdFpVLi+/jmxQlcnIybikN2NlpYiPOCjLzT01IY9HvQAXu0m3jU
kHI5SH+g8XWpVa/v6NUW4OsfML4SbsFUQK1qDjxMOp/6ZliAx5t1T7CJdhKlaZykXYh+YAelLt5j
/U5+qpaywn3j9GovA/oD33nyL8FXimBeq2DHuK5E3PnuTVTh86/uLa3aVmUmlHzI3LX+SVNw690U
vTJXIVJME52+82GqizGr9eNtEKIK+gSbIV3M5MmT4xlATJfu0EiHsM7JojEs9ckdmLRM5P2cmB2U
eiTsH99A1H7o6HGoXQPaEI5y3Og9x0/vmCeOqFEYxbTrx0aObLHZWx76yIGem3UJbBIbjRKLc/fP
b+bDYiAKgDSro2HdpW3wBXf4bfDQm9XJjoWtpza1ojvbFIZbdmK5SO4bEb5aw7NcSFLICzkh+V9D
tksjoU3jetW9mmgkS7sJXqHEm4ktkdnDbuGatThRapZ+lculiEf7hCH6o1YvMhgJyKf/p3SJPlaC
SS+g9GLJJkrueOm06v79vmECCbeXk+46ICPcWuY16R1F9mXIZYY7l8l8BcDOz6KGy5TmlxvoCH43
RKjnSEAgvZJn8Jk1kuOidxUk6rpU0Bb9NsEghK4NBA7RUYQh6NHLr0JIifRh2VWA4Z/sAudl7ljf
c6WS4nZiI7VBmKCzEyauCpW3IL+m8IagtnLWLJgEwru8KO2WnuK+mDsv2wI/PMOmEoZDgz3QubNH
WLu8jKY9Xs+B58bBay3o2EnLkeRknu+T/evhLCoL3EwOXD0LYffuDYJKibCue9R2F9RX0e2yJpg0
HHawWT0h2BVs/PSzc9cE2jZHdikL4ferwdnw67tjKc6iEno62tGi7N2N+1c7V3yobIsnSl+EnPoU
4D9N8OCja7lIKxGxvhW0+RvseNEQBum3oS6z6oI3ZLiWZ66r+TSUiG76A/u1YBto0gIvt5/LvPLF
LQRt2ARDy6LEfOi6g52VA8fBX09QZULMZs2Dduv5ru9VAUdej2x457yJ2zBWLcJaRQ8ovUFiFbEW
YWGcUyvzGpkEXaFnhL5VNdZ2mO+ZRetreTJiVwxyFmbKBxdPtvG1TERAizx7op1jgB50lo1to1g6
EKclERHhnyvx5/vYGZb3qsgLsyo5yZJFS6vOgGJ8IsJY5VrY9mujcGOgnotjN26u6gupodwpycPX
zH6vGw+0BahZCmO++OaITqccOZvD6S9iz8MyymFKpxa745AOb2oAwdSXEh54n8LGZi/CUZO7sIRQ
n5lOI4yMGZH1KWAirK0dl4A+58IFFs7+t71tm0XqgDLT2t/go/NC1UxVrl6fOzElq8SDw/x/M2GK
Q1H8AjDn+qVWfJek88UqRuWSZSV797Y/1e3lvj3PAhpRNh79Rd843xMoAQDZqTlW+wrmnLOH5Aai
nrs2GGZnApSfXqgZPWtl9kEsoUiy41Pvm0twXij78pUpxrNNFQgxRqK8r9g54fiTrtbIbnDI/3am
MMBqt5XdfhGiAFGamWxj8EXU4WcATwXrWkpePIR6u2Cc0wr816FW8xEm8AdixHtjPipRHUY12Tif
iiZWRPOuCEG91+lc3+YDO/QlOg7NzHurR93x1YEChO80fMYTu370oQIpYP9Rp9H6JDWZ3UMCQF7t
Jododv6r8eJwXu4qhswBPfJ/bID54LC9uTpwZq+eIeXfVolYwtW/0WIwZMtXqeSgMhQiaaLQRKDZ
JyyvfFnttLAhtYZlKwTQI+uwKKbmxIgmg2PNm0TSlR8jp5ZNAkAlmvcJ2EHKm7XG2PehPyMdJkYr
t3homo/BUIoWEwAk8qVLfNbOV8jJjffauzab9sPplM+1zfEMbEBb3e03eF7Mjfq37SJ8Gex2m7mZ
WcRL9zMDrOP1s79F0erORdpu5aMNYR8jR0HwJKiRH+O3mqAm5vtW5uldBpE8pzbT6QvBHXXh8EYz
Bo86k/8lbO0cSUrD0mpT7Qk7HIxV1V+dZ8o531AoOOfkRaBGeB78935qjMjSw413eY9olNUNtDEA
sHWKOvTzib6DKObyNlwkEFsuhCzgybawiNLSOZvishoUPV2Akc5EZ0O8XbixglcLkU04SCLlTzED
pDpDLPP6pZ2ybbjAj/VdJj3OZzFc4oJHvDWOb/I/MED2zD/Sh5mLXUoxn+JMROce8ukOHiFbMptj
rooPl7/ImLzvTc9OuGnrDBjrK8V5xaWq4CUjlzwIUjxm+leCu+DKXP9wg4r4CRBhEd4JeevuKosl
o0M/v2QwquG0EFcfKjX0T7ZxNIovJVYKZiE7jI/7e9h/ZWpNzNi9WSVuHPXtNUYE2dGGf538FgYF
vL9ZFqNnwEMenxdmErLuUYcBGLuYvnJBwM83utRIxkX5XraVnPTHGpPiuQqtXUEft6/3m9Y+9mx8
fR6qb2DuukrDlOIVJmhE57TbN199gGnrAJ/yLorPkzpfNZ1nAVJRGgUeBnsC68Ti3nmduf9SiIRs
3OtxN8Ee5WEoTWbVLRJ2ahR7jTfpoWktxQ7cSv7gvnjb98G1v67fBRBjh9k+rjUxJAk2kWkYjzcP
u2/bULdU7J2UtMM8yaysUvdNd291i3MQgcbvzc0KA/Eh2TPvbywLvtVNXqlDPTAEyx6cjPQIG+3n
VIdqFbQYY1+itZo/ubIZSiJazweLX4xu89aRYG+vMgAXuk4S6Ufvxb1hoWywKEnd+CWd98nGvdSh
wbgm4MHQd1Tjjgzq3MANIh19jejbF82WWuIBcZuzhasmH9UjG+sg7h+KjFIcp9RuCVHHI2wVqRcR
FIQa56DubV5RNxdUon7GzKLDiIFzmbBiA+bs5jAFFPdaRPq+sGjjSws/M34o7/Va60Z9ToXrtIAm
bi0C9R4oUXtw06PseKcsd2BB+tqW2eafy++YOXsjKmz8DHnCRyzoV5BYaIeiYuu6eYg+pL8xEAbp
lC7BKbiya6dO1J1eHbViwZrQks4WMGcUz09I8aD7aXXVmd+5laWOH6htyoi5R5uSNz6o5h+CUmQA
oiKyNvFqvAWvHeGQt2ATT2rZqkFWA3xiCXIFRPLuZVHfEl+gKzxM4fS0upzwBRfx/kah2NrBnKMh
WK0iE/Orqv1iZZQkmhT13lNILc3acTfojgX0gFngpfjVWoXP5jKTTci5c9IpLj3Lkwmv6GtCJJE2
bXu6/POCA/paL++O/PblJmzSYgbVCaCBAjeHaRkox0DgHT9M7tA7J4Op9VrzyqDO0cb1O+zQV3Y7
Xf5uRt3UT+KJoZbOg77XXDisiDIb5WPMm5GXh8VFkSCKDSLIKmgTXsnnMWR8Zz14lIOQ7is6Z8Gq
Rz57mskTpeMdvUuOHJfQj28Cg5lAbgXbOPJ72lWrCDoqo4ZYL8k68DyPLdSWKc+Lhst9yfjS8/jz
JYRL0VHQ6kcbQuUqpGakhENMpeIB7kZRtCu6Exw1wJUsClEFIKFtgibZAFPqCyM1xm9GfZi9xmZP
FKJ4DmSsckPsKQwZ+Js6pbLFMmccwBGHE22ufu3GTavKdDcczYUOSEmVp4gzB7UdGAc9mYJjrPHL
dWI+0sZwhfXGGBwnH9VzvztqbUojWOO5d4D5Vb5htfS5WLWujTBMntXX/RlJwBdpJFPYgUFEF3GO
FueDKlf9UiPrILKUbICnR3uSHtlmcUmwRqHer7nv2R41mFQ849bnvyX+ERwKb1lXcrExuEnqLpb/
mo27ptDBPjrtzum4bUfdgU+qDcWC5ZBhvw6ilBIFFzeMLpbi4ywo1qHDRuwA5V5O53A269osVNUQ
XD7OlgRxZ2Zf5ldqUqdoA6xGQEeN3vumYT+n0WajjBKx6RHEdJSBnI9ev613RUNaXjV8Yq3IVYPM
qFH6DO4nwHUagbbjC0egTZl0RC0MJhwXLbKE1NV10RxFujtKSPQC9mA/hYuqli8zvOk7QrwfbYLI
d2Gq6DXoWSCCXXekqtOJu2+WDv1Hk6igYHsZ1vRxV15kZKF/CLzmtWNG7no3yekAtoPz+ctR1hFd
Wd3b5w/LOwE8ef2cRcpigsLUe45wYPPnLAUa81xkJQ0ckew1AoGpQPmUjpJBgVWn8wbj4/hAy5A/
3aQli4D75R4Xt5+f/rYIKY3q9JkDaWainRdlLDXa+jjIIL8h+Et4ISEF1S+vgpdFSUTAQz2eB50h
/ESFWtaslziQI6fETNp6IMLP93hgRnF5LK6Mgm5Dii5ox4zaWciyMpzr2QsOJm06SsFS77Leqj+6
yYDuYcgw3n6Ll3cBfxvizpoZ1U4ggtaTeeYqNKbWb0oP4LfjDSf1PT2cPzn0kHO7116iIyJ2RObu
4NNLe80hYSXcKbmKIi3USJRfocV/lPH51GGPx8lp7EHyT3yX2XZOK4sbRcOMSsS6KGMdwKSJChfd
Eae4065QJK02oeZowgF16nYg1mIowdeN+2dYPUL+jaX7MCnGS6i3hWG2Y3pxwRc2jbf/fxWCsKPw
wofhy3HbxqTGp12D29qaS+ENhNTYeMbZMAflwihpQZrG+L3OMjSD+C5UkjdzMtfMvSV+tt/g/B3c
RBWgJkEmtAjGHM7CE9hg902CZJ4hjYEnZdibYF1+T31BklWWe6lAMFLneBhoW6VjhcgJA5rBafgN
jySO4tsVfeBysciSYSLd1AAco/FpxTAnjLrG6CkFA9IK9MukJYVY3EnB91tfwMRFfnvymKt/HaLa
inr5+9qqN5aMRDoXIZys46LiXX5KMSGqOqpH0Yx29NxRvoIuFxwHLLYPHR93I5rF71g/OwnnHqyt
pErO/hoW8z6Hmr/Gzuovnqf4o3t31HHqpx59/Nw1l80jjVsE1xjPDx59wBerZy39kBEkogaUj61l
AvGE9mOyjPOhDcDsLGVe6FEu6gSzRZIi7BdRIB97AbJyEYwPbYNGMzINJfCJPIOlWdk5KTfxXP5E
O28EzsYfraIo5bifwPK6aIPwkxQRONtoNMEv/gcadrXCsnyH4TZCCUrXYpiaZeR5G3ycpNgtmWjR
AGIU4EdVps/04AprSBcX5UlVohUE5g94suLjYLmNfVi6wUac92WRX1/sFKwjKKUJEL3NhXYBVtKc
1FgHwDbn29D9wMapRONcMhH5jy9FD/B0BJF7PztE7yraycc1iv4P6StZnk8Ny4eVRkM4CYA0Pv4+
KtWabalVxkdcLnONEu3gqdjw0aEovKdqDV143jXSe2Mz6dsaMQvcy2xzLWnTwV0wsx/3CQeFtbMH
b6Z2NY5mueb/wBUp3V/A5XBS+2PTv6RZUEA6YnUE4Bz4381BjotkW/g3I0gzfk+o0RgCU4waiK1J
p7rhAgNXnoJwXTL2cN16nfNtj04VWEJ8XuFpB5sG9OJE7uT7cA/2CpNks11sO1/uNT3tSrmWlwh3
YZk3hp3y5JLW7HX3lOjmb+hgpUYEOawKGqd425F+CUp5Hc64luAbCUiyNSzwNpndOtB36fesl+cN
I55VNdNfdEwXtqCN+JWxPphqrQK7WlPCTW2aL74S/qGmCSURAFV9G6C+NnjjrlnjHFs4HVcEUdOI
s3fEEXfWrgpPFKB8U8gTRpcnLmxSJlggqzE0ItQY0w34qV/nnX4HWUnM4LXnommVsc4P1kZ6FwVw
OX5VQDP5yP7C3gXErpHJAmT0sX4TElzocziczlOqoNTqExZ9jR7epCuDC7EP85egsIX5fJ+YKtfe
5dnEfTWNiG828cCH4mPr6rYqL/Qy2j5iU9ZW5ADY+DbFi2DtASxk92SlQkiHhGpHz5kHaYoKxyeG
pYcLpXBqP4xIGz4CPDJ45kCh9QCjiWYQ2HR5vhPL4lle8QFXa1kLadj70zSNI3brd34fLl/UoX9m
w/QsB/DUFwnLK6bmjku9ctieg/0RERGixOuM+Rk8EkVM+ZrIUg5FlfQw3wpD2k8VTqB5518GyPOa
kpOqcPrvIB2TyEXYYPfPVjtyaTmDjWawtmeZqt7W6c+kRky3lzQOZa6lbercer6lTilg1Eyj0mpk
hFfGvSHArxBsbhvgoKyCNf03PyNAOxU32wX7zdryHoZykoXKfJU+do+T6XFSAxsOOPOWxzWkuBdY
6mvEGaCkeRfalDwN2N8bSFneev8RXx/ynEu89KlSKOFdRvPabF41t4IvAimpyIv7KvHRylr/G+UY
hLKvSffw0uSHJ2PKrOi3EiObNn0h93mck0oZ8/L1SetGlO/eMpLLxnZZ/sAFOGZ/PNgorjEJF0CO
hc4HJkrSUF1v7dEIPFo+aASrT+ZcYM0S6drRApqe9d3Qq9NrVLQCy+gu9+xXdqKBiRhJrY1r9wvD
fX7Qu0dreJMe5H+gd0h3YTR6bxLYcjfxQQCW5pQ3yjrfBSEWNPlOm18h/KzEhNFNIogo3eTzUbeP
b8dRY34i6vs/nLvhzEhHifZM2qdDQhMbbq+2AMrEUheOpZ6X9oIEBtFQprNDf2emAseDdoLLEpXi
u2YJ/W7azuvT83SFqlplr36V8p21/gUGGo6l7yaQg6PRDVTPi+p8gnaF1jsyf1T59OlkCxsJlddq
O5U7fSyheQqnFsgabR+EBv5+p/MzyDV67OaiegCjs9/VjMFXZFyw34GmegDSsAqEfHI7vxnrrQwN
zKX4jDRAejzSqFX+jAhULAGWjHWcn/dmS4JHYcF0x2+17FuO8qsm4lL7N+0PM/lX4XrQHJXT5x0Q
X1HXTRxfjpDsvrW3NNGLkUSrGxtxzZefFSfrKMSryuQOrU7h9JWZO6DspRAqSAvPQdollzthP2ul
GiAjqgaBh0NyvVUlwXPvsq2HLOd9d2HiWzHruelkMOzxderRCPkp9WmeUZtlAIfhklMAN/ObR4IZ
84Kw+/PfdCYXnfGcA7PilRnTqjfBgQER/O0/dcaJlknayoMPpfcccGCPgDqvWJYjYXf4QTgRhH33
S7Ys0UeJGDewpgO8Eo9y1BifXwfoBAKGVu04gheXb6zAaB46FPKM+0T4DTl6xl4h1zIQuO6aj8kg
Z4yOLbzRSSA9oI+GTd44lI8KGX4GaVmUziNAgrAQ39BUCwmSZd/fPQBSzXMfjET+nKrPAhn8SUOC
SciG5YU96LEQLKhXrVx8nOoyIJP+G7wE5UCHDMGKG2XB20JCxFVocli0MGbvPa/QTDE2H44js3/r
W45sVI+yCSnK2igQJbkOiA+khKTT1vh5xCC/oEt0ApnDepld9/8Wwe84I1+Vj//YYqz5FgxOCHLE
t19YgLD/O76UziT6oskiHBiM7KWr2G9bXNvgKofhzeIG71QlWGXyV1fnkiMJ1sBVaAuOi4Z1wfvW
C+Wssj6OKEE/5OwGphly+v23+qePZ6nw7uaACCXCdyHAvgzJiUGB+6c7vCS15XLl/r2glS6L7qO0
nnykfVOSCBj7fGPiQbfZ01YcyxDvC6OXM8cJ8HO67hxDcdF29efKZlmBXp7FNlYj7gM11xMKJOKW
t0hoy3xkF7fOvLmj6EVrxox05z0bVRQraHwF2UuYH7eVnScuPjsALpqoHQh/xPLGu4/VHKjzBYP5
DzN6b3t3BbLPNJ9/5sBzESjyhUCX+qzvBFMezXrtCwebZfFCygE+Z59lQ8loQ0yRv5W7y2iUPo73
jveOngb+9pEsWPKuYskU4Krv4Q6vO6LB/AU5+kEzmWH2U93h313gvvlSLPjBu2fo/PpGuhTr+D0F
ff+X86igm0nqVZuo6RXbn5VdIP6baEOzb4PY/pvplUCH5ByXZGtmEJr0Jl+qOEJHhoMlr6GimX1E
jL74//sVhrbPgMsbATlsNOEMgAZypnlj1g8lj8xyp3KejKZVpqnsqWxp3PSLPGe+npXnfPAz+O5L
G/yP19+QZWU98qKQzghvSxSzGPzR5VaioX0IVrtNyN3ZIJEnUucT9Ot9rH91Rm2zth3jgvrmGGFX
m4qb/FP57gTlnLfBhB5yyfa3oiY2JuMgNXBrNTSLi7fVRiELK51Q0bog1fBmRQfM923woBVsCtu5
l3Tk/BR7Q8sZI8JJfqthT9+GlyLbyy+OWJBffq4Lc1gtM48jLCA/72ezJvN9466SAdubc2RS/v7K
3sdXimEyccc5g+V3ALNH8P7H6AmvbL6WLSNgFKn1coLodcwWQjC2vEIza9K1zyiXl2bTXVkP2txH
F56Qa1bEKqKI31EDqpYNn+WvEcOh6jB6hnFJOcCxrFtjzg0F731KUi0g6YPjAaqKSMkmVBeEwaTg
F02hK3oo+jv7J7jngb+Ll8qb8C1fJyiwl4BIkPLQTPWlIowoGNBd5quhddrESVrcIvPB1rI49geM
TvfbL5Gb6qB5XalJdHFitbVdZkKxeMwF2xWrhhlzQXl3EX2XRjdvL0RQuOJNxLWJkW9/C9YpdLFu
LuvARClTJWZUBfxZw2HTQjdI8v51y3KBLkd8vg8KmUzh6KpJsuEF3XoCuPO2W3r+q02kTzhboqyr
C4umH9Q4ryBhdi79mFJSERf0iFETsTMlg7c1BX1QOpgZOTxwhDNx5PqkGzEL0oh0ftnqnsTiJGth
SNl6m2wDI6HaYIFwLgA5mi4uYlZWjA3bvNvDTxybs7KTXWsfbpRNwOVupNfa/L4BRRxirJwIJe6F
GDa9AFsVP+7XoUCOtS4636cNGJb5g/lDxLjdZMwn0WYpaULH7Y4EbF4omatC3zH/vwCV8sf3ECm4
hMZQB8DwgPYD8L/8Bzi2b3XVGK//TiXqg18gzSNuJTBj8gSPafwnolhL2UUh/YPqECvJPJ0rlZ/H
05USPsZS5g/E87ZExZ81e0+G+fs92ssH/o2tGxbjFa5exf6C6eFRI2uyMeZ2R5v35B9ZsHkxmQlD
mHPjylEcf4u1lkSpCRhp39raKbJARBqjmV/FwBZzcg/WE7BQMshsb+ZRk7qb1Pgfdo0fe35UiQAw
AG4hD9B5AaOkwhcR2Snde8zgh/I/vrTqU0wnwREcmwpJS2hPeah5NdCSD0H8TgwZB5HjYUCqoUUT
GBTktZxGRloOGQ8iLJFwdMRF/iQfiL9+usxr9Ric3IlR50p+m0zZZYpgX2XSUEQVzvbzuxiGV5zB
fO1LtxK7iMD7j/ub3zXIF4LG564eG0hfjNQLeyHBbunOcc8HTGnS38nWhSDDm5YpiAIpAX2ghwCS
6xYLWR4VolSi6v5zAabvw+boJmMXo8+3RrG9294v9coJkfXsAZH8aq7VDZd3FHDNQZeaLcI5/Sl8
NA+j4EmrmWxELKwZOA8Sq/nqgU9fxCgjbxjS2X3xiKSe3V8V3K6jm3Sbaz4Hz2SQGTh+LvmpB+25
os/vsRzgJNKD5g0rgHoiFOgSUQD3EL9cC/M8QxLKqa+HM7t6PaaMtwYDLpYkmlKmwcw4MSjDc3Or
MPOue4wt9KtSccNZAY/cTMwiFlvw6G5e2IrEbYqDitvn0GmeZ+k2rDTg7IpeEDCTf3qoDFxrIwzJ
Ayf2xn64xmjjXw5osIr728K8sDH4UBfePufpjfVf/P6uCuWVhSd5ajgjGHF3GQ81HCJNwpBD/3GB
rijSFq+5haBHrOarMn5riPiw4WoHB2GRXUwKQTlEOlpRewOBvUr07MFD5/sD1Ksfn/d6xNWOhoRE
briVO0V4aAQLHQSzBAcy3Tpp/ifsQAMVw/+97xWbHV/Hg9SzitT+KU256bDnImcG2MrqBDMQY55E
0L/Jn6MVWDt6AT1aMbWsZrqUR3YChk11Up6F5606plVzrxsMkpQIJ9wKfar6y5yWgFnPK0eHd3hr
p3bZ8DpaBFHhC4t4oD5HKq18A+AIi+4rqse/gQJxfJf87J5OfJGLoc7J9Kzm+CJaYCVJ0vukhnGY
BUHDr/cez4DnBfjUMqIjTmyEhJtMmNsF3MwG131x6SlpogmEgt0qFh7MCSIy9ta9meZS0xjoPO3Q
Hcc683NIT2vHf3u9AQPkbPxHAovRcfTZmTgZYkjwgSu2wkgZO6VBifDC3Yg7IMBRla5IGBJgkKQn
O/yKlkVZyjTwp39aWMLWXBWcIWfKT4z8ua9evpQBo9jfr+g0GVVpJuBmonZHCZ3kekicEcfHelOi
UJWaJDYlgrjSnjam+y/sd+t5NwM1G2LntJNGgBXrE+w3+BO9ee/y/8oCskz8AsKOj0PL7dFNlaYM
Glmjy5XrUvdoH9xMUB2oawoI7WsETPxrfEUioEwZS5crJcDbFadxfkPSeynahETaMiTGAlWmxtnQ
gsk1qLz6irnU1XDJSX/CGxWBQD8pjt4NEKysVgjfGibNZs+PgHo2+K8ulqDqbDiJ+Bx/RDOFI9Lb
+BS7lX8xIMr8/pmw03TWCc/xwveocqdwapXu8tIHsdGrpXcOcrkCtsTXwwIeW5/glcBF21JFBqW1
zWzZ251zfYWJhCW+RIxM0HBpByjTgLSdeHE9tY10Bv01Jcxx44aJ7YuKV4hNh6EC51xha5jL4xoZ
DhfEluoR63ITw2thN1YsP/hP171onnifgwhsrU3QKaGAy9NU57AZVru7j1/kVegWKhzjtTZAxF5K
vLuUkGb5i4O6aqjXsuCToZX8kVxYWqqjkoYyiYjuZMMtAsyHwLKPdyYhjDD4y9RIY7q0KZPBCHcd
ct6RWQx4Xv9lMez73Pw11t3+x2ULEnEprjBju8ZN7qoyZDqwbcPzSgRSOIhkDhm6j0FQlySPcZUq
TEgKcW9Z8HxV8AFLru8M/1cy5IuQ9JMl+7Tvp4xyqcP93lb1mQXE6DMOifHNG4w5FVZQ+KRDwG3U
5yqyopAcioeE5aorPW7m8f6sa+doLfOz7nBXoF2NMJ4/ECmRwAqOfgz1nph3d5idN0ez+0FBqknR
TvL8C5vPCARx5NBYiO1IoYlTgRy6uSIjyPCLjRH9Tyvsx6HXyGWrh1jVsVSRwhTAAjpo2Agb3plG
o/B6QpQyxjoixTd6EkWSIONqT5HtPgekOQZMoYkZGb/lARYe6luZQzU0i7YTIPukgEQNkAlf3o6s
NEe7i5216eqbs6WGaH8hXkjwDZnMEWalM+hFwBBZETkmOKMlbW75zlGgB4mNR6EkmTXWUkon3UeT
1aAhjiH3BSxGq6HyyvzcUoMqQIq7duydJQBap7gMUVVKA2dThVaejIUl+u0C45ikNMuXqmHg6Fza
CrdehqtvPCjCMnB+X46k02hUClUuIcpcPNoW+/DYJK4M6RnbiFIME6HlNTXTe8x4O94xwzdNDRkE
3hSfi+7wPMq4bAav9DczcMI5juqy2ZpnuO2iW3eixAXPH9vg3U9j+ua9HatuuMjKjHJOJ6ERtYse
Nv/UDAYNqEBcKLkJYA27OwsYG7ZdjEwOPawnd2JKnmqL3Nbd2xfgVRYgnErEvVhs539rRV/snRyu
p9PMPhHeaaKysinebKMBfEw2E3hmZpyirVNgmKuhwN5eAo0t0/nDgqcQiG6Gt7nhIngMvWXKKerx
UBsizQa9VFtsMAxkGcgp9Yiq8nt/LiPajEvWv9WvZggoLI6qly452FHf8kEnl7Q8XBVs0Rqs2MI5
ESYoh4u/EIXa7wIs7NWpX0J0G5nNLC6hvXP2qHDY1FIo9tGAU3TARUxH71oApM7hq8ER010IhCCc
uUkvCytqAU+7tbo5jm2PyjttbXbyJZF5F3ZgoWmLd9QWRHxXPCueLjRo1mBijrZseI2OjxJjuxCu
nllrHtWyOdakCV3311espkcChkcDA76Ol761RkaFPPTZ1LDH+DOJbyVH6vVwF21taDWvOO9s4Vfg
GjzfNJOWQ27RNFnEOYDSBMO0l3JSfqVswAT/KvSZI5K47LxZYfRD+rEed0dUuwRSU5CfPbiw48cl
hCjLcm8buknlY3Akm20TBpqIrk7Q6/52f3+dsMEwciimZ+0BS6H+1Jl4w0t3TM58O0MrJSSXZe4x
BP9syGIaCAL87xzKee7s8PGlWhVKfdkgrzeDOlRkj/8Zh58xyIG7VIjq1F9GJKDuoamZba2Wfajh
pjxQa/mu5adNzUOlLKPpMaRdYX7fXr+Zxjht3IS1+KZsOPgIYJzOeMJipqR3lPIERvUwT4p+MdBr
6G1trl20+8gktay7+8+bzFWAfBl0wbUfw2So2P3lVzrUe//Do1FJC3nBS806j4hkfnSOinujpJld
I7XAq8/6yh4n4Sk0bDhQ33TTrO48FqIzWgnWSNW87uh+xP6V/j4M/KqE/l/kjN+NpxePC9lSWhKl
j81/p8oVXspqbZczWNEuuBWFQMYJ/blDf19BfY7XDG5Hza2ajQXQIftPpHBCpYxuIBVdKnB+7kqG
IfID56PmB9hJFJOkUqyYML7il3m25Kg/2VVv9CaVy98z3zKEvjAiAM+HPaFxTZGH5JPyi6xVblUz
3s8OZTANEEwqjhmaV+AIx4u5ELCmLWObKkssGuspXS7mrdtLGfPPanwSgloFDIsn38j0gjrMMObr
oEzH5719kO3xMVNEnnfqJHa4EdMJEDLhW1K4K8pLyj1l/G8aUhfarQelQeZq9yN4JIGeYcxitWch
KcLApWX2tbF/+G3yCXV5NdxcSx2fRdDJFFMFG14UgAENIEhoq/22QhMfRaQwH53sWJkDReh380PZ
RLz4GJlo+LboBEd4MOASaelAJ/DVlqVgMHYQFwRysHR0XxSMQWoV5nn2qEZWU0cUbx4Di6c+pPxA
PtA7tZ6tJ4fHZyZs0qFhaW+Q5p3LflpnJNyfh/riynt32eINXgHlHx676zSB6/i/nKaGL0mOEmAb
iCtfp8mh1Ml+qB0X9OAsI8I4fVciESDCtOS79+RXWZrtmByDbSzUXttqdoEzhgCvyvyVpqX2D8wA
5R3ChCDO/pCY4QcVpP1ej7udPleCEuIb1J0WZ/wwssTPYUD0NQVK9SFLWl6EnEd42UiErWSoS/9i
W4pb1KLehWkCs5vM4hiUagJ/htSXN4V2IBH19CAZkLcAQt3tQncv/kOQ8UNhQ5FUTOyPe3NJ9WEG
1odwNTnJiHCh/NSlV53wkL7FFGnINcZzXe2BlyNASgKsE/Q3cTa3pK1yROhVE6eV247o1lhvhucM
4+kYLqVUHpmGLHzLhdFMvB02mHx2kJlsCqoi2uhy2uBmlFA/UD/Ppw6qb+ugSB1N5IdjBIfW9any
EPSMgpv7Nrym5vPn/E0wPd4PRkbbBHQ+ytpluIjVJACJvJdrctv1FjjRL5bWeBPp2VimS0JV+9u/
F/4EXt3jsQdo9vPJbp2xmM+/lpUqO0wYCJH9f157nhq1TVltSIAkxakgc/5bDJW6WyN2hHWba9Km
6XRVVNkmyotnaMvzrZoLrgreZ2VEAF/vF6n2+NE/Lj+AkVVxAMg1avWgDayx/JcyAj0SfmunUha0
m1bvnHjpSQCIaWBl473QXlBr+t3Vn4SsNmITzeeQzh5g0QVin1yso3mL+m3CVBX4CJgAMS6Xa6HF
wfvQBvOQzo5a/I5ZJmHEvYVyYunE9pg1nzBTmWwBJ/DOmor8xbOL6wllZ2eJUeqOS4wUCnYDOYOF
A2uR9nc1VckBu6f4Q9Ok5pmthVKT0Uik54WIscaJHcNAxHFr/WDfVWLUSPHbYmD+9SUzvnDOQH9b
qBPbDg6IWw3roi7UPc0lQZNlcmOS/I5F1Z68rV2UhNNh7EKKDRokTDT+CzyeXtmhwxeN7BCDGngc
EVKXcUcJiyVBnlvUd9UOYMcW9knUQty4JEwgFWqerbD5o8j7fSUJrWzzCxv59IvzHbej4WlNtctJ
ZfUTKFEGRC3H4+wIzJNaYyXnmsAHtmN1S3TImvNoZpkMCnFNd5OOSPhbvBH4jpl05IbCD/UwYBj5
Yy/LvQI++QyT9AVLOucKBMhLUw/8+urASbeGbapPtpNuRT4xls07mLTSY56OfzLWgsh7utFUWLOT
bUAgFP10GotCc6v9zql9Gvl1oC23xyv2DDmU4T0ewaRiKSF1JlBBrUV/uXNzUajoduScaG5617MX
yAORGSy7w8Nff58Fgc5CXl3YyDby0O5qLJcJKfNMSu2WFzn1zUg9DooLH0AWFRC55x64mpdK40Qs
sCjH0h1HIQHEmt1rDaJGIyfgKZHhMNDzqgFElDN/5RldHL+VvQ0RcgDw6lwPFffhqxLre73A1p1m
g9CDC/bTo8KzELom/WHJ6ecM8qc1pOtqhgczYsR5T2z/sc/zT2/h75XUCPAQLB1dVvzTjuwpNBFt
acTsl4z5EHaoKYYMcGEeTT8moVmdEzG8JQV1qKO2WNLpOBAWtn1BGnr9eRVO4qPVVdo5ZltoYF9q
BkmAy4m+2WxLgBhk5Gx13zFS5cPaZRQYrkqN77BXkjOCooELyepDSSXh+RvpKy7EcWCqVGPckHYH
nqzc/NElysf/IQDZqJIkVYss78eDHvVhTCRUXzkmMlzlIY10qaYsD5Q8gonHg+VMKJiEffDy5tPs
BG5HFeR68QmSu7WgOH90yRdowvTuKAkUEHHyZJeTR39hSEzI3djTYOLUfFqTd7rL1SfjRsa9keWq
HcQnBol2qz/ttVvMF3m4IoxyINzTeMnPwEjny1PPN0uNMBU3Zv600j/ORuu46Vl/ZLTuRiXH/P1F
pjxC1tyMoS/kX7X932ZrsuokWucfqo3y7juH3glw8kC5Cx9iHcz7m9BVQDNwxo3z+wCpd+F+mxM6
0CAA/84/crkjvlTxJwzOCf4JTiQLbAMwgk6RhfCMXmR7f5Xk3RSfizAbUgHxt4qTUBwA9uUdh+Pr
BqnEuHd+mCYxV05+aGeXAQn4RS0zJ6EmSeXNKQOBhEEjDnljfL5d6khV73mmNyazsWnCSaeTKxne
MaKY3dLAO+5s4aOrY9J2rDhSRWh+GE9E+GkooDwG6EIUt99j/naZixN4SCTtjCFKcnjvosjuqq8n
01Nm53EZodwvHUBwzT1+0BvP2f2soxyLFut2H4zbjEb01gHhngXYQ6MvIyWjKeXE/TuXy+RT1p2m
+OTTn9iOz8tiAwCzIP8wdOvObMnUKwqTGH9JFI2Mr1djh4+ImzpEXNFPEofkaGkVZN6uVcZ+5eF6
g0H96vGpHnvxVDdBJfUTd9XZb1Dg91JNu75u6GXpQiI38/akIVC3LKPJKAxS8OU4xtYtbTSxIood
gijBevKfvwIwujb7qoG1cA9A4AiF5dsp+Hl1tl41CC3E0AzGoAfE/bUDEapaPy2YRj75+UOqPk2E
VtkKBC2jPCsc+YNonYJjDohaMIn81FyI6P0FFQWKesJYSc3TQIskrAw37oKtVY/D8WaEZqMACTRm
YhgJYrzn7I2lc5FsKjxXrUplxZZlhqPqgKFpihG7eFmM5qbu4sH1+dbQoIQUjRmA9kPOnSSJJNgP
Wag7apLVXsSIeUB7NfKtvcakOv5DJVKnfiR8T/j44FALVB62yq62ZJTamJdvUlpnURUv4AcDTz4J
TT8kM5Wc4rgLLfLl85Dzm4qgiykvHI+FJJl1Rb+eC7VanLdPWY3oexhAqtwJ216jIqi3DTm/JaqB
DG45KGDG2nGDjTKFMiWbmKpeQu4ramxxZ1ZjYJSPiWe/PjoR5hnbPCrlvTfURs1hLehtRaYMjtlb
RIpMhy+4/cSK11gQQ/Km8hzavop2+bUiT+tUiOkXHZFZ8JjBnubaygfFwhfWRwYfydZTG3V8a1eH
TSKiN/pjXI394U3RxAemeaWU8UOD4+V6SsVHJS7SWlazdM+J4w5J8zv3sgMuwKUS0c0hJGV2avPS
eHsIMHeQbnzjbGWfa5EsPqJRDrPyCXr0NQR3L51DYX7arIf7LiK9sQWRJUt0vzY2eBMfRL5wyhvq
TTFOmbUwXnaCYZD8HptrCFCrFjnOPxPjwFebrhAtfOg85lfuNHzaVZWjU8tu5r/ZPd2NAN2V1jvN
WxTTDeExpKgJ+FybLSqs7FGtO6X+76gAhJHxVVjIb+cxhaz9JafH9yh/5XkVDNRW+dGQOCCGMKtJ
X6me0OVDleQrzWtvPXuePbJS/42Vw485kPDLkqHRI98Rcg2E8LabdDS6fystjKpPfZhNc4sYQCTI
5JT1YXDgu1FnD4ZTcaoB0GN9XbVHZmyft9lk1loEzhchAt3uTxnaNumhB2h58n4Z37+E39biDb3+
LZA76W75WBxKp0CWYZ9DpG/7//S4a9tJX1aujj/cqTEdgDe+12chX+oTDNvAsN0YcZ4XD0KJjrMb
kV1/R5rzc8wauNHJYsi2/eWLxxnxSxdzi+tUW+YiK+QDkkKkEHf3yd9nmgJ0LvmneLnwLLYxLONB
Q/k+QZQGrajndRZojEvADH1aM0sc5WVZegL3xTNkkyWk86CRpPH6osH+uTzzTbF9Uv2d3n6bHJ4g
cYMcuXmcZrfQHomPkxogYjogtSB1hsMwB+D09hfBQ4jGuNk+ZGicISYt4MtiNKzJt7ABt8cTN0ok
ZI4U/mXSHBKt1BX8xQeZkR1fdoIWH02b588XJHOfzEhQ6L//UJXZPn+UaCahqkKWCz+cticnaT0v
iXsbWhCtHNS7PwR8BV3om+Uu2qiRt0eQ2m8JiYtSbNHkkXdG801KJ0wWaXIrdhpKHQi9ElOB0BR0
Tal2Pjz/krWsSdfHvdcv2aGwLdvoestGLoMR/c2jDulLfeTEm+0iDurjeCGiAQrE0y4Pz4RALbmK
lr6uZZLupaiBzrYn71x+tg+R0MvwzHHd6O5Cpq5OwQF7Wb5SbtPUZSmZhoNL9rrYiJAL9sYUxf06
zvus3c/3B+JVF1wpm+k9rQwjMb3Wk8fUlGLoSY5Tc8eP15cHJdLn76pTURFPTe11priS36GMgw9t
tYze2WxZS4U1TLo6cYQTqa8y7YFFpUiwJrqyqd3AUDqJV17Zz9qypntoIMP9Zf6yRYPm/Ukql53k
1SK0xPKh2+F4NPijxjdUfmV1a3CExCcq/9AzDDXyR/p7Ccu1pd5WOFpnFkcoYilCZrpqEUwSzgsF
K+agp0gSVCt1G6JbJP3aZlP4rc/NblslAP2q1jtyZVf0OJyWWYqbd064NodTG/3YP6lDhX6i60Iu
MN5adqZp4Q/3qgdYdO1DN60bNlbCm/RASih7sSLTST7rpkWDYClP8vlyf/x14ofaH1toepWYR9/8
nXClvSFL7vGEVtk89yFBsTieF+6pdq0EBVNfVTP3KrOB7W+1ZJQpUXyqtvDtAWHr2HCJueRsWyDC
JBDjqalZY0BGWwBR52fhmYKsequAn04oKn7dq2bu6OL1GT6x0xp1QH//yIcJ0LR4RMslVscXcuG4
dhCa/L5oj1ZQWJ1oCD88+XZp8m3DbaI2+7P167pdjTagYKC5iuo7Hk6Le3KYnEZAOO5ePptW2HBK
IqW4xC6c7RgosuSOY+Ledl8imuAA3Zz+sgTZ6dTxXwdEQ8ZRL6XkYtyfrMHYAf9+BwWjTgyC5H8b
IwU1clG1+IZN40uJrx4QOFBAXiolIGk9Nrs6yU8EyFs1/tksl1P7m5XVrp0fPoIhjIzr8Ap1zs42
sbmvjUNTMLWytsTZU/ns/n/BIKQjX/twRsU9POk1C3mEpXqVQ51zJMqBxSUPAAsRGOT/PI1cLEQJ
xP9uRjfR8IbSkYyCMOUvAiRckJZF2/ZfInGwqFgH2fJ6r3wAJcWE1gn8x7k3RXETpym/JABz6YUe
nT5STJG06Vmm4hffLmcqR8kEXaHzCxDnY/EthitpuhQo7R6nsoR8GQinyQ4ksampTKKh9ZRIlLas
8tl1JBA+gv0y4sG8GVUu9TzVw2kyy3txOeo2UR6ZgWqA2S2QnAXcra4WXUdPV5I47R/3dmIrszoZ
Cg4CrhYQmLDtTvKsDVEsT4tl0Jlnx22496RtVSl6uldPcDlCwPSxgVrIJDgC6ZFePgVl9/MLKcR9
qncm3zmOonn+UDGKSGn7H6cooUProEpzYldz8uUuWXTdg09YndiUo5unpxgH6mS8R/+RE86aAk97
5Qk7pFx7cnLICrjUHfmutDnlADY+FDqu/7/sihLrsZ6NxVdMXJA6ZboEaw6Z36bohcBkrZcfS6t7
+nTXcXP/8UWhuaSpBEzs8N2wDYymcpy9jBontJPfgVdAe8J2edkqW4EPMIcw5W6a4tnZQ1McsPS2
LcR1S9EQaSsPBdU8y6wnVB6BwYcp86OjSW/SQLYSAYdv+lLC+0bG4/aQTpoEZxMvq3vxMslSm/RW
TDrvO7zQ9zroHtY19+J3tOIzHKim8iTUoTVLjTkPljV90mxcg2sSbbEP4C2riyBArA6qeExMLc6j
XJbKWxBhLZboZrTK1/TiUtgRVwR0qRKm9vA5/AyPWz2gpv9cApoiJ5C85Vfr6ecQr8mQWCJE4vGp
jGF3PVvCpYzDP29auUqrjXha3ZFJR6naEKScEWJ6RiRZpsIzTQ1mdek9g5tN+T7iZCtp2fL2cgqo
Q1z2rVtk+VE/MQxpUwk+UxzHsDQwfERJ8tVFRhSVk1L8pk00u+yLX7jgse8wHn5bdR0anowfEBXh
YsD6i+ZEiqktwCcWakIm5b5UGE9LkFkE8/WQI9qBH17aw0gKqO+7yRxv+2ySjMEWv15rCeYRVzCg
5VFI7R8VQhMD2fTdsxUsO+e0TuPxJ1nU4HSNoDH8Sxa2BaWe78mWf7ECmWjxiiyU4soSclGtlh/7
vnxNu/jArMnEo3ewsOytsKjTdjU/kugFhq4aF4MDerfDbS69OdnC3m9BTieIo4lXP4QVYoLlo9Gm
QO/sxiK32G+Q2IfQg2A6ISeKHgnBh3jMCdnhcnkYEQgQMtdORuttYCi3bp/w5MDOZG7uYmuh5BSQ
TpMdbmoh0rgak17LYolQQpRHgs8Gk3+pWx24mDQI1KBQhTW05YOYkKBUS2WmxocqnVKqRBu1Mc+C
b01GegChr/4d2CDd9XVHDwoUWAKANCMNtlRDOz7T4MsuTQYmIGsJAUjYJZEDemN4GLRsv53d0kuz
HH9uXXNX8otrruxH+Gu114ZmOTVlm2CbsaCJlgVs5R3jCfyq7BDRUL/ZF0+vo8bqaWmC4x0Agakh
uXFOE72qb0khndH8mLF07ihZ3vO5GAtl2fHrmefRKnbQ4GjDaYk+3b4Ub5YPHudkAbqjzxAvsKDz
88DJ9u4NFYwV5msUbgVnhi3WM82lEsz4DgS0882XXZZ6502mX1ypOl3lz77MCjy3Fr9UdQLuFVCd
tKBJII5JRdt5lF3O30A/wAQ9gYCYwkVLGUYI+T+mySWm6C1sEThyQSVICLZcaFFxHPOuZSvlJBRr
KXAFggAwg13mLn9KZZLlwqCgWziosAedI7cyL6/i2rsJeSHvuSZc7Ci/hUiHvpyhOEadxKUPcgez
g7tFWVrmOJpQN9Q9dGhOPPK1nJHiLNdSWyuq8W7YqhCJj1OqlsRirpqDaL1V2IVqXkM5nooEF4p6
Ssz/2Sh2p89X4B9+CIoTFxAW6hXStNG4hbqyrG4tTxq7S2RJO7GDOw2cVT2VuAFPLuL67M8pNUWo
KaCmTfp4vTWuPT9KoQEj6JO+1PCT88E2D8HybMYScWhOzHOErULC9MI8pCUcG3jMx3NRL+Hv6xJ+
8SEydqzoPB4JCjStCUR2Rh6ydpiuGQscOBNaAr5Z+VNT8OoH+XjmhOqV6g4NP/xTP0N76ZVjV77y
HsVbl1Zjlm4kHpzx11ZnExmNgJe3pSU96mLjr+L61YLN7YBXXgEE6WSxoeWjKc6FsGo1kG4gynhO
J2NmG9ABLvY0thVkFLsHTzaXz6EcuhAJInkjZ/F+JUh+EMSopr7rvm93pfCXK+1x78Ld4DAMHwf9
T2O7M0yyjJmlABDkihCrNPBPV1y7j4T1+TXAurSVXCBzpbKl5E/TvhdcvaIJvpUmLG0fIFsTNh98
b8NUzsZjj/VBddJQzZigNXq7PwH/g6zF3A5vHX4VRWeJ+z9CxBgMoc5WW1iA++5iLmXYbiKQeZGD
LuwfICpX0tErhO8LOFF2Gi+9/CCk0i6Ux9qczX+ixMwPzz2n7ZL27e4VSL2e8N44ORUvf9Ej70dQ
fIiWykNrbLGjFMBuKZEFvD3oZjpOmnMeLYgmLc81YHzpsqtOR630Au09eRrB+/FQZqUQuRSAQ79J
Hz5uM6gijwg60BJoX0cPSsmLvDI8ov0ZsKLx7DkzPils5Hn2Do7EG3QTD89jow0aa4egDC2nZhhn
oNSgT9pIlwdw/T6SzNg/lOyjpzXMthCb6x5byanEwd4Lyqtzguv+R4xh1ZMeDsbYX9PKbjUWFUVS
8xAVWpI6PaDqBfycBzAVQXq9UuTNW2WZK2/EBTf0sYr2ZmjeWf6T7il5VWm5hUK25DRqVww8mKio
hGxtA/OqpWgzRDk2Hu7Q4FCJT/XG6ataCB0vDKDCnfDmbUObcnSitPKCbus/A2qH0YFrb2ZrjASZ
Hk6En4iFkdXS70Tv7ZZTF3cyLP3o8gjx88oqHhM/VFGooMnMXYz2vLVJ/4BzIVNCAXzpj6xRW7qQ
IKBKM6SdlW4KKzcYkme3kgRlHo61/Y00r9QVA4asv5OclvTVh2zlh4LDQbGVxoloP8f4c2FnsVUq
dnSywPvYDPVY7KDt6G6DE5EkoNCO2YniA4k/NBuntMfNjsDrLgHwX5To9Fp5jZRNB/fAHDbqF1Qf
2HyCEA0X9g13jPhPFOevyyl1LvZJE/M+vk4PXGVjj/NNHsKvuvGnHCoJphe+EMZplmHcjmVwbeWe
hThL3AJeSbc0Phjr4lYzb7ElNSMROIJWBegoblsV/LKJZWe/XegmfFZkhb8pDrEO+GWdKUd9lcwV
3Tlg5AK7Omd8o0ups5gsdBG2EVX6PuhyiZwbtVr88IjAk0lFP8IWC6KdLSc5PFo/mQK/4OnDO8q9
eVMVq9BRRRM6nmzMpY/eBUZyWdRl8RGnRHVTUtRxKPORvjMFg6QQ2knxORaHCtXVUDUW9yxk6hLQ
xM5v2lnfAUtzpquE6PhGIZymeXGJSHVEY+lHRGs2kJrUDcRbcM3OfIL/yinPOexZ2sccFm8Syfdh
3EEQee25fXGtjoZ41L/apZ22ba7ZcBXOt3PE/jEEJbvdLyoip4K2ojNm9bMiaienNaJf8mGYDpfg
faktPtwLIPNBm2d+SyFYTvgeCvX/VaEns4YsJxzz/JdhIKUDZ2JroiiHZeUAvaGt1TZ5q6v+3FcT
o9jmva/LJV0ibY77wxNFJ7OqONp+A4uWtiCNce1CBPXfaaJsl+OpyozTU2ns5bAL6mRScha/veo+
6XUS29eoHQplfJrmcDXcHIqpU5Pv+jQ1K9NS+HhCikQLvJ0kOd6ofVbYBlCB9b+zlvkacLGt9bhC
fWe+IZp3gjL4Y4HNeEGjsFnx4a7U0R+MDz1DSe+VpqAd5DUOuabvz6gRCYVb7T4SFtpfuWpY8dyw
SbcdMbeP9JAf19KnFDs3XgOQrQqzwpUwrX2seOKTsUJuMIx9N7bs9lAt+Y20rY7BkOys7xRQvHtm
YUCy52A4XeBkLMeT0tGuuad/xVqGSfWLyoo561l0+Uq1JCFeQVbhF35vw9/IwyTsWOQP+MxzNKFD
qriWig0xQkz2p7Tq0SATjqtRpvKxjX8yLwxP4/+x2Qrsftyns6c08Hnpx4LoXAKUh/XUmPdeqXRT
kRdrqoPtQ3YDNRNAGrNqA/Hs0Phu6Z3V9YFCLomn95B17ispBqNTK5PxEHd9hlh/Qa/QaJ/uufm4
qgLLhUE0UOWrDDCsK8MfshiPrLCU9mxZZttqMkTjXG2UpRkyMSmhd3mKWv8YRKtF1TizFyDppnyd
sVzcmiOkVa/jQSOQKqMe9KOJso5ovDSSdcRDxtx3V1TApA0LSdoj9XZmTmleSW1ASF/5N4k/Cw7f
67zWyiIO2oCNBS8cAvpuG1CiMyZk/VcWz7KNsnlR7eZD5L3IUO2L5LDu22YWVv3cJJCDYBTyfldk
/d67iKbssPaNzVSlvtMYC3Q0W0aNGE7WnCTg2klXdRdlHlDwMUyV0DYOZY3UU4/avsLt+XOB91rF
M/cNd5xfFpgOyVu+NvqkVbDGR88eKd6wmvs8whTY3GLDjd5Qs8R9JqHQ+VWbYPuJgyWycMYrgXC5
LAE2Im5plXgoJmqWI0yJn9y3AAdymh54Ox5IUWFQMdUVG/5SIXxMj5N7xPGQOcnndpGWQblQVVJT
ONCSWiWGmqxqMlezayWUlRx/l7/XeiblbU8pWVas8f4NnW7fpZewQPPBDo1gK3EfylMJ8AzFfjOa
H2nohkH4iHifFa/0nfJWhM1zc6RrKebdMctuDf2zjcHXmxpPcn4oWesTFJbEtkZlHfqMZSxemAnK
FRbp/bEWr1PImgBAHR8Czb+3Li9+9dKFMKpATGDOrAEj0tmEGvc1vpK/mAWBaxYM5IDpktDHODxM
Pfvh/bCJZQsNIZq3jk3JFERep3VRWCekLIjWkT3SqBZTG5IJv8gSqrAbCSu2LPw6X1zcHA22Vki1
x0X+JfSLEoZbKLyF1jCIkIIkPlHhnnPUPmqG13CwrSEDxjqkdbRheoeGutNtkF0kjbjZdI5f7ybm
LWiaL3JhZKqVSruXxnih/y9Dn2Iua/CnalmZc4gYy3PqB1xVISP/lF0Ar1l6TAdStesKU708eZ44
2yp30Rs1yEAsmH8ABsFKZTV9oQIXipAdl+Qg7HYuN376x+cnmuEC0TEKkMys50wxktndjPiv1uk2
QoxQYoR+MB9VJJwZ/RiJRuwmuNSoBpcKyOtgTxDryNsT47C3gyWS8A7e+x2NV4o+t112uuNtzttZ
TF5AGi4ETT1rHzKTQx8glfjS3DxEHtALvqEJXJZbsgUhoTiUEqusVOgNmY+Gvf6tRz1FRGcQzS/d
dfDyllnin2nm82sCrDqAII9j83aWHXiE8kNhXpbsxqvffrEOCxjoshwRb0+arZXZrjMUWYgZlUbZ
FReNCl93lyKcRilhKnDoVc+ZlWsYGGq0WWAK340OAWAIjKtWUc46zls8fa1GLjNPnz4rEPTIsf7R
Kn8qv2us8eRDMLlSQ9zGdwBblTgZUGlcBOgc1z5tpUHuyeX1u0HIDIsUTExOUmWPjsVjcOkI6xKt
bjqd6Go3+oFMaPfCLjrvNT8279qnttC5W0URKU8Ueh30UduvnzpZcaLlA7z/Qwt0EC06pSG7eqrk
11C6epDSiQgLQlm0XlPFmJ+emHdReS6EEau9RkLMiod5W70gPf/iJL7P7H7qgFoXH0sKHY2Aqpbx
W9LoE8mGBt0ZNBIepr4IQTOJOza6wibK4upqDtjHZvm83Ut5HS+sDFZK32q/jzKo1h5N62xCp8U+
oh2hXtyFOECmmEcgjrKIjLrHBBGmxRH7zpv0GOmn8emxutjPHEcwdKMqadR8Cpjm/vmlhzm0krt0
7UASH/ofjfOHjViBivdW6KoiLQTfCz0LmCAA7C32zlb9wsmksThYQLFyDwKGoHsfUK6dpCB6KmRI
HZeKxQJzwIIogwuseZdOGUy84AdVuaQnk7yj9Hc5fwZsmPk3qtFov+XV9RHZR1RTqOlkKKxvew1F
Us6OqSAxqx5RE3r/6znKjMl8qFRgI5PasGOj729rdGTEU5gCia3beCKRrzwnhGdTuMdWLHLdrQQV
u83LVh76yk2HmsmXSDYjQN9H0DQL0UXaIxdVx/SDPxqiHZaSgXUICZ/5iE6Zcx94L/R1VBalGo4h
Hxju+puNJIXAjBELMr/IxOokeWTPUUjGLq6RgwiCgVo2e779ImyvaMPJ9coe228R9UjEK3yGPXWr
qo2eEIfzfVdAP1giDDGod8q6TQyCwCqaAjBB/wgmjCFyQoGXOJKI9kF4npwDhEoi/ySEmJHexE/n
PNQLugU+WRFA0sQPxON2BlrqSW1YJStMqVScwagNMzJEXDDB8ZaUciWLpMFmYSZ05pxXidz1L/iz
0LcgRmOKSUECKzQ5CE1DP/sKWsk4XgYWXBGHKp+VJZ7PTULm3hDrvG+IlC+B3t5FOxspKtjyS7Yu
it/JKO725E0sEKq3GNySHsWXgo27ocPagOHx91Rka8kbe96i8oZZ7tok3AaNNrpggilahX851ODE
id7Y0ETB6liNOTrkb9sw+BHnMKMMAd2ted4bDlmzKuvztgy/msSItohpMhKC3aLNjZ47hqVJ2AKU
Llu0icrtU2N58d1jn4AeGwyYL9fASWrdFbNuUSfTlyH6gjd+tfZJcFAT7sesKUiMXzfS1qxMewUs
l8mluywz76TE/FRjIzyco/2KeiBlvt8Ypf+sG47CKYdECampAKXLqFr8/ZGyLvG5vB2xwV2nNqwe
+bWGr5nrllXckJ3Fjkzhj1GLfTjJEqi83nXhH4fNyJ697zcVeNPkMCe1+rWCe6QW76dAvxoOWwJt
l0qYcThyDgB0/9Ode+Yn225NK4tlHa11eEJWBn0+JE4CyhvtkixLsznL5oHJIQX39EydcPWauiUq
yxnBGgdJVLj99vcDVRGUiBw0NnSbkEMPXi0yrBKXRxDJ5GyjTt34czyHsOV5ll49vh1eCAwNmMDj
GmFxbf9oH/nf/Nw1GFjY2ai04bAoYvsb10iZ5bqvaXed5RVBeNIpi2fU5eEzpcATPhO4uhQeO5et
NpyrhXJ3Ag305DCmRPbLxXm6mJff3ukiCSDaMT86wAQo4EdGIFv3aw14tlPSMYnfO9LTvRil2COW
l17V03epLwtYKZcWs1WL7bFxSiH2oSGuRfLUcpmwFhlYPadkzloWjvy1DbjEw+nzVhwADYQQ0NJE
Hq4cWeSO0JiFTYnpmrjBKO/TyLLOQcXmcRKsAShxGHDBChHjE+miFfS4E1DWX/LoIsHp4xehWBcB
kTj9Hd+JucuDIL5Dk/splJKUED+DYbK+dfHYAqXWxjKauso8xEJlVY1aeSdTBAD5zxs+k5TAc+Cb
n5jwtU608wluHNrf67zt/DLouyqbKpc9EZsuXrbI6M4nKwV34lptixgxws353W0boLxLBu+hIWcQ
eXqG3/Pun5B6uJjGffR1fZWdcsu5gDW9b+vDPFlsvAlRiL4Kn4YbG3KfnktT3Cs/HVyJoqJx8q8f
l1cVk5xWp4F/ZJfRXlPu7BB0ytDzldf40cUQNk3KIj+7+uDVCbhi7NXBcf8cRWrPLA0y53szGQo7
WM4lxN030unAGO0zXJS6zKmwgOQFw1PmOCS1pjicidrEFSLYRd3/SN9+bgO4ifw2w01uZm3VxEVt
ahkg+1CBZTFDD9jgvDKryjvIMFyOk8Tb9ASQlHUr31A9b1z3nHII6HMi38zKW/fci2a5LGq969uN
pPG7dospy5ZneJsbkJmnlwc0/LlLUfucBBa2qjz0X+rVk9AeUgGYt+f6Pq2GeIoqMB53utWruet2
PMI7AvG15Em7HY3KDYN/Yeeb0jiG5PbP/z1fNY1KTcHRMd0IZvfDkc0bMqjBCnTgMt0lYpEr7Acm
OI/XkI1W1/b2JkUn8Lof2uV8H9OBgUQ2NPhWNg6YBKY6wxXBZFsGUzDS6eTy5VPs+sw3/sCnpxx5
loPnVdxXXysXIPYgYt96tOoFSCbVl59ziROSI4bcxZ6uw/uuI6e7BPziJKQwtrz+c7yMfUZe9dMD
xYBCx2CLUlftWJ26GIAkmM3k7aRcqaUwtoD1kynFiXXeSKGA7YV1RYOGrXfyvUt/OskJrSDMw4Ky
QUEM11wdFbmsWcZon5rTYK6Y8HO7ZY8XL+UpnGXBwXi5WAeRCdeoQWz4gldPs7sssyDmtbq605W5
9hgmEVEypEOU2q8/3q3WyuIxRPdikqRlVm0nN1UapY3mWlyWZUqD3h0HiIueiAnFlWqFYveOo+Vf
nHcYZDNquX5c464V9B5jtD21KJoXUA81QhFmiXa3hsremrS3O0CStaIP1zWqSNNDXZKX1cbMzrN8
yMQEgWi0mFZjIm2mPlv9Cd3+fQYl8VqeWHib772i3Tr02f+hS9uUzDPVp+AzRXqHF2gx6psVa4R2
yzaWfoWCXr/yr+FXYxSm2sCgW0BbxmcdvfTIe12gvyDkGQkcUP084Ju49Ih04/TFq9bpjDtABPiZ
gMHq0wPohgrZBIhrJkx3Bqz/8FkMW50Drxo77NIsbjm2CnbCVDT+ez9nePyOtlZyJerdUOWigix7
ypNYZfjbfJSJ3/2Vr0gu/mIs79DIIpOFiztoD37c8wQhQiiu+/9EQV0OiqIFKyNRim2PaAoDznI1
ma8WtN12iiv06M0WgCN2eH5aNGd+fAwA7nuf6mqaXl7zET2TE8rJ0URdA6qtYf+HF+0Fbg8culLM
kpe7QCPPDZbH1KdhMdD6lOCe1L6qGWJTqeako3uqIJNEG2MlnIW13RJRQb+2j5uII2E3d8VQ5mEp
PfiifBqY/wDlQUBO1qskm9Qp6fsCi3O6uN7lfQ25iH2EX1D6jLqBR0iP/nddUd8p9lx6+jWrA/O2
KyvFmf75G/DyrxCbvUV/uIOh5kaMaMIqFfNJmDUl3oWFtFRodpc7R4wlASZpVXlyvxJfRD5S2Mu6
KVGBJsMHvgJjm0HoJ9zXhOPHRmZsBASNfHEpkeDb2fySGBt5HhvW6QM/TgA31X6ClcvfHnPWfpiV
U+1WtHdV4FEmTRd4UrXhUfAGFNFCqW32IKftXLo5GXdlvCY3IrOdYb+0U2MX5Vam6a2pGnhq6iCK
oQjmnkZq8MXGIaLlzKz3cgmC/fwAY9NuTrz0bfqE7u5tBFIaakH3wUzwMbxA75MujCvdK88lTyh4
AAgP7bOHJ8tQtPc10e3FfLbAurb3K23HLFxdxLzIFJGDhmDmU/jJfTr1kLyxkVZ4jmDG70oqJxJg
qZcg0DP2eqwp2e9p2JKIu/kgHeTuqyynR4fAS1FAtebILjHy0z8cgQNwPoJLcIv8QTiPo0nXYdQ3
Eu/e7YKczmMtwZvyHEWAvcLf5Ky2M9DBi0bKDz94YIRmcM8+b46heRrrmYaPGM0LYNi+ZEvGRH1T
VzCRD0SKqGT37Z4c2ZyLcjQTYyIXaONpVwAa1tTlaghK20rb/eUdxKWAKg6a9OR4lXmZHZ+ubzbK
E9NOQihldHod8OCq8rXHAO7aHhLxb3A9vhJs7zm/7AVJdm68CZyKg0viDnRrwXs4u3Bn7dKKl7Xn
vbvufn2eaoHRAlUxnkcWoiM0oc6KPR4QyhJXXaGyO2g+sclldUSFgErQ7D0PYgkzaqCUawxCrveh
LwKmJquhP1s50A6iNVeagcEjZSDGakLbIIXip6MrfOb4anP+H1Uo1HyAR9S0A/QqmxEU/AcOazr3
5F8V5khHIRmKrjqRCRXkocja3/XGHs5XpCjIRWUkCOuPdZIChgBgK7/xDAli9lMUSSzDUPBppLi5
7uEsbq/PYv0D1az5GWwxsJv46fG9weoPfFcAvo1Q7vaFqw1VtjvrGZgnildingVl3QMfUk+lR6LM
X00UJW9bbSWmTHZpfGAYMLL7wy2IxxD4+YOcGzI0Of7TZxVPWxE78ySLXzWEKtHBzbXqNu6/Oken
xMj7lwCeUV6zlWNgsMlHZXDwnKjHEDTiqR3Tx0DGX3xlvGWQU4ciRCpy+lxhlEDenbTGweZyMwMA
jbYt3PQzjYn5/o1zPyeizNaICfkBJ8UW0YXqTsFHQlFr16FjLqxdUFIFvzOUGHhYPft0Yaa7Bjsr
NZuQSfKK49PJZk8htq/nvUbCZaZW7oXMjUblcdPw/wPb8Hs03mJDu1AQMba4tYk2f91d+DRLH44b
tb3GbrN2ZOvBW9eKeBvMt+/5AnnYcllEz24ckz0DHXinpADn0uOk2Jq94A4w/OSB8NkSMgqUqkhA
Sbcap2f8nJHOVeBeNKBdOihc006qTv+LLypPXBN6zC9sYrZrULSsOgnkgsXly1m7J3iVN2VswxSA
luIi8DvkcNZOjETyuaeh23pA+OS89vRiyUN2Z+IsK4BztrHmcPaN6yGBcgojqMQlz0mhydcQRtI9
SqEVK3y62c88UXmlqlBM7aZ7lNJANNUmBIrAZXCxyPbK3SVQS16Bkrpe65Lfvj/D7VbMlIPzteYs
WmsmxLRqwS/xbuZTFnvp8v+7SH/H0Bm61u7jPxf/QN0bxrbONviu38OLCWEs0FYJ9jYFAH7Dc8Yw
02ucBex2Az2lR2HPyudbJ6e+TzMQ6r87Nzyw8s9LuxSEIS7KsoZEWP07YRe4uEEHhI1SfqkKYP88
VI0bWWESB/G5wm/RWbFUbgIsXsodxFu53IVODtquwGgD+YYr9v0ksJBS6d7K6rwBJmfOJ8DzjL5v
3lD2LH7h48kF2qFSFCXbUc/c72QsJ+MGJIR2LGJWorkeExGM3rY0EqoijFJ5OEdqkgEhwuUeRPN6
V0rmyETMkYCYXlQXFfGlKJ2ocNhP8cv2Tm1cME31LCuxOrCGOsEFKkZfvULVQp0bJZd3JX2BhCgT
FSjCekBVp4DjiQ6UQg4ypE2keNdgRz7IJJ6HPX/pBEWcibuMzVS7cGHqUfdhX0u5t9NvbnMytHe2
5zoKDLlBkSnjh8VSiHHnZvO6pEMyRMpeDct+GsSCTP3L25r5xxZu2U8RsBLAtPxM32siTtYbHvvE
Rpw8+HBfy1jUl2MK2S5erjLLJ9vMy6OqGIqX5fYEfrrbsRHA5VpAqzKZBhpgZSHCxnbtudNHMqVE
bUlq9Ya+FT1bCnYvqq/sFfRjSiokYP6WfM7AuviJu11Pow67nyDZ8CelK2fIXiamB+YIGEVBY/fw
T/5Cl/cba6Fqiar2bAr29zpUiS0RjXDGWhWTINf9wYsWFJ0MfYYY7WRz9c4V1e1EyifPNmbAUccj
S3+wQ5YN/U4YL+k96V4jQIHCxmg+H+0EfrOjIi7lI88i7EVfhjusptMX+e0g7vPiH1P58vyc4zvu
gRv+jb/3RvpUvyrNeZzQSEeqcSj0Xnp5/uWaFHv2GlYPhBk/H+Mox+0TCnQ7EZDFtBt3J+LMYIP2
pc+1KxNk3SXtxAPjmAn9KA9j9UZwYKVKq/Q3EKmPOJYVUdQJU9Bh7jy5S7UgT5WkAi4y0h6RCKgI
qO9fQMvVuNRTj2oXoP1bUCttpDrwfTTRHMWISFwXJ/BBM92BjEz2fB5VPD6MzGCHK/24dPxazJjE
DuvwHEOAMLT2KpLi4U7SlOLzBMUUG0ADVPRAaWtjpuX+Chl9OhpeAXlhEd6t7mgDtUn7JWCNkSZi
u+kbNPeF7OHqGA7nru9USOCahvm5yQTFmlIx02Dlh7vTk9WospiUJOHeX94ZTQfc7py/wT4cyr7F
wy5Im47V1g4eD8AuZHNVkRYL5NtlF/rC22qxTYGE6fVHH+tO2YlF8rkbFT6b1aLMQpauj+8IYcUr
j0UIy2Yjv+FjMPzNQkuOHq5nCUeqHJ6xm4sZ9nyvGB40vauQSBBbogjVRc27TwhZ59k0REMer/hA
Me1kmX+dgvhWnfeSQGjaHRPMSdqOd9IlQOYmL15GzHs1Niwh97xrBuBF7l1eVZKU9dAquHCzYZku
fjP2XMmbEnKHvU7AG05pZ2/z9GCexFDcMsXeH52+m2DaGOZopZq1wW0peXq4y5o39faqeZ6RBOlN
q40Ou2nRq9tN82ZRPzEFCQMyzHyiI0gY3x3rVCHowFYs+UX5tlxmRCAb/EyCQz13B199XFP2DExi
jjFLxesjhTyT8a/ZImqXpxQlR3qjfOftRRqjdvbbAtaRHLurMEgkEhffj9Or+ElOMwrdNiuBHmsJ
qypOOBqm5Vb9UiLRIQ+XRqHgEvJcvoGMEpqela4JM0lwbGtSSzvFR587SoQruq3yLb9aN5+ZMYII
YaBqkNmPTkicl86NETo9juJ3qhGpi8bIkoYJw440d2igLPbDt6WUNcXPJoWqcXJtV4s+iNSnAbL5
r9zXTSVcrvBSda2/S8uCobuS4SxiTiFoVsWvPl5R4UV7XM+tyG0INj+1En2Iqlu/4gGJQ/YrRsYR
6tG7+mTlIjX8HtHC4k8ksgUiUdFeNXb9WazblxgYKqsspsWgdcNNL8QDZAeZ0+A765QcK87ftzT6
fxi4uXcuUHihSYrPtGVIGdAiD/SvwJcMVtKgyQgKGOi73lS4awaCRy7QEAjTYL+pi/vnRFxvqz5v
5eV8HZp/cxoPcafhcBRoDXtsCSueMAenzBrnVxgBqoNFHxAuFywvXdoqaT8LeITdMu1R+XjNsKHD
8MOhNOerSEzP6OpOTzShqI9jSRY/9GN51A/CWyCQirE8hfBIs7Vb0BP75pZ6i3q8GlQDtbl2ArZ1
qhXfsxgrDOrshKKR2wC6IP7RNb78X+L+22W3gI8PGOrWU/pargMuBgwY0aPQVNAB/mNoWUm/rvvm
oMI2QATzK1ZUXL0Hk3wgjxlWHalq2DZapDa2sEOQJyYB0GX0LtkGU5LgPGwPGBCYO9UjfeNMN0Rv
3yMn/vJ9MpmYkPrxGHcDJWQ44+CKniQ236XVsCHaiSJq0TowdPgRRqUsLvJwGyGQVXtaqpqdSPHQ
k5m6dXm2dZG/ks+yF2RzAnPlQs47o8DuuzKtv5VVH4xLzeUCQQ2zdw1MRzTclsJW6nkFhWULiakS
tz6QnN6r4MTGOFE9HkXTOmNZe4qFFAp9DTOuAwtwbDbq/I3Rd8gC+y/eDDrnb96eyUvXrAlAACHa
q7HSAqOg8S7nIrVwqPsKK1omOnAy6lE74Om7vI3nA9EYQ5dlTp/2YI3swcTkbnKciHq1oafis1WW
c4cqgdHN/wVtXGZRa8joA+i+8ZVw0RRPm56prX/s4PIgS++tblh2bt5gDHy8qi7PCQRr/5/GA01I
wURaT4Zq8KAEouUr1thta4sJuJVyyf68yEYcsE5rn6Zlqt83/+PTkl24HobsZL3B4LZ7w9badSt2
QnmvvudQ1moL41+vmuTQHx9u9nmKHKxeW3HzqVuX+ZVaU2aTdDsjiWEMvhcbR75WBshrgNfHJ275
ucLu3LjvoIAM8FzvKriST/0NP60uZ8YnE7MovLDzbV33x6JLZih0GjdF9eIndgqReCExtLaa+JLo
6pSIq02TI5St09G5zJKKZTn+CVzLou9zM2YR0NvSurTWgsRkJR3i+oTA20QXSUX+HGgXiaUkB4+0
wojtyYiKK1jNOj2BIt4eLanJuTO1XYtLuwU/lGcYZlP9xAXQf4W5weTnj58h0oWXrvk6t2oh0KbS
ZBJDxZPlm0ansmJxr1V6Ydg5XaowKqZ2biu8eTKNTadSY50InpGMbIpHqe26TF6gF84adtQS2T7l
0OaKzf3SElW4J2QxtT6VqeG0DmLZrpc5b/iCWTWzixTNKzkHZTkaNmawy9lw06vqeZV5p+FaUNic
YmS3yEPyvBMGSRmbXB1DOMX0Xvrh6b/K2oYCsVzb1XCLlJypQFR2qzoI1vT6nRbjD+F5Rd2odh5M
4AX++pqeFVFPXOQ66lB0i984x1QIL0i0lKEWb0NiK1hqoYVIDx1OnTKNwQpGz+ULhaVRcCLvIGpN
5uI9F/ioKbO6wpQ42tdTIQvWT+a88vcxC8Jwhpcz9nki33YAx86qk7rsHRC7Rvq2tcMv/D6klhvV
EeVETca6CzcKsyLAfnkaLTiia7MViI1qklQwuQ8O3OQsH0fdqkxjjgAYSbB95BlvEjiawjoYA2ma
I2tYJjwsOvWqjAoxfBdJFRW2Kgegmen9dhNvzQOVHQJIZjz7iX+xvEYeDBmvKq4/bW6c568rdqRI
LZJPVutwEiyPJx6Z9PffdcnBXDq2RozmgHeZ6Pgy0mZTjNyoQpgzq+/stXeHE80sbqG2SbKZ09eo
qek3qfVEoWkSy2NBQUw3xsNdTyhPW+qB0CVf5RvbzV2QuwGcVBJcm1eZv8Bfiy5gjAK0DkjHtH/M
wNuHG7ffqzQXPThzrFYLGqMP9B8qKj6AmqNOgQ9bQ2uJlQf+DcbyzFV1h6yT0mAl4YjVYh2I3j37
4XkaZMlJuTzbqlo6lhHdsbQpkblT2zG2hGWtscjX3H0j0u6YTgLAFH1gk2BiHbFHmsilURpQvTJJ
rb8ZR+L0MwrHwzjCVLJI0TlA3VQIRPQJjyZhh5H9r/BNAYb++c7c9y0sLJCBREAGn8RRKJh+YVgI
9xJsvbykL2f+LcV3gTRqT2yTG4eJy/LnS16O46CycD7GiyTE1eErJIQ/JDWUvW7Do0HWxJrHh8Oe
vz3c31RKL5tQC7WDN69kFSpffaNF23BDPfX4ylnzCu8pYCP/buOnN+SOfKCXY2QjKmmLE9T4Hs3t
7OQNxKePrJi1Lw/IbIE92S/6/hA0bHS/+nKRub9OiUDWUH1gN+VfrfPwsUnld5RvD5P93Oc+3NLL
GrNStBh+608mi+Z/rZyPmaBk41BvX2IuZZrvdNDFDtcLkG3o8TbMZOMIdylhZOINc0I8fox3qNrZ
q7iksH2WTudL0y14yOnDX9lKJR7zs6W7/47iWwLXhSwWSSG2NJZNcPrCfd+YAuoQEdKlfBca20QD
0DoZqoGZjADHdHZpcJ8lw+dx4LHVF0ur8M9rl7hzsy5e5JVbHtVOX0avE8FZHjcAiKe6dXQr0u2G
7ApFkk2KyYKOF7m4czTG1McYVQxEIFayOhUMYUKhnFHOC3MH4c55HucRzduzFANSm2c/C9v/BhYt
DUYMNuRIxfeH4ilLvm+AanLDu0oNZmNUwED+2bMBOxPa51ap/lSgbYxPZ9deWhbmPuxCfkyNhJrz
HfiTRdWW3zTRhTD2MBNrYKgGshW7/laIw7/Zg9TefZL147+ZO2tuiVFq24/Mj7lbGKE/6s1GLYl8
vwcYoz5IzW2sYHQq3Dn1ODse+m0lKp7gmshy6QHezZQzt459L6XgwWDDJE7AQyCMWB3dUujEp5Py
ZRAwy1SpAK9w7ikhFeq77hscQom0jkvOWwQEPTkKo2ZkO2eF0MVx5LLrjy5+mSXffeMgk1d8HSMJ
LxJr/omltOAb2Bejc2jEc6pNy7P1FXd0Kai8oe1IRTccptD8/NgYFAsEYeqXVl6glIkWAM0Po8HN
8nIP7yX9tIPJFxldQsW2b1NB+ssDv2NfTa0EItsEnCFMNLgXimd1QQ9QSZZXe3K/MVsuFteUGy+T
A+iZ/n5UODQEAbJeD6RtV0jFehLll26fFI5eSw50BAuNNxVi+BQUdjw3EDJYAjnLN3u+NfBMTq6b
NNgo/BKwnhbkLJzOTHdxSIEWyNOvYwaVVnnQGL5bpAiyDskeU0TVuevoORGMqK+YP9m5SYLGhAUL
3tbaWaWq8spXl9jw+sgCNte5AJ6IcvUjFprbLecrWe1BHSt6ubpXQ2yLyaZ+S4orzLcWFrmRQwC0
qw0pDGHACSP9bzprdF05AYEZKeXq1pNxCjslBMYz5y2CQI00j30tNurokHamPp0x4gYcTffrImvS
DzD3DdgIoRgq19xd2q+XBav6IoyJUaleRT3P00ZZoxgZ41GXc/cDu0fGePMMtpAm+CumzZ8w3rwW
0TcaM8rmVbUitvQZDkEAFOvciaNbVbs4AjF8RBD9vdS2OTSNGC/oAFASiFaQ7tFrMrJF5dS/QkQG
TyllSa3ld8visi4BNFoo5bKLPk9Z4Zb9mXWgKlhjIh6e41s+PZQx6Ztt3uLvJpikPDldfLxi5dnM
IIBwko3LmF86FnmGplmFWYGvSx2rGj7X+sin8PbCmIt0PSJDadoMrGFypGllvjoqNOFEQVw5CV+i
edzbYB7ymfiT8AVXVWjEC0bwqQweqv6OwqrYDB+/7RFzkl98r7n5OpZizYhw0zVmEmkAJD2as1UD
2hI1ddSCjGVB+LHiw/EjSjDQx8fpqcHVWxSXMNE1gihcmDLCMVzv1tUVE7+fXKOp5MCDfEhQZpts
qW5YU/hFVLDc995/2HaRVBiPw97LTDixDVxJlTaPFxKhxPCWND3gw3RAieA28Iti5LGAbK24Me93
kDxSAb2mOXFNSyQlGxTCB5vukkR22Fa8r3ExwHrKa5jDZpxA2WU2IKu8J4qTMWtDgfsbSDC3B6i0
1OSlRcNGDxjqIz9DQC2kv07jnwConSdkv6NH/y8OeqFA2rEkDJrm55a7g8l2RdrqXKN6vxgzHmhe
WfjHWWVRqhh36VyV4TbrVuan8eVe9eg0YIBdvWhfmb8XfZgSUXoErc1kC/GcOokpA27GdMIh37PP
V8g1pAjYNwHABSKahdUnlJLaSw7wpyy/VyafEm7efEQUr+bnto+hL+HTiff8MHgKA377+aWks1gV
1+GQwZiIAC9Ort37Qvo5xujVgZLIvdIwnwzyaOURZOHVYxOMroIP6Z5JgKP94d0YsQDaOeEiCqvv
J4SpwVZtot414mA2RVZaFVqv0JwTkyVFKG0elaA++pFcWWGyjPf1yqNZ9MGpQDAk5p6yrGMT1flk
2XCud2kLRXBigkKHkECapkiXkZ0UN+AC78718Lnv+FNi8RcEhCSpKTSl5AjOhGpXdtGF7n3INshr
gebv+SbEIio3+pCxTKBAIpVo8R+6hM7/4ElgO/r0f93nA9aEryZjBS/WDTqTHft3WSJNoR6kLhWN
MTTmTbMu3D44Iy2vvlXVLpUHqORml391NW21ssHzqlEeiWlQtHvBQQDSSwo4GAxWxxUjJcuAupSX
8elsPaWCYbS9MDdK0CLh6VcgXqVvkNa3WtdLSJ4L6RaVyc2WcipgvGAENobynw2Z4qcgR84VPLiS
xlKTKsRB49XXCnMP25K9xAZq/zuq0wl1QTEh0QV/NAxbs+ftsZ4EzjgGw1eQIIsKJgX/g0JkkH8M
4sTp/JVG0YA6H6waWFukhFUDnhSRb/7w6UAPeIwD6vDqhDRr6q4a/UtxDuAJRppqxkZbm1MmO+w2
/shIzc4KIGf8hxq94O728T9ijIQ5nJRXYursfPjKKD4OL/Cd144ccZEUH0XBVEGpBQn1455sykFU
GdxYiTniQMXWi83JLYEbLuKIGlsxskBmUjKMZBn1WTVko+1z5ci3PQV6hklyT5zI0om8rV7+1VnR
bHuNa35Qu6fP8sZ3Rhsa3lcZazk6mZ3EfnwFhs5v+zxKcKu219GCwIiU3kGsmq35qsWQmPqE96rl
rQmHDIifeiihOXmvLcHbQ3OlCNyUNEIivD5FCx5cWV5idSNnpJhpEQ6ebvWd+tBZ4OeLBq8DcEGW
zFQb9WdD7WqfHM+49YVwlKejM4+wCwOGqDUVC/X+/R0fj9el6ZXP1shvX88HcGsvxmHp75yJslqM
iD/nZlBtb9sDdxQFTQNb3OtJpvWklBKuuoMaxF7G2aGWWfn/g3T5dxihkNWhObpnwXxIa5LYQSMK
39/IYStKKkdW10k/OzXaMc5tkStV1dpPy/qHK3rB/LcGqMV9t3lUdLSy8NCYaCog3mO3mWgdBJBF
GZECcK39G8VYO8JrRLwO4zmLaiXGRuxwGI3XPaHE0Z8EUaMHF+suia/GbjEPg4vKJ3yKD7+zVWDH
dhapDs4ZOR1TrUc/3cHtjgmxLRxSsibJFBWAvXhwKHmqp95Bg0pjVS+5Jm+FOIZdyxzbKBgjpOyJ
Y19Z4IK6QI7tBeVVKh/w5EhXwoE02J1y/tl442+6oPc19go3lDOfEF+5ZwrP4xHtAFc+woinIZAq
osxzAEx+MNIQO6zk/QWUNdOvYp9sPeIKQLykpou4YFTIz94gfur7Z5+BD+r54Cp2A84a7v30aSML
dvsleLjvdf+BQdQ8itkF9bnHbQKGUuGaX5N/cx4niGFU9H+qk2ZtP0rhQ+I7H5ZajxWX9tEMzaSp
ctrLxMFrpyKkzAe23wKhD0W49nWMO2t9KwXLkmZJzTWNEGBcBwuWdwzklwRZJr6MqGCSXGVN1F97
KNo4wSYkkyEEqNY0cE/tED/K3w35RzJT9sW/f5Oa76Qc6teio7ieu32TzmvlZz7IZKnOW3zB3lOG
LWwOIvV53wVAB1WtZxzyh3A15KR9m3d2mEWDZ8hyIkKnTyxOs4Q0YOaLT+AQ0Wsdq5+ZeHoTur7d
1d4ZLOWyJ/0GURvBYKYH+w1ok7Plhszmuy+g14y46HcygjxlnBE5btvsQLMU0mWF4ThLHFjoVaH2
osbNFMlrrQF8P6tOrQ/531PMEuUAIuhqppT1EpyI3xOyO519u6lrHEa3K7EbYG/iQaVso/TIGg4T
1GwGHc56CM6UwkDxSPNKIETticvPzgbzS3WdPyYHd4ueCix0nErg63h9KhWaH5sVxoxRGafZvPYT
6GU91Gef9BOV76NHn+1OSRKKOoXML8xUDDFemldxAEczlSG0bqcNKfLrSe/ftzF59ha/BUf/FpgJ
UbN/AvTDA+i0m/TIrAQK/ydUALzjVe31nFnsFij0TMK5Pknclg6YDbwJqLvpD4DBqVktkRYFZn90
TEgJ08vTyul/nO1f+5bNr+GWLA29ahJOEn4EWooyBAT2V/hyIoiusIntTW+fc4mnkp2Y8iaVdkAm
pCaleEyEuIOPHd2uNLgAeBm+nBMg6pAUJWuQu455JQUzXTKd949KLJopz6QffLuvrvlhvPix+7DV
65vloNFaHUsFtORf0Wgv55vd5GxgrQJPOwmRMs17v0VeB+8eoTfX5KXtuTDlPfCtTfZYBf77rZdW
aX7gWiqf95f9ZaQ82Q6xd1/7oR1JH4kXydEcUjmNavzm5MyZU5CSKgj97OgCFh4seO1g7wtJRhsF
jCZ9v2a8GsCwVy65s1uI02zQYllT0YNXWzno3bTFQOpYintV+SblMG2qrxVdq3rfTtItm9dwNcO+
fhR3Sf2uXOqMBZ+0SZwNx4JvIlNUg1DEsBzL9WOBIws+EUUduUmjUd2kOQ8CyJS1eArLGc1uS5t4
qSSX1zHCs5qgddjZp5kAwp28i3grr6R8MPSMbz9590REMICIEUZMLKZVLdo2xlh85xARMv+UkTi3
afTcM6DyNF9B+V3uLO06GTsArls+uQxWiYSQuyQBTaTo9+VJ9BQA675q6Nb1c0cODM5f0rH7H11H
U2OD6uNr7NQvHaRzP6RljASftu2YskWsu+zIrwylMvInrXAt4CmOZNylrj/cqA5zZSs/NWVavFfP
t9wufIBLWEr6cvKklydZPyM9M24hgwjvkF+paeZCPfKOYwM2IKego0xiwUZ59SsQTQ1bwakjBlY6
p6BnTwMaVQjr/1yfqArydBOMTFmDao6J2FSS3cpQWR0I8xpU6K6LZjOIykxM37tQiGH2JYMDWGMp
8zLDQl0yaCU/qWkWxoGgKwACV+jVvEHE3SPdapr9QQVQ9ZRg3234eh0SEWfVg+qn6SO+0YhjqbYo
t7L0NPesJWmRdHfWuf+70VCtooqgmPz/QQxEKe9Vwc9qbJ8QSHLH+5gB1Uj/SR42CfLcxBMfG0Q6
xrSgg2LgD5Pwdv/9K8+khN6LDi0/rxI+ENli3KWTnm32YGugLdbXJkEZFXnCgR1q1y8byc5Ewk/E
N/LzHbaXoBoGD2H7wks8YehIOQxI7v2ineSDKCxJ5/rVwtinibVePc8XuSBph7IhvMnA0GBSeIJ8
YAF6yKrEv7X1rCiuoboIwJLf2mtWucCNXwMv1eZ8b+uvsR/GRLUT1KK8+2kT/vDCAoAysajCDR0y
5LdHQ1gbPsTFVtEpOhKBA8FolQ/zPPZLk5HVIa2kMd+Xu3vRqYkWoPqka+aAROlM0r5bHFFJSlpp
b3gAKMz5LyFXq3eYYrWDctXJ0D9Eo13U8GjgK36L9qWnI6KOWO5+fdi2Kg2YOy8iak1IuJ3BMC09
GBWWipQUOJWv59JY9E0eht8NLa0cGKdksJF7GCO0plHgnIIs8PaUKfgkhCdKThSyz2GIwr4A16uS
hY8qmZG+oah9JfGB7JVMszcKfeDw5vMG19RMLU4XCx+ofCCtCA0KXiiYxY48XrmdtxySXLGuQxmI
hsEDfLa5aHsXE3QqiKpK1nmp/HOnzrTpCZ2eEkqQ0UoSc4Ys7XvMa+MxUu/AojbLanF3aC2dZN0I
FLFXAEqun584YwPoltgchZQfC14sU2CULyfEmmkC6duPvY4gHZS+hSfbrK914CFafi8Jsg6PeHfs
nAVezi3wESqB5/D65Y+JFkgU3ibfnDbAbxfzeiVmQ2IWEVL/Faql1bn4g7qCXk1NUBAcAhKWRUai
JsieaigK6rwo5He/y+vg2hmQgKsyMdr34Hgo228MMUgWolDJPmiWNLl54qQUUJCSWmqyLZu2L+NU
R0CkKyVtQPVzDxzE9CrmSfbyRkMVSCqMe1PNNVm4DZ7yEjVLZSqfDMnrAEVOgvsvcHuBARYoZYCl
5b2f1O4LCqdDSzNM3ZSCgv8CdK1y+23P2K0/otTNn85me0tVpuDVSCCR3l8ro6H0kbDwMulDn19x
KdOfhR//WgVCqCMq+R71JjCq/mL2FybgMkjCVNidizLydnT5Sw9IXndWc/t5As+ND89cCu6ntLne
kIpgiyDE3EUUkIXkQG6SZQxlY1kJ5DLKLV/2LPo0aQhiPC3onS8fXiBbiKeMHP9NA8Jhdw5EIqFQ
0sKgVnQkF1xXMG95fozx7LFWGtQsVZhuCKF9SA/vY+rG2R0q+ad1oYtC51vFGEdcYmP07QL7K9Zk
PbOGtmKYO6+TsHQ+nzpWYrQizUcJdVUK9maIpZUKA7V3s2w2TVNmuKRYKjSm9gCjGTiytV5mu5K1
OGKkj/0dvfgpVFIKG5Ce9BdB7GPBMxtNnEFLQ1FXzbkoU/esv+WCWiJ1rddzGQlRJAPP8KYHimEw
Vnq0e4+8BLpAZBmKcVFbk39HqU/XUJXrQn4yxeYm+LcFfYi/sxFBT4LBusjXBDyKeQnsG9Fu7RUU
1htRUaMYLQsrlMfxE7vbivzmHvojptjAC5b1w5iDDK3IiI/owEO/zWBhTNHhOhqAFNH3aryUme5L
cmOnTK1KFnsU/B5TKO+4RM7oi0Sy+s87PMr9nS1S3TDNp4P4s4LOonWy0NGL1+rY5n3affk0cv3w
g7N9WD7eNzBjXjnWKV3gkG2jX9oglibrmtIC+thbGMdH7Sn3J2af+3HAVFYkfpsqakt+PxdMIU/x
I8NN00FBDtCMm6HPP6imoO3ZfQSv4erz6m6xOmmhxIH1OS8cpIN1Ch6lrMVO6biJnkVDT1395jBg
1VCjTJCk3iVcxV37e+6yxphQD2J5PO+qpZieaHTxB+VbXfD3T+AEITQxZbGOn8qEMLBgOqpDDeT+
JMTpE9tMKW/DJPNoX9oJcatKzk+Rbv2PrUXOeEfGmb0mGP/mtY+Rrqcnb0RigVmUkDFFi7SHErZ+
hyP4ip90VCAUl3P0fbB/BuEgmmuMqvWRKnSFQBOKW0GE8yKeMjnuRCdggQPgXwXsVpzNp25PUFXT
gL2/jui4D6ele6oe599WAWdTRKjMjDgDXi2do0LE9Bbio4BmZ31bagOA3S4vX6JpZlFn63bAOwMH
VefGVyrxiDlDQlm1HqQF2TheWfFdg3DpYl1nHC8OyMivnfGbhXbXanL1TDfXhYbRL7PykvqolWU2
PnZJssPTZ6mXwUAe7SZLGRK3Ce7TR201lUKUBq0ej/sAsnjizRxySF4uHrbJpTwYHc35d9C3/ryI
uHHPa3WjYMYoRIT+6/sB9dv1G2BUm6bYQqhSg5IpUbanK1nz8kkxivD8G/fpCj1xBuli/P2U18Ya
yoV3wmCTVBXUEWOM4hcfsQewwUpjThPbbAe8lCxElsPpECZVKnarATMTg+yItLkfQI4HzKMSgrfT
Y7GZyt+3n21CIkSHrCb5w0sBhFTPwP6FXhJcJ7nS5ci/Klzg6/mQsJ4A0NkoU8Gu2Q9G2/Tog/A5
PlBIJsZDXMr+fM8MSk9UFt/yW2XdHDsDDw9R7K5O+gl2tDa1+82IfHFavc0tHuPAgZucB52MKxT6
sUKkZs3xBJ5dPnHfHAF3mQ4lvjJZw6zMFVY7OfBw43QCrtOE3yeMy/pPwVwSR7dhzt3+lqptbujI
srLvhZgdQZHoB8y46vmb2JbRYY/NfSEC5+ndHomrfz7jCJvs/C50VBuGZS03bcP8vxn3l4Dn/3en
mTYlaYtFP9Mx9MPw0QP7Tr47zSjtpHRL9KFcNra8fA1YvG8pKPH5FjEZahn/s9XjDz9BJ1BHYMa6
IdDZwzkHwmbzVD1E4PyihoIGs8Jbjg0RwiLTqJjd6NDHQiZS04QqB8sb6gLSjK9gsnFSumlQ2n3r
xb/7pZLxf5xvUZxXhScQcVUvgH9gkYExQVmkUuq0VsV/52J3CQ7DSiSFr/kUxxip1ZFvXZixPa3+
cERprIzBCMmGdbL7av0W+SjCCMkUMlTesvkf60e5HFaovli7Zsk7QcdWTRkLbKpLCQSkiMlkytJ2
baSLzE8HVTguozt00qRwCeIgD+biM+m0yV/AAe9MM6WMUuNoIEc3896VxpiNG5ug1SgCy7lcS5lA
PbZZlgm31uYDWuR1swUIjzfi9OPcmMWfHDL5pfY5TiEgLCjAmjjLxp/YU3MTu0IC7n2bb4fnKnDc
04Gre1Uvv/FqX/eouaz9kyuxHOEl1AXh3e80eudATmE+BjBFoZRzfMjOH3JS9bFHbp1X623Puyu5
oI7MYFsSRjdG6nraKxK6i8woWXoPGsbjCTTmdYRaVaGb/u2btZA8AK4O8zw3pUi40OaGyz3id56r
4D68JR5DDoz8v1YdEEbmG8ZOVrgOpjulyL+IZaR0Z+Z/J5MpZAFlQZZKTRKAjPtryfDXrvyWA4kw
pO57dMegHCh9ayZR87jSyGMRE+eOfoi/8wMZO6e8qmLxjPQ6p4vGeX1eRdV9oU/jQHaVfToqahtv
ZtE0htwpYVSDUTLSDwJOYQ085FoKiMgAMYYJpbWsl81UBgvziyf44ZJzl870gzZxK5yVNdjVKinI
EWHIhJsRQx00jS+YoRZZ4CGZbbL6lup7C6i809ElCSTofpG6tpnKL2xr3dgOqPUeAA8YFt1L4fyl
PeG3vVSvhm+bSsjUoyBoMo7e3yQJ0OGmsdvHwtdyUyVSNfuo8OV3cY97QDM3QIvoM8ueKJzsCyEI
ZGepxRnAHVB0Bc9oVNStHsLa3NShz88JwG4QPnQInINa20Nzoe+fbJ2jWMTfGVzkQws/WN2C48AH
RS2VIk8PQ3mM/oKSfeEExzgOnu6PUjQL8vU6BdmyYXBbuJF9Vdw5sq06HC2mVZxO+c8rDcKpRXhP
k6rSJRD1BF3nygiLQ0upxlteZQdq/nllHcbDrdumdhUIxDlq0F7NfsKZEH7Xse7E1sEMHOk0eLAl
qF8kpfTEJM34YLnz7TCRfCC8f3A4YQD0yekO8dxSOIKr9ZRyJtg7rg1AtTbB4RWtQa6dnzKdg6vg
ZfbEQHidoCFlHPAPh15oSufGodUq/3c64aigH6RBPW04/yNJ0qgby4N02Nn78PAzsXbuDKi4cR4z
izjUlMOo5gVX5q3W1B1VxYl/fsi/jLkldhfDkZZtkwjt7tR0S/tmJ+1BOMbcZrYhSlAH4kHaKiV9
ht4tzs4LbOTQyJG+sMBh66FQZDJUtzKiOGlXt6Es7EjvCQEEMrl4M5YRblOwi1Tv9/2UtJ+Qh6GH
xdnEE1kpjzJfBsft3oanK8bmZjIecktTdbGnJ55tSzB+a5nLtQoJIaxkbjqCkQo6oYMJTBADljfN
NDEQgDkhBeLlv9ycfg1LNPoeUbok5l2IZb0SsJcoU2NPiryfAC7xKZ28W/kJ8nuVnk/7Ka97EpeY
HMpo6KG+KRLvcTe/hTcAXPc9ZTB3AsTb61Vcy1bMuuxLiVRgMz5G3MwthgmsdLGVIW1yQN+hOOUo
qaxP18cTuvfTl1nIThyJU4t22Yn8BNq4by0Cz2K9OWFx+3vYbt1qIX3M/yyJKCZZeIms+A2FWDKD
xmbCBxNp8zkIllbgDKJB6P/ISSs9WUPubNJ855P9T7H1AqwK432mtG7n8L0CXzA3TNNOj464AMIM
XPkjgadFOorOAmOPCPp+S5+YGJOFhQWUcRB9iDFk3yFsLyBjUkNR7Gu9TN3I5XFkL5a9JQBzvVgo
3X+8seqys+5D+AQbLp2+3lyJrir4QeZvHRN/vgwxay5+ezfWklI8dld1K9q2vTDja033/dWLlZDz
MosrvKz4j9+UApFyHz7VbUetn/3D/skdyMkX6DK+dD1dnhbLSkgsYtVu4p2LMD1A+bDg+iQjnFVw
92KM6WPVJAjxFVZ1TsMDTw1tm16FixXfoKPNsgj1yRNveXZe1XQzah0jc2dkFqr4uyDMSNvciwvx
THMWyaswzUZd/l8fbMWsVx4y2JDAIVgCmq6rqYone0zKqBpn9vMIDee52BJVJXFhRMX1JNshU3Py
KA+KYwqJe3Nhg1Tci6126ObvSP/e6sgNC0lWSLsolGxBzRmrRHXMKg8Gl55iQh66taPpX4NA6EX+
zh4MWGg7Q2P6gPNQJtYs7UnJwBwbe+M4uBFf62ugkvyjmwB6LHR9GmRiDa0TJ7Unt7qAFx5FqQEm
60nX90+RfYL2J41U0kHbDkrn45n5YGOZcIK/vWEKVqqKOGInNevo5lhery3eSYPCygtCHrspFyss
MXwXiakabkyrQWOaZDaKfxhKpAVyjfWEnLFSG6flI+TfwTfchKKUJds41Pa/5ezRGGcOSswm8A9C
00CZOEt8GRxyioWIQ7o4u80Sk9JjVI3mroeJMCMUCDsMFqbiwDyVld82Eznw7en9lv6qQCJea4FO
jSo9TSlefixV4nNsqBr/iHrUDVAIVe3TXzZFDdzQ+nrTEjiPUMeEUQWTC2bhhoZ4uLEI+BtinRyp
sMJN5E4ptzapSXB3wi1OJY5fUWC/UPlbthSoT1LzywZ/Jt8lyHra3efkt/foAKSYK2O+f7d99xeX
AspvgYOG626NLh9sEUhYOWCQSdcmNH3Xh0SEIHJDKXDCUGW0PbTE1WJWWqEHfIBX8okv1yf5jAIR
nYJZHj6M5OfLfeVh0FbEnoLU9gOb/B86lHFytr22dNL9Fjl6DUzfe6aCoObcA7lV4nljcsSe0rnc
WvXQR0PHGUNVulMFy8RIOgNEAWVsXWxTiMuqriLlQkzhydupxPX8B/BKMxxgBDu99ar/twp5Ex9o
3lnQ4vfmI1kYjCx4yK9vX/MMdr/fJ4ZgtFcNgDIQSQj74crnVPocSikoECJVTW6WzYH+xLA3o92d
Dhh23fFhFxF7bEddla7+pIwCRcNCU4vtJEqubUR1DYzsiZ6oocy7hrbGsEAHsyr4lUnaZrKau+IY
aIpCx7DhKQKWxNyY/PLYtEkilJVscEsJHkiwp1yQw5JYRVqLi5trnzWWg0hAc2qWXv+GTYxHP7iR
ZsfQx4gJuqO/+PxhwyDu7hYXsaGg4PVOXI0aJ34yov9wW76t6c570Jy8NXtjfZqG0wpfS+uDyaVD
d9txCreTBHclanoYUMMuREGgHlMu3QfwHDV+qtae1aVCNtcS7ki2KM+/2HDFt3J5DyuNjuMph7Pf
zNhUtmuGcnt6dVITkTsru/IkRrPTy6VnKEyLpY5q5+GWbP+VzPKWGpZJeEsJZbE538Wa2JH+4WLT
VbenfZSHrMq+Wjq9fyOhWbQ3aknzEBHF4vLzEvGNRoFZHJFcl4dvjqbwdu6jpzaWuPND8qlMN5nx
z/H9buLxpgPVbSe9pkgfVFgG8HS2XT0gTx/blR8PYxZVxDaHKACWFpjTRTffxroh+EA8/eaYHBem
i50EV43irvocxwBaDaph1fs5Zfy0kJxH3va4KM7tsrxy9Hu5FdIgEovQZLn7sXl8WRmhjUTmeyaO
PnGeib3qV8BUbaTYjTX634TWq3f8fLcIG3NSoIMe+iTBUx3lPC1g+y11sPq2bafBp84mqS0V7AnG
lO2rOcmILWmXmOKK2ezLo9WVmbd62I0Gy4Q+e/dpPfvdP4E7qotrq2LY+14B6vnWArh/a51bRbZM
uz9Wh2v33s/jEX1MtwPopg917iPQAVDfHot4QVumbRmD0ijaZQxJXYgo45H/9qaVfoqmdXqW1FQA
RKvnnSznhQZwIjZwLB33SvDSp5+YPBbTVRC3ACcPvQE8VXI04hMO8ELtohxlNPoy+yp1FyLJiuev
rc1TW7w0LwXJRMYvVfkK8FLPLUxdj33wB8bWB0h0m8JjgTS6VlcsZPUE2xbfxPojvyvU5gE4PuZG
qpDcK33HBhDoiTMjPCG8k5KoYmB80JHwr7h/e0xAN8cEFc1lpRCeoAmI322DV77sKRjkAMbe2C0G
ydOkt0XUdzrHpOtLUvJ7ly1nkdIDgXVhttNuY9JX0+wiiOIfYd6HBhO8z6gAl6gQER3f2te1oG5e
fmgenWtVaezRWRQI8hbmsI+CofOPImZldggejGTQ6nzX7FcosZ4V1sZnL2WHtRJNXB2fzJ3CF+1Z
h2s/eYtZFUBKqQbT4fA1wOYmCP1tLx2W0kuxfDduIEV8vrDOTffbZw7FEYlkhLDadgS/5f5tUb03
cYp9I5DzByrrjZsOiGjuLPhjHl+bddC+Y0NHqU/PKidct+R6c46+gpqxUaBmlqxlzUxnaUAAjFJY
RIAL3czoHYASsEhl5CaS1IP3R+ctpI5UNWd++8TItl7dqfBK7q2Shhzvpi4bPAkl8KyP06Qw32f3
Othk30sqO4HEC5iVblTud+/NE8jdTsb5TuDUV0ZHvWVBa00ZdMo1XwyQahJx5vU7tIG3jH01AksT
U5kD5d21zY5uVqtVsHySMzjqmJ9jnh96vzvSCFLPweOmy9m7P5zxVrarfDlgGwNTMCqE0z9qc65E
AYDYokjUhCuCPBeySfa3RBZyqCkAZRkn0OIIQjGBGsAdGCBVbdUkcLzMqcSfrG5G5mvYkenjxRel
OOnJynxWmDzReiLvztAgpxSNnOKjCCDX2GBfWrIXSAs7xURWmmvYc15XwaHYgVkB0uGTLCKoFHeO
ZOfIENZJCX5WHFzZ7a/bLhW0sB/y4EsuSZGL0sqFjhqXyXMwNrjCvr+FeiNxLCQosQhVUNm0kiVE
Aywwweef25fZjr16gKL4+9L/S9PgKkXjqvQSz6YLDLRIzx2cRWDfZEaGQFYLqSlD/HBg5FMA7fQy
f4UsSuAyxVd6I2IwgH7qrVE+DoU/7uaipTQ+fHkbGsty2jaCWU0meaXz7spuCYPwJI+tMhb6jE2S
JZvN6UYFY6d7G/unlXha6nQQiCawDa1eIzQksIyypV1jtjFnMA7tBt9yl+r1VI0yOpZM66vv/WnN
72yeY6UjxDhCiosvPMytBAgDcwpN7yihCHmo7zhjSlramMgKSFLT9oRUws1a69d7mq2+nW5jFWXH
KzyjhHoV9wmGM9nsUitfu6fiIufKGMg/0vuBReZFmc6Hhsa5TJn4IFsEF59XYTrD0lEMotKD/iTl
ME3dpFy6GTk/zWgluFzX/NW48OlU5KsiscGhfs80jUNcIBgdzSygZQqljkVBqJc7I8cUatwYC29k
18Dz85NwtH4+vSm+0j/k8DuYRoaYIaJdC0S95WvjTcp5A/Pwmq9G8/Lk6/mwjgeVc7TtR4iVjYSn
qrvUzyzTWByrj1Rlgy/X1fH6ZiM1eq8AEB1iuq+yvuNjpMVnm4RBWUtlg3IeSeBcEb/dXXK5udvI
jEXe3gWw/xO7JypSgJrblEa78JUig4FYFRhbaiUbxsWRyPc0QvjJgW/rd7R2e079SjtscAZ+pQFO
WGcrpW2hRXNmslpw1CyNLkw9A7OwzarvbzDq+6VATIMlPWLXL0Zo+ISFYTLaZnZUPXrXo3tAP6+D
nECg+bmptbInQELd+6+F88M/Jm1rBVgGC55C1cJwzKClEcQ1lKSXg0dQGOK+2z+Jr+3wYMIsFziE
UvFWYdmlBeiyKaCdREjZ/uYbn0ABI50YFPsd0LizuNyzFsJQhQSTESGJGGNS+b4qB/SV9CEhafJe
jLF3ur+Wf9iPKpPdea8f5WSCdiUTpJHwUAA0/wovhf/EQFuQjv++imf2D8ouKR3AvBw6l8QZKrva
rm3L8SenM3c/17L+753hNAjsPW93/O2SP8qKW9fS4qY1Hxxh8wbvAeWS/eUrEYuCagy9lNHr/JIQ
02ii3pqFMCENNDFkgOCV1d/47AQ02C9GxgiROhDOV+QNz0TDKKKqRO/H5dX98SuGcPQ1hWTJTHIO
0IBH24yhwpMuAFUyJusbHojXt8Yq2fnNEs6/LmGmsvIzev7X5h8YYRQ/ryQ9r8NUb8OIMCDtD6Hf
JPn2aVxQMwdqYaKf+zGPjpalIQMOV1X/Z8RwTAl6b9fsn4yHn38aUChwoJYtCRyQPQ2YY2/+Xpre
BKgqWJnmqqD+0ZoNZnsoQa7UKStHkkrpriTE74vIA8TlhrrmQKAKM/DZYKTkn3cqRSHoixYCAXXQ
7XxzNWBJYjsGKWE3noddwjP0GyQZQZhvbAHloJZkifPunuMyySEcDJ1ErB4JJJIhzQd05fh76Q1I
Nc4yivhLuIj5W2q9SYC2NF2HkRVuehkFGyLbQhu00EAfZKtYUxtwHJ9kaKEZTBNlTlRGRLp9WSNL
ozR10RdTMqosj5SPGU53v3wEISUp9UgZE9LkjOoI5cuE9nxKUcZxo1IW8zRm9FsFW5oroTMtnTRV
UGlvWaHppPKDb2EQUKjBg7lVbUxigTdLJ28A6JwYXtA/CW/MSO5vJUtI7QeNVwnW3Kiw5aoqZUbi
I9lhi30ia6T5LL57Fgb/mxYB+B5584WZaQYrJybNo7LbWEhliQ2XjZIYfQSoRUaQiCvg8OfrYF3H
mX/F9bKOQpyqJUoHXvO7yAFdiahojfcq1EbFpyVsfnF3rKV0DBht8FxMmFvK94j1rclEp8bOANxY
N7xhxMvVR6gaMQ76bSPsLRNXz0WbkbSOAfD47EGIo6HFJbXO5erydhj1DQiD9ovWgiKqJ5D6q3Mg
pSDL6ae7HUyVIZwHmSbtCFm/mikISEE0P/bRBI8V9iH26hp4mUbUsh2QMX6PDycp8ptDnXsOx6k3
fz9O/62fr/g5zNJOkV9RRqhyPC/DWQw5kGSZMXUNYo2Xa6Zz8SknITjsunT0Zd9omh8Hlx+/MwsR
xHXFVJznRXw6dsdgwJjB37uu1ktDXOLYENlOizyGU+cxTFyeav8EOV1DsCpaajpHN5QMNAYEO5on
XXgDsqcKYvoQZopqYx7mHGP9NeV9EUjAy9dXhtmJ2UmrSwRWZiWAfPQa5kEZug7Iw4Z1GxxCir3B
BfR6RRXVIYuDmHbMsfaHjcjYDecToIJLzwGA6QxfWcbRuHmMsXQiWR2v3cqbSBAs2mfh+pbopf+6
1ArZYx8I4BAKnvnqg/QSNkhPYxT7JYCOcrE+MRCdGPD6ncnESSF4G/tj1vp6lQlT2pzg6YUWisRX
HMT07Ihw0eRKb9Ywytc2ngsAKyD7xldmJvpZNQpHcUiboe8nxOgeJbN/iz9GzjcbDhyurvjhFXHR
UdmE2p01um7wtE+Fv558f3UX+evKe24KII6b2YwAToIRvcgqiYTzNSyCd41uysJuuf4DdNw0R4le
LRiJRxr20jc2/72bGGulqA5Oxna6FdU7Iwq4sQI4meG/RxlcmhvkHM4sRzFjhN58xY22pqm9TOxn
IQmMNNX9QcFsSuks6W56n7yCGaGMd72De1pgvtUbvjOMgNC6QD7jnt3vCAotHd4SksNZGSZ9t26T
G0ajA3GQ1IxYdNSyH5upYjJM/CbcHGjK3nUQesRVBlHruDtAwuob7pDy8GN937LpqIk72CVax3Pa
FmivgOzy7r53zsnIIjM4PB4hhBU6Xz7KBsksR6CwSKXhSh9ZZ++gvQArJZFORPUCrJKnn9nlG7hS
mX9E/qbxrxu2wfzzAMarzODk2Sz+dIKV4M3OK0s9PQM34jQxAFxffeVXr47CYJzGtMFNSqhY2vMc
o/Q2xYNmzMI52s/WYlnLQjePf4MFQ+dzWyWcKWUIhp0w92MCAqJaSYFVQ5+VdG/weQf2+5NoSb2n
8p4kZ8X61h3UeOv99nQxcml6rkm9UFlsfCnAtioSZ+b2dxXKbdda34pSXEaQz/j5QJ6MZiIYslMv
ipITyP5ku1Wm9FnpHifIeVbGtR1Ae8njsnBb+ou5Lt0JNXhTCyjkqHsPJdZRB7VEDXVIW0C0g1xq
GVk7eUlMHPOQTCV+93mqPrJo+/EcFMHCbOKD+pKzdFxKHM44YI728R2kzMASxt/WgL74hEXAvjL5
7k5zNFW63yil0zmvi4w/4Sx897Ins94dkxFibrsaRhnQeC75cfMHpMAPLyPSQZ8tRLRpYQwBl8TE
eNmPN/liYMwmo0L0XoYlbMhcazK+QKPKSNOOKUACQYTc1e7BWcpa7I75s4M/12OcnkCIuE2rENPK
CaOR4YCHjOhdJXaCmS5AccetWrNXFemOCHKRjPNbg69PcdftMvlO2oQvQ2vFIgav7k7VwPcQx3aJ
h0sJ7OSYyITW2MPo4GV+P3FKBLDpN1FSNI/lmn58PVQuXtwCpVN8YlDIVFIG9oHiUjsP/0YDYYev
kBtOlhzEVhpgoo+veKT5uCffdtRtI8jDg89W28UQKgnhM8qHQv8or/o5R8vMhlib5AJChE9Ixowv
C2LZR8iA5marrCkryB6mDwu7uFujywbHz8iyFlF8wRVwjTSQHGg2KGucuIt1lXsxJ445dh4BieIl
7p5vlEV8sZt2U16jGv8XlIV3tla7t8dw760h56ZnStMELRuztwiSrEUk/uVPYu2LC+S5uGaqjh/Y
AwpWoIwZs8ww5QKDEV4cl5C0boyoT9xU7g0xSZvZzlf4XTWlNw09aj8uBaG4ooeItmIJLuR6qzVj
bOwCl94RlvK3mCPpDJrIBNRt3R02KQSjPXdzlnTzcc2o6Vy32qsgKHOd+3/+7A9t0FuPdnHztkAj
DnLcir/T8xszyH+JkEXKj3VhDmLRPgJ6Q+nKjqF6k362qniB6fF3ATvfRKowdz2uSq5EvLkCPsaJ
qa+hTqCb0BU1J4ZZKU1/Ca/ptLArfVNYcNL/97ZvZDjWhKh3as01VSZESPASBmRnP8anTJSM1bhy
ro+hTm3TjzVfcbhH4Mz0NMsrLtQIgyJZAvkQHSdeUpjriMbNFNBPUpwbH9p6P6OoDNQI6HET4ep8
r2g7hkwpFlsp1e12TvU5Q1EKozsIgeJACStgggcUfrJttJ8/57f0zNG4bbEOLxj+MeFGJcVNcXRr
gvw2NqhWd6qzyaNO/aVd+m3kHlOBDwAIySOwDIr/KpkzWCoIXQxmzYouIElTDnYteYg5HajeUFYL
pHFEwtVCq7xyZFFD9PAN3uXBxCHI44W8mvYLGGAbigkDlXxm7o0boCOyh6L1fC0Ge3UOYC2FfpCN
0xmglcXVEitQm4Xe7swdJ1Ys8VknN1o1E6Op8cPnuUcaCeJAsMPrnL8isV2GaRRi8L5vBgFdPFLd
i1h4BfSj+tEkGcRhdgAi458CQr6mZzGuFI25gTNjtOUnpK1aIMWEgXsc9OPat7h3TuaN1/rFkhT9
GrGVUkY0z8NmVMcU8qB+CYZBL8gUj9hdH/6dwv+8F7NFzGht/xDwXD32YtmIkE0A9DLKDx6Eu7gO
YQFKuqkinyf8dAM9/ZWTstKkolsx+oWcUiaVtvoJ3xZHky9YnvgmNSfkgqT8ap5nOLgVkYiTKSnX
oTEd0SYTQwd8EArrhqK150Ky0iJ7wUwGItOp7t82OfiWoda6n7T5QczpTQ0enRq+k2U7pN4ANd6S
W6v2SYWlZo/Nuo7MvesNl8TFfRULmEV6/9385ELOYRvtcDDfhHf7NvKcHPWeFswxZYpFWlk4RCRD
NajXcZLXBWfuLLr/MDF9p37R8rVd1U//nNooJRtPd5l1/P0hp6enq3ap4WMlr2CZSmO7y4UW7+hM
ii5yzzKS/SCbu+jpNOWWVIo5jwcb5rpfTZkB1rsbslMgAhx2cs9LCswYiuPC04JArkOQDM4r9kea
WJl9vmTHIbJRH673SzDFQN/7uoFeaedmrSkPBPc9bjQrOoW7AiFGbKTdQeX4mpMi+B9bpwUkk3KQ
pYhjU4asMq4WBU6Ip3g+xNskTe2oexVHsxirHsg1IrfxfruGiy+jmbF7ZhMIFhdqeAuFc29YseXJ
IYK/WnafizHqhXlA2H89KPGGhw9Xqp4ejDa/vwGZUnDagH28+j6jABhGcLVG6RJeeFXjsDMdZ3UE
vVl3wV7jXZMwTVNv03BsJKAMs91v/A5sgO82sTktWwFN5VVlwSubN2h5b3pA923Md/TBUZ+4hyZ+
bmPi/LQiTF6Vt9pry7ov8j8is7SFcRO+jW9Xbg0l16OgK5srRZiII0byGKe59B1/xriJ47k0VilH
e5gq9YNjiRSqnAkeKSJ4U582owx0p4jsB5DKuqYByxGSMr1YQyTRD3cO2w85TPLFume+m15k5YET
ytAfvuxJa8ybqxEI/w4OAFRFTe6ToA+LqSQaGjLWp7+8yOOgFvpQyH5PCN2mZ0liYHatSkYVc3vf
SkxUIaRbSUYNKeeHRxuj1lG59kyyd6LX2U1FNqiLlcC1Y+yeiYYPln07mts0Aea7AinFe+8f0iS4
MsmDnp76I1QTj4DCY9/ndhaVZS0xEyk9e0s7V3n0q5hYAMaiLJmStwqMX89amSNSR+OxLcpmYHXS
mAAGA2rX6S1cQ6qT/Q/YGJ7ns7SSyiwDZcEEaFOwLsjYzH8g4R5eo4zRJnRx4mK7YLYuyzhkSUDa
Jj5//N+Nt4Guq4XfE55bhgiqoGK+4M3LgpJK274cGIfObv2jDSse/GOkxm1V4iXvCq6jRwBXvFl2
7fSDQoc/ZjHGzfQu39X6Q9rpE8SHNjb950l508qnz7/3s3pZ1fFuBmFzI/bNkR8gFKu6A82rTUHa
ybDQpgueqdBTvXJ88cWdsPfn6iPgaIGU9VAFLlEuj0s9Vs7fAa8OXM6a7yEoWQ5i/WZq9v5Gvbgm
grGfSV+Xs8hgouJYypoCwdZtIufxrQuQdwxxobGQnZoE7dFfCc+dywju5kNuLuXqkRe6f5pB1WYw
UTG0fGci/60Blkolx1TI9WWugkeFGwWGvmU6DZrJkwWDgYhoEcQepu9EEmIyIq8Zr78ARNWBtabz
if6VjvpbI0my1dfBHMHUqs4PSstfGY4F59U5HvHc6WXs7MFukoaHI96loH3YXthkG7vineGmXxxz
kuaO8qY/5oy7PyEjLHBfuneadEW2wqeo/FOac36kCPL3b9LwGrFyrikse9T8tgyW/fSNwZOtc23R
nju5UUzfRQR7GUyGugPJDSJPWSDJNlWKmDYaVSkx9rNJ5rMZZZEDeJyLowU+d4OvKzJ7n2quL/ec
LzPDD9X46MW5AdoThCxJY6qvuyh9UbL/c/+0Hc+5jOieN89TIIxnujSUSn8P21dcPMZCt4tdfQZC
LmEyOS+EHq5w6O//SNTO7m1dlU+pptvFDFlPTlVz+Fn8IvpAL7Q7AoZUeC5HQQF1WkG+MrbWqLOw
N8YA0zzt+lF+JG9P/Zq+mfQttqlDQFgjX+gqPZsMRIzo2y/SoBTKB0xdT0fGXHZLjIzh0pXCDwFk
CahRtpXedy40uaMQIy7uRqyRlvvMKVoMkc6EOy7OEDMxMWh51TxSqvS7467lrYj2Qj1sZAdKCBDS
p0YOj5RxCoEiN3PRdVx0aS8Ha1TXbUVHonlsGArPli5TD9QSmsvp+mTFTval4laUqaYBGOan3sDn
Lor3nd+DNcUMJKEa7qxMFIf6VBWXfA3ZAxHL73SEil40I3z3utzoo91Vo0sKsLxeXOtzQaqhXGIZ
eAxnskaVnnu+oppStmZMOg2cso57q+dp7q7U3hbKu9+Fkei4umNlPlCTC0aRjHZc8YtlJnveZgNB
UgT0IUSuprme/ElC2DbaTLam5DhS8VKaSZRqL+0uM+gnhsYLCUQozmznhldmU6e3S2eGGU1KqdiO
g+FCCXKo+D8jSF+FMHrFJppGdFRS+pOh0uZe/uUg7Vlq79BdW9m3Q5p0nG+MfATEvE4q5kBdty2i
uVpYbi+wIPOxpT8BFte7xbXfOpJX4dEoSm5XqWWWWmhf3xwmtSJsL/kwix14iRfjKpL/QscHbCFJ
QNJOMJfBVJO5Z3av2fJpbpGKZk7xr/w0FBJ4H8pwVJvEEKfoy6vPYZ7wGDa58/3O9HneqAqydj5b
2lqBY7758gGnfaaPF5eL4uLeZ2kK14BvWPbu4ZMLvd9cdhR9A4piBYr7ZLR8NHbFs8WIiNVpy8fw
6wTfyiN8OW29yKSY7gz4ERWBYjLgiy77c3hUbg71G0hbfGkbGBRi7MuVB+QWV/ZlXYvF8D/ApU1R
vNuc+XWIFcznOyZ0AwiXxtGYbgtc9wGANak04zjgMlTiRoJYhd33KvsY7SNT2MpggdfnnMYQY5fj
r5tORhDlibKJXCcaZsjc22GDw9Oq+5kMD+zQzeSGEc7wEvA9ii9m4bLDY1EHMWJI/6t/x2U9Glxj
FD3JO58vfFNquFhtqGFfwpcGSWBHW1rjkdmyfvwmYiohb/tDZNWntXIuYfzSrjO5mMlW3gpNLpee
HGhWFHWrO/YWWCF3Ut9J1N3/eWKvEj1KBHeAig8DzfI7mPzNG5POUrVYedC4pMVkUrklZVWuMgys
d+2Fp+A47Prp6RULqpI/Sm46fUrDT/rRr4SmScuwYX5XLoVPvmIsjExo2ttYEpsEvb+mVgABeSkk
EIUE7p/PBLuDwcK/2uyzwuysShAm3mqx4+IBhFbcBqkrTbU0un5S0V4MEYEfnyYjko2tQKuf4kjM
KdWd66KSf9OhdCrsz3dIiippAt9qD7udEWIPJrjWmKbnPs2xtBKfo3pxGBq+z/dhYYVgwfMieiZm
drO0rh90l2CfDacQw12+6wNSc5ZT67EIxcAVFPGmHRjcsXF++1w1EyHf6q7mjfmMh33ceE6GtS0r
fsh9Vz1iWmjDZ+MsIHBxRkmRrkPvoSWE3iQhXy5apMJSbXjTXMRH1kwQf3tCCaHBfq5cbPEp0Vaq
xPHuab2nCs9ilCXPwheCXI8RYY4EEzKkQoX1rN0BFrs1NkmOvVJfMeMgg/iHDTIOBeHit1rTe6Yn
Qc7bVtqf/Bhma27yIljNNlJVt3XSLIRcVzEwtHnL+Ws3Fl8qWwxWtEtqeJ4gHhuNBhNlAProLEEU
g9fhCoBlPtgAS9Du+XtLoVsQulDXW5NhZgmCOYjYW2GJXqd5Y0A15cSqteuybankoR3d0JNCsmE0
LO9lSsLYo0wESp/LkXux8RdeKEWpjekXjmmG61T1evZ/xFbRw3LLl6qchr/YmI4C/Rv8EQt9wISn
rXyI4qKBLdFF12r/9s1sQq7wS0Ip+lONMXkTPsTyjQsrY5+PeQ7+9A3rxwKdpFB2zmQ+skbxApAc
f+OyTAFHpM58/RG93JzUlMNnRL4YR4Xd4G0aA953yf/49TYoCUYxveI8l0BkXkDAdynIuNdxs9Mp
HgVdbtdoGWIeTSL8yNmSynKhbt1D+7Eg6F2m12P9ZVCFOSAd08adqM75RjuBzGYuIKeP5XHKM8hv
sFsLROOZ2DaUNhPJaflMlpRuA2vkleG7YROuzxuef6niBWcf23wrlSFp6FJ+nXM8ZsfKAv2kmgXZ
lYoh69DGaeOk1p1ymuGiQGz5XS7UXzDoHQrQg4rr4eTVhvfbR336FEMqrpptczdEVJzpqJUoqdDV
EWF5TlJX0TEyIPmIS1SPc0wAmiw3VleBMymUWQtzwSdoJcwtCbA8n6Lbl4+sABtLUCB46jTfYK6i
3y3ejZxHPTaakSzc9QTGUt8YQ1Ao5ztjDTFAc3RaLWonkiEux4M5WO/PrdFSfh+InaUwEiq0Ttoo
tC3rZQUenXlugcqBGu/YktIpvc1QUSvAYl2X2smOPbzYgiXDWMCzMcDIJyGsLmSpVcQ1ma79LPVd
wjVR4V552fihGeViO1ZOgEirA6eUHRO0Md+ab2eiG0b3Sb3EE25QYSsvE668ZR2EXJitF1xOzfyY
Xz169ldD9pUvwftnQNlyoS7jHlHcDVAlJC7sYd9HkojOHzSSJxvWqD9IJsGm18bsMR5BgfoOXm8a
3on3XFvuBl2lmeKYVXzb5OGwWr96G1Vp554jOlVAf+zExyDMzzv/8MSWYk/bqcI1gg/X10o0FWEr
AYnSvqKnYXhoEOY2SntBbPfB1Jmhi/0b+J9VQExZTUmlt+RjJHVkMbDEHjIpjndqV9qXLu+C9jq+
c0kNcabY8O32cvNiZFwkRxyRneZo43zpMAyy8ulxTfxNw2Qiuhy3tHhj5vnpsOc4FSJfp9gfszUS
J4zMxT4WYXoBnHdzO8yrUbj/OKb9VZfTmzicXH4u/wdukT+7Pvcp4KIAmIJkA+3plysCUgkVu0wB
GDOYyQwCKj9VYXV8wEkTHocAZPk++RVmdAQRvLh0Fa6T1IMKGBSpVNj+He0ZZS7Zcfpe0bykp8Vm
OUMsCk58t+ygTS/pJt7CmTFAjo555NesgOZt6FXgMwp6zwAgNjt+pmDatX4ChIzntCEoKSMbklc+
0M0MQTiqk6krQwENKCs/LFDtaOzFZMABneEWrwW/o9OIhsrcJyLARU4swv013PrvG9gJXj9OkmPb
wm1JPDhH06WLHdK2Timu/8GUpJ/SyiMdotZlf0bQdCIlWkgmaSVD7ukZQ07n0kSaMIlbcIkCc3sx
d9NInjVl/q+vTT92eeCbZMxO8FzDUJZSK2liCajVWLiZyeJn+nxoVJZsmTLchoqMc4UPwBoTBElf
NdDYw613FhPtmg4ssOuaHF0Pbz9kWyZNuL3paClDtGIQLlGnqyZKKpmWdMYH0QXKCQWbfh/J/2tw
0mD9IXI3uZr6YIFds8uK59dph1jAj5RSrTiTWlEm8Rt/q4Ymt4URSXCvhp8IjGfFYgy7Vr2Jgg2p
MzIqmXzVWdVhtneEfz3QhK7It6C9K8Dr5G3SDYttytkonnrTls77ifY8Bolt4/YD3S0ENNf+/s6B
rXwIK9OLfHxv37IN3eLs6SotvOeQlvctMXYC7IkzIV0coRbiARM6KAZWlaJbgzWTtc0i0ioeNjIK
AaySENaMTL4GqE87wKVOvWO4v75g8HaVOFWWYTv+ZAHJ05mcUCRVz0bt7j0IQHJM8/qFc8nmd3+X
8Ra8OsDL8AYPHp/tCfZoRbUSHFmDESyHal5DpQu/CGEJwvKeqKxaFj26f2gaB5+Lre6EYB3mBxzg
buC4QVZEIcm/n0hfTjv9egYJkBD5n2Y/HtiAS52x+iXnRu0rGTsRfVkhEyN1GjvGnc84o/+/A4Em
OcMLHFyEKqMcU2ZkQR8Xbum0XQB9+k868cY71kJ1qYbfni0JeAiBzkkr/c/qFp4LhvMLvwmFoivA
PmMpYOLzvkaXgnDm2zBAOt6LV8xA4xaDCSPVYg29GSlAeCWtJQ8W9EnnEyMiwjE/gzXLqpwo+b1r
rP94DlQqHcHCjTYRFE7guUYOHBMJZ3z9xmRLOI48Az+rY8w7fp18bXY68KKQXFv0ZhbpP9G+74H5
nvILnRLHuOnDb9QanBD7X+pf8do9NjtjGzzTKKxVPXk/DAPW4q/gF14jH/a9QXeNbSfK9V8KY1u5
h479BLxC6F3ka1yNLiaW2roX/elgU/0omk7uaWU1U5cfoI8wfWLRUZOn03FtivBdk9Mm05m9WAPY
kkA1cMdUhquZn7x8bgh5gPaolMIrSRyIe5UmZ885u0q/GHpVUuNEi9X7sZ6egcsv6h+iZ9bTbisc
3yfDB8K3ud/7K2u0SfoJgEus+tnC2bG8bxiOSE5xpW3XnlCb69UIOa2zVEY2xBAKStoTMCZ98diR
WBfj4CL9CEWWUWXHU3Jcb5hrM+hoSJ/til+lM2fNNHEIjua0o/yvH4on9JaRPwchPO6mJYLyrVW5
MT6hFG/cG/pG+tRjbSdBa5KolqTv3Ijy+5gemCH4uYjDtbnBEvVkx++nPxI4Sue3RUR4jRPqBQQm
G47+2hoXYm3U+TV0X8mvsa+wT86eru+gSqaztpSUB729Wv2YCkBRVTwRxkRWLqTBBLrgcydSgvqS
AvdN+xjwCa6L9Yk5BXphaQmZfMbtzRe7x8fqEDALzYxQXom+fKJd9eO9BUpMZtt4tJF7U75hiRlO
MoUhpE34muJ2JzPuoksCM1b07BEoAnSZwLm1h3Jx5QphmEEilsUEzvX7/mlppRbOPVZXOzkSjZ0j
gJjkRV+ZiiUfSzie8AHpwxklYKp8Vk5lPtizDdCMtNhFOEUeYpY/pL6rm+C6cVhtmTM1tCIIQ556
RX28QSvvb0xvCw/OBEg8L9BCNd7JSooxT94Ib/VPlt1QPm6EV4QOLuzeJ58Kna4kCanRA5xVky3F
A7uW6NAXlr6hT+HMNL8gdEcDqQvOmNHWLil5yL3dkb9Fx26SGSKae4Jp6oYcjEraA416XNBXvIUV
rPB5LZkjLLO9xZxrlD6LdoU/EC3295vyWpMyUm3m0E/Dd4k+DETnncmgfDG6DtNNHqUSTxOWT6IJ
fyu3EOr0r0m/c+O4XjPf4A48K3PNUKlo3XQ8eDhCtKklOwmiwgQKSLZdtBVeoM6GoeWPli05XNv6
lB8HQI+FYO8yywwgOrx7w3arIFnq/7HbSbUkFciPCWGJmWG2VnumLiIaTlpFW7j8FSua+CBgJl1G
kDNSPMVvfMQLQ7yMTLIrRvXuSm+j1C4wCTJRvKsh2vQeD1aNQwLfsso4mX7kyOIqxWW/sxapof9W
J1zXxEHINcJJmhG2d0LfmnPMzDWdOFbfB+PW+m/8iZHTrgdq+SNtQhK8hNPVFfk/ETkSQrjrcozH
0TjrQ/sUMSbiWwYz3v5mQjMYO68PHHtk0iEBtcFvxgozvoeaXElYsla12IEOtle32tknSjfXbzpw
ARIxK37taZPnrLvK5xZGUu8r0LPRjGZ4jth0p8zcaliK5C+fD/RjGqFJjqP2w0CJu5Qvlage6mRC
tuTT/Re7CBWD0+wJS482WRiMQS2EbdbZt68QVsuXeLImLuS03alfE/X5BdBJ/19WFJg58DQluxIB
qQfm++CQpF/RPfwYY5oICvbp2tZz4GgR4lJOOMW80viqJXlCXaL4hKSVUhASEEiwVH1o0E7zoIxg
ErkCEqmw9jjJLav+qhi3eJgOHE2EN9HfV0iEOuHmu6rcbo3iZXpvIf0cs6B75EuIsDUqrfilwiUL
7jR8+sgvuxJfO3+oJxnZ55e5/2T6Jh7wYBy2LhXwVmmsSxVAy4OtRx5vfcypEs0XKRP7lIObShjh
emlaj54eJ/Hz5zi+3V6+NtdIOTmfRIf6lgZhnUWeGqbpE0RZaFjo9bFI6pPvrrFctqCs9bKIHuES
yFvjGhbjpMmD5o8RXN/jiX3vm4TQzwIkI+pQauj/TyddLcTB1mA3tuvaom+Glavn+UFIIsbY8/Wk
FuzcTyx0e9zMrxk6eiqRWUKqTYZtcuINZkqTikLdCFoZ/CYJJmhLOsMTfo1IaPMtFZNWj3w5KXIc
LFFtosoJ9WhNfeJ23Iueh2/Q59Iy6xEOlXOYoK4NTDGQrOBn+d3+19rkMi10WLr+NIS+92P2cjDm
0YGfhN+RdQffmChKFEqzFLQuNy6FWQZWQv4M0qABdlrer34iN8JfdMhFiXKa7VowCq8Aph4ARSub
nbEu45V6qV2S6qZLhcz9766UXbEUPLbw2trn1cvCxegpO/v0/L6BUrgP+uVBCHlMjJs3X1aEcIcu
oOBlGIfBkUsLqnIO9nZiFIESYK1WgtcKqKIJPUDgNy9B7Lm/N9FHU2PjKIGhaQbNvTfE0X889jfw
fehf6tWo5zA84VxUELBMgXVcymGBS5NgDRbxCj/6nAQJ9s+Nxd3NI0Vndkf9Y2E9v689C6sbSPc5
k//cMSR4ruEAlW9RaU9q9oRE/bKH8WsaUrQdbcGeHLxJFJnUCAgucSK1r6KaHjasL5xcd9unX1Ma
3d2/txrnqPxtBccS6oWL9lrYjsSL//D2zMlcYkoIRp8DHuFQ+xySQkpo/is5h87JcOzoVsz0gk9J
PJFYqkdMwVqHZBwQJ02CHJ5wxQ3i+9b7T7549T2ln35FhXF5/xXeXct1RCDVU01XaXpPKq2CKcaJ
jYNKTP03yPCTRFNiFdotNhGtl2+S983IH28Y0LaQFy33Edb5zZQlCrGEVIuMFCWvR/SaILbg2yIE
oHa544EmiRZYABuAiWqW/RnmApUT+ZPv6R2eA0WEM7SISHZyToN+On1EQsukb5GOaelAG10ZKRCi
+TOs2D6cKvhuO9z3rYxlMwMS/6FdFoybtxARyffpnjB0/fadB/7qGZpQrhWMHOq9XwB0coWGQQJQ
OWVXjlLf4BEgCou/cle3+Ffovj4p7YYCXECfIck0kE7gPKRV+qDkpqJGW6Eir+lfkLwofvTg2+vZ
YjuyrCyEJdx+dhRpFpsMR4hC9Hjapv9hxcodCrdhtevkUcQTVitatB5QKJCjLUBLf6RlOtjrpqEN
M1dl8+b8X4zm52l0z43mbMb2R49FH3U/42X2AR/+hJkk43tSG2vXESFY6CIaQNl5RMYG5VajjxTw
217fjLcQHsc0fnhppkUoecD2okg8/vQ4sJE7vauZefzBPExrppj9DOsEAOED7cJgXU/kSxSX+wqp
ofPXc8IeQmIY9s1gOh5NEiCcj6nGApU0Egsx/dOJCksvzY+qHVV0Ydy35lIl5QWBaUqDQPtI3dkD
hyA2+1ZG3DcZomz8Z14rXaMOeAAoshoX62r3WSPPBWdcBU0HEOzbzuFJ1R0CgDXD2i1Llk4yUiYo
ZJNFHmrlMh6IMuJkxP1x77CW6IBtyNqS7PXnOZx+CA+h2kXvC2Uxs70xwPgIjEBV2HYS0RQpqI/i
nPnfM5lUmQAGWZKt+35/JdVYP7IqPGCFdjFikiFjINMqK84IUNYHLB/BpeLOyEtyIT/RId+UCYYb
noe10QgSUGdVuNzc7KyDg3MmuG5/UNOA52XoObUSpi1ISvnWKxg5IoNYGCaDtfnMkby2q9fPBXoa
vQQ0lsBiAUuqL6GpVRfXsCWGzFtQUrqv7H/3Dn+RiwttuyK7k35sLzLv1FHMzStacM0vgMSXDQPq
Ptl+eLDcx1/hE1x2l/4YAKUJpxFQNCPBF1PVEElamWUa6lphms6KDQxhsWzdy01ecdqt5QsD+v7q
wVij61Sqrnf4v5GGWoZUZMxTWrw1PO3pdQpXZHRqtHgYsMJsPzR5iufbBVdXLxei20gvemh3yPb/
+RfdKRfMNToXHdhwqL5G9wKg9oMoj3jOh6r2fTURxqJEIcA7UVCFjwA8zsPMf7+5xuEKr3CN/58e
taTa2lDfKvo9JB1Slqv8l4/tFmutRu1997JdlHGTBGqLv6gwur8DQ429QmwAaRTZKN4ldvGePLnL
Qmha9xIcy3nSlFJXNBvCKphs35gwmudIq7eBlH8vwJ6ugPrWOKSdBJOClJLotkAOH9b6DvBJyEp9
ooR/0hhJViWrF9953ueE6SPlLjrcHrj5z/IAVCVyok729Twvh5NU/pUC2uM7uaScgRRZ3UIpj7lx
b3zIfiqrutGoAhJAT+hKb5deCkaBJqTkyGrkwJApiMcC4R66KFVGzmQ5/7DnCjL8YT/57o4+tK7+
708DOIEGPi8x1KGWCv5b/rCVbXakFTZ3bSwjFDxl89SOnAGgrqpG/I7pFDmXa0IJgeRjzGcfLh9T
jDY9053A6MtWLq/QaBvpgovavkCjSzlucwf++ePcpYFABZnOSd2aFnxFGR5fYXXwsmZQzgd09Mkd
uGwdIo7FdaL/ifmBnJWDyNTB/wykxBnHX5f3KBChrjSnpoNhrXNwlf9tSU8Uwsa65MaF1cvvlYqC
2CFl6iU408+BjNuzR+zp5uFRR7cc6EgYdqEORTyzJnDzEBUU6qUmogcNgG69KroRqMVsAUY1BBVv
AmxC10utRb/60R312HrotOOcAaWwQvaEhsz5uTLD0tF9eElUSx3uVXz65rxHTrCEOfPcG9S5FIxH
rA0AlRIq5YLHPvDSe9zLNU51R/7h4fp+XLecuoyYciYqA5C7n2hbE6T6M5ml2Uq4hCQ0vaBo2ZwY
M77CDjUkFuA3RvN/zxhq12ay/P+KE0xbh1YYVffifk9nEyaay2srVmdI4SKJmV0BCM8XO5JrE2qU
3BT/VyGnYhNcMxMwIccUZnBAaZhftd7rB3MpGzjBGl2yiHD7eAUHUR4oSRCrZfjD6kpV+LdlxA8z
US20jWj+R1487ZQU/++edi57OcxYC2oNt5EsX9F4PSCxH4REdFp5QsUVL17ovJ/1vmsIbMNdM2RL
k2Cu+1fPCPcF/eC0gT0fXjSmLkHAWIwQ+HthF0z4Pyp8+vtrgeU6yYdiI7j6oyu/AIYsTtm3X+Ms
sZUTIftpLqOgMSDfEXIMcLaIBwauHpPmbQYa5iSO4ULs4vY9JKxxrzxCNLSxPX07rdXUAy5aya3t
mH0K58cLk2AyrcCVhfkURkYAqTmkBT2hCV0kZ/QkF77DiSPgOzVwjdVqgkxOaGGqB04U5BDhZZaD
sJ7Id6ZEHCNH8cGztJH0zTQYGJ5obaXQk+ytG8JMv6hvkTgYrG9ZWBBYvka1kK8gY8kVoG7IjzqM
S2pnnjNOnpOJ6HUDneuSqY6lBHovQIP1Ik5FSUOFikdX97eLuJDwJDFWjwRNuQZrSUI6jXanHfIt
ndeoYrvkifwi9MpCL3VSriZu7BUB125cPqrlgu2Y8/4n3V9sQ7puT4OLTOIqCRO/7FCWWRvatL7b
QiH7NGzeBo8lanBC826MA1rjR930+SYnwzkOQaiB7ouSsoZCOUT2ct4kkZNujGrFvEKCqGTcXt2v
pVrmafNDRfSEZI1IDqChg02/O2siglrPFItgHsgAkwbIC6PiU1n5kqyqGmXdy10qsYgcrFbgVlFE
J4lJzG5z8iiOS6/ylnJo3PCuPBDnpM73iJj1++hjwxKuKhPH33xbqCGV8QS8agQQZ03Oh3o7sosk
Qj/kYdmH5eqR2aDx9s+Ae0XKRsK64SwP6Yxhe6n+SdH3CqE2wnMRMWK/PAdGL3KeI44FkREHmaum
KVI5czTJIk3cPaTasUF1lYOWRpyC+iaHgWaQYZ5b7JHSCCfTGJ4R1oAqoGjqxM1mOEbFZjon3vQq
YeOM9iku7XwbAZwXtI3KNPKTmCaN5Reps6wz9nIob3zUg+13kosTubFJlvyzVK96Yhek0zKSAIJe
1zBnqQwXDt2IIpYiA+/RLl/xOA5MZQCRT8/bog8vrHvvaUJXtxc2vybJSoqvl00OFYHXhJk+L5QN
Snt+ncmRAfp7wOw82miQLaj2sb6NlYsyv7lpEBK8JOYMeAUjRluPX9KGwYQ2wJleqbZR+d8qykEf
ZlLk6os7iElu3w/adnd46Lh2Nl7jdQUbcr0ZyHexEsjN1yynN+AlrwHLdNABLYb1yrfx/NLe2zOq
A2RnVpJIMlmnxyOmWIa3Uu5BUWpE+rzgULi1U9MN00k5E6QZM8mQLK0XVG5g4QUc9sJQVVBkS/2c
kmmXGFpCRGrz3GOyrB913N/PFTdYnWnkJ04XhI1zRlkkByQurBH0cgztj7QOu+PmqJTwbsjkjlib
6jiGqmhTFhMkXiVQv74lypDwD5qqdgpFt0j1vyuiJY8Dcfk/UmZhH48SkhP11YGc4oPith1IX7JV
+DpoLY0MhKa/qNBTOjRLd4+f7ijVhw6tTrmd1thdtVXsIJKVvTlU6iugAJZXBbwWUtq7i6/EL6s6
Yxd63G5VU+RxMBCXFlfac2hLzVmv2r2xVVNzhJRhm4Kgkkq5BIdlr+lcH3PbmpLkjFjeOPLJDBRW
WW3078KvRBcV8E2J9+VZQUZ9MwlzKiTgQwD/HJarKLW4YSANA5wADvtNSMNCIejZ3PupLFp6NqhD
OmvHnjE2Lye0GaaEXF06J/rFrPo2S90GR3reG2QgYVmS2BLfXkbDqjKrs1vo0LCwroLaC70/Kkx9
6Y3KLpOCzA6x4oCPAaaOgBnnNHvrIKnptGr1lUwCVueMZqIKzzVgbA5bJ/3GlQQU3TM3F5K44zWJ
xk0KxCMcdFOPKnU+gXN5QkxUbP+UXU99es62Olci/BXipi+5HRE+hsEVkjzPqVpMDa/DbjWTE5CL
oR/u2K7ljAByeoA0p/M5O1HoWKeb0mkqljtZKoVpJZUWwY3r9C37amJia9lbG0BpvXbdGr4QXk0b
gYMWuoLHYl/mUzyUOH324hK2wowmAfLVyEdlACLuyDeMHI/Fuw+ou29x/r5zHD7YnAj4rL5LcKhA
rOEwZ+UYWLCy7s8604QKzpdEm3tbEn6u1Wp/Y+TcQs5hKf7JUuXfwP3nQEofuMYfMAvQekW0izMC
47ckGSN27KN8gQaaqUF4vVX/B9NkhEcRidQBgbNgYARo/rZGqumbU5cOVWjGCo0boxejsN3oVt0u
Q/N+C96V/U4/KWzqpeFOmurL0+ZXtEEa5KxVwY6Sb+122doht+xnpnwopgkspIPMUwjbGR3Y/G09
/NZekMNJLBxzzFgmKkPrbdV4MeFH4pddPQQKb+QPdOP+ullIamx5duNwMSROKP4mwIe0We9CE9/S
94ofVaNC38ipQxwqR++neHwGs1J7rFz+2d2QGuGsDLdYKL783AAXyJpYXmNi2EcK6N9I75w99Owv
bAgWeMl1gb1krpplpnakhjMMLl20gTI7ApZbhvJzYu3ep0vTi2lSR+Uh5lHANrgcgWOjgqnrXIRB
8tSvONws/RNwdbnSMNV+Ft5AgTR2dR/aIGnEam/C5SZ0ANo72OFk29TJYMQCExT8J3AyjFemkKLk
CnH7ysU2MudK03GceNA8hl0SOfEtYLshysfOtnpe579rRMMdwCiTELtW1qvtdMEWUt9k1o+Ci2rk
LHQhZJll4x5DDsA9DyvckKNlGMS4pSev6076apzIQm+i46xkXaQKbphYlT3+aKTcakcMMtC6yaL5
OZx6OgQDJUK0gt5WTSgzwcqaT7/rr4VFdu5cw+TV933fGvaOudWkKKWqyGR60hkmiAr3pB3UUy4m
10zeD/uX8DR9iv2n7qczX/N5sMc9aULlJT6hkmF80QrcubCclgftTNoE+VaTw32elRDmUh8uZRMH
EFlPMVkHX0MgsIwkbSIkZqT2sH74n1dssPcoA4mOs6Dwn12nxr8ZzHf5QXVajPkrXxU7pt+L1FbU
mEIz5NKW+HUCavHf2Tx5DPmAgW3C87UyULSKKeioT3wc9yy9og38RiT3vSbMxXAo9ZuhvJfq86Vn
+TD5gf5YdbWMDonYx77F6Eg/7iS5gVG+xXhHTc4z41mYxvZwQ5EWx5xNPBalSgP1NjXeJlZPFVCS
noX0L60xM5ZdF8JVarqvy99XxqfkiwcSSD4bCTSQPIf2Fp8H6m3keQIP3ldGJm4mPSClk4Iw0kE1
hsh18Zqhb8Dn+/7jKt4drxWyQaKLldML3aLT2BZ+WnRFVjnb+SXhQtSR0nJ+4wGvtb9FrYEilsEg
Xubb/Vr3WOAIhh3Qdq7lhBQdXDNSc14KIbMNXUfVAdip1drF330+RNhmCDqQS5dgonogmhqNIKJM
0+sjC0u9x8TtRG82dpF9oIkUbyiBPUDSbYy5rTCgXuBYrRJjhLaD9yLPtVFtA5umGMYx3B2WrR5j
nogXuN5doTsBU5VFTti0NO2mXQVSaltE3XtN1ANYV2YSnnv+MJdRZaiarbd0vTnr5Nxpt0qegzgv
+usDyrBgS/sfDMMkpfP7sk/N/Tw+RpiGbvvMdI4ZXNS39i5sX8ZS5DU87ifSqd0lriPeS0b9Etuo
x/fNr2x1P4mlWaUsEbOYHR9sMIQyn1ePkvrf+9JObWQyCDwerLIWHDwODjth2MZ4JVfvTpibV1as
oELT9k4+z8ojV9BRz/pyxAmrGsUyE0n8AuI5fsEtdwiIDq90qxma/UdUw9GkjusQ/mzq9U0Qp4/c
kNQB6J6u1hYgAOD4JP18XZ4I+kshWNGn3eVbSYCrp5pNwH6VYcsdfRuOzKAJDQR3B6KhONfkJDCk
UZ6g82Y8YCrmYmvyhDO4ng1+OLbh/T1+SIq+jRWYZEiuHpdiNM2Ml/g2G/EthD7TWKN1993iCR89
/SqwM75gNWsLZZSqGmNXU5e6a1fl2m9FlJgl4vhyr0SFzRGrTxgA1zVNMkorEaU0027gKQ6COg+Y
16foB0+AyKsYG6ZC8QfqS2+dbBX4ngccwZJDgiE6iextBiafYm4Yqq44AF/fi2vmkX2d3AI3/3qI
EOiSFPj13oM9cHaKHRav7QYa40VmyQ9EyIfsi+CfWDfE60xi6nuwzNKzHBygOE2eD8lMFyoqPLye
ijL6iqqpVOi/LgyLSjND7+dDeVoXWYvuBqPx74bIqOyDBZeLE0zW+L3Vg54BOFdwKygdGrQu/9X3
y9eZ4mRL+89L41Ii40WTRMzshfBl/HFkBQHkcswJxdqIRWETFzltIcZggnvaomc385LHh5sbfyAR
o1MLnFXVAfAFuyXNiSjooWARubMPfk5svPxCVp1jJLysmR4xcOv+mCuQh+GgOYV0FquWmzz1TUUA
LueNrOcvzLaGm7WkH8fPeNvJwYdLvPRhUli4i8TPGv14kBHuqRY9hFanSFtJEufhFgBy1nmfT+MR
a+rsfgAYnv/Hp173fGxoc0dvfq1FPYVKkoDOD8pnnLODtaap1wEETaVD13k82pWHVfNPllO+zX9J
314gM0sm7PQ+rcVtayKmuGa7NaLGx6fBRjca08jX+ZVkI6+aW56CEskusI84Jsi687JNmhTmOkhr
NQth8TlpzbGkCT8eIKThcE5Ra7H4QP0Xq+zm9OlgrJp3HfusUKx6LR0FgoyLYpPRf8Fu7JJAUlTW
+4KFTgpfe+C7op5cu40EnmCNhFwn6IX8JZuB7NnqcEFTU2h4bhnXzwGSW1vmGFlbVZo62U3xnUlP
0rAWokMPKkrF6AmBcIGDKgw49d40UFEUEs/6Yi7NwAorXI+xATK4nEv28TNiuEfJwpFMgjQqlTOx
Ut+noHdXCE+4veRI7Z2iK13IlZ0xEziVCLTp9JqOsct5Yj1arZfKQ/BCviaq2FHN3Cp8CrWzUS1u
J4aMUiZ9uk6IREcMldsK6tKSIA5fciXll0krrVXZQZr7an+6Uv+SMVa98jtKg7xcX0qAM27kcktx
Og7e+PuVtptQ3oMolT7Efd0UBbnEkWuDizpVYnCkZBXq9aIhwB3I4zQuo8I9Xf0cjncwkRtNiz2T
temg+FFZ2hpUVXu3tM1Sri+TuloOxqgN9HtT06lFvtsjMfOTPRalb1aW29ZSHtMkE1EjeqY/BIe0
z1hvFf9M0bMHTk+sI+Nkm7vKhw9nqEHEDNVmTbg8jtUnnTCFGSKWfpQyZx0JErjViisVMisBPmhA
lKtlFQXNJ+w7QvZGukqYrN1J8BSZqe9x9KO0mH+Teh+ozTOpTbdFpL9ExJGrQl93+DaEyPhgOqqB
Rjc76ZQJ8C68QAjXbx2heFl58bzk94FOl3pTAhmzvjXlDyyzgRY8SUM4ARDtw0ZAXN/kF44y0Z99
SGSo5bPCmD41/n4rjd5bLNLy88b5tkEXEwDET0mRJ0IoR3GqqHwvMMB2qqJeOyPSs1CVo1otEwrv
c2ZD8Q8KyGM2ISqaEQJS06jVWyOTHjNxGCuUdL52afmFiBjuRVfE9S0LQZuTHEshmnRMmzg3//iN
ty7txXQX/PDs1KkLrWJFmsxIOtilgIXJ9s7UcJ2z+HJJHg6Upvpgpg9527o1gOv/6UJ6hfe3rJCc
d0/fjTUeBlzU5x/uNKLc/DgXumQNMq6D9nqXTTpPlm49YQbZYrJTikpb4czHdFZ9S7MYg23l2XA5
FrpgM6ql2t9nwmQEbuh5se8FaYdpw5Hqw9wrZSfhj4rsy9Ajw7ezUAQLUFV3An7g1vop1eSD7RN+
kolurrwpZYWJV6ldQgGUny2NPdE06/GhyGUo/mLlgUwh6DBFm/FB0UGc3WpN97eVhTXxsmZ7Kw4p
JUl/X1zlg/u87zxAPOQyGFmdTtiu+88nggtC7iVMFl86jWys3TFM9n6aZhc1wrA0o6658KMAGEiO
ALQQsLs846toYqsQJAundLTrAxbcsjfI/FavsLCiOWwp38xkw452eCwDExIv4oNY3xnAhD5GoaFK
MZNtX8aHBoaDO/0/qyW/Y6rvg/59z1uZNIUYoMMwDV/k1Cby4noe1LBgnAbIYnYX0w4MBsou3TxG
9IBRjv1awYte37v9N8bxhLC3ZQGNB2U9+0h8M44iDQsINrcxDr1bjGBiIwiNjV8lsyJm5or/Uxoj
0C54smhGOUQe8mj8EqWsGO3THPhW6FUezWpJmSCqXkrGOWNBmnVEeeNB6eAYfPi4fCTR2XR7UNPm
GJzDuFsKt74VF4j6vvx4cEdrX3GgYXKdI70RUxBykGraxwuQT6atntsm3CCNTuYpfvCl2YWTnMsB
1J0SXDE2ddXl6RnhA8MU0oum+gPLFvb2DvTlAXvw2InS4vjQFLTxzbs6mV+9uBfxgNeyRZiWaLT2
T793hMY0epGJoargCeJ+fi7VuyvvVl/hE9WVRl5oqSFmVDV5Z7yViIebFEqCbmn4dPK6l7C914/J
DIQJoqPwBkdY5ZcZP5PfQ6fClE8OAXaHT9IUiiA2hRG769bDR5ONs2k9wSgVsuRuFvm/6Y7oEtPQ
6Sv8vPw1TdAVpbt/HA7hxghTdM+T3sC0cKt5pZrnfS2In280F9zO6x8kyXRRk+aB5fFOXRTw7GSo
O6W0Dt3NqMq8S+Olo81VeCpOeCeIAKHiDoU36PbDI6lGoIQTZYFKnvPjb0xWahidGfJNfZDbTF31
fxNmueQx94CgUNqFXYqnVjadL85nsO2ex2sddOiY2aCccOVpcawVQCA70f9HZFZUCK7IzBYyrStA
Zvx5Iuy5u8cJxL3wm5MC7n4Lk+LxZIG09PLp4MQ4+Ue3YWLr98XgAENz/O7w+LUZi6I3b+1nTg8N
csP4SP28ZeOJDjGeY7vTMfydh/ylPfqppFRx0TPUV32UMfMZKhSDmrEWKqM9u2bFqbKUsH+/gDs7
ADb5PTf0mK1nAFrbAckdxjFjCL+p86MHmyEmmcwvLFQpyPCidYORoLvy/N5KOzHCTNUkdb8efkxR
mnGzqddZlUB4SL5Ddz9l7LzMoXyz3U3x49Lh8uxk5iC300Wx+jKBtiK4tmkUSIlsLaRItwsHx4B5
9aa3TLXJQc0nwuGF6rVopNT7I5Ad8TiNc/Ak9dRdg+LBdeL6Vj/7wRujTTa1kNbs8j9QS3+0n1fF
wFx3usHxonWQo8zhbJpMXFGLc6ff6p6XcRKAEjKUA4TXHns5eg9oYaLuR8Iv3pc5NQrNDgaLM+yK
Kz94bfvcu/AXZezTf7ugc5a20sin5Me3mCt3AO9HETSxH0sXXAuoKtX8R6Bz+AbPua3Mz1UI9qcC
26vOYQLtJ9tOBd9hrVVcOtwhEzKmulTuOPTBwYAv4QsswqO6IajNXBKjLtyvEcatkPEdICbeWm7W
cdDsXROJwv8y31tuyKXBkG0E9YjeZxOws5Nqpaxc/KcssGKot1RhF6g5V9uoJhvSlQQN6AcYtCiz
08nCV4r7sH909pG0F2XAwwYXUbOboFKJiR6yvNKM6nrij2NjAXJF1r6p3Avmuejr7jhrxdeTkRRc
llPBzaCgOw8dEzOKN+benLrFqxufFSMmuF5f8sv2HtEduT6fYc6eOTujI6G6Ni2wIOR0gTmgH5ne
XIV6uBp2iTWliV0Wnyy7kYdzCJi0PX10t8K1LLkI/mwcPpZ16nHMS1Yk1YYayVjkO4bekzKEH8Qb
MnT0fA9XQlpukrKml3nu0FFvfiUdEWWSzQQpgxuvbPbW/L+PI6ICXKWtb1JXH6IfJYSxQyX6h2lg
HgJfd60C3piKQ7gvtU90RD0lGRpvmTIs2/SoPtLlsnQ4ekfEz7O/KVC24JRLG6VTCy41KG837Ncg
0h75Pzf7gLn5T7V8bTC8Xt4s1dwl1XLvmlxYbmU0phhm7KvlmWWPqfJCuSi5YMWlgjpP+8p8BZcA
HlF/xe4jVh/CGXCe0BrdqRy3h4PbhAjgkDXhaUd8Xay0H/ysuvUNV9HeB1J/2BgWzSuoVPR7FzHE
MocUk8BtqA9TZWsfL20ByOqanOWwZWHh+LyJwtzGHnSD26w2CRS1V5VvC0vqp6lgPmfQ1+gj02O/
WOj/WlEO23IX0ZjUeKR8ueH+qKa2OYA5XzF5qU3pAIYs8hQQBUxH31O5eG/uoq8O4itwIuhHnoTr
e5UEDaidB3cLXU7H1eHvwU7CfxNPSMOlivepFOMSgkCg/7AYFpaqvb2IxlMQDcn/+27umWkjsgEd
25s/gowkIV7p7wJsI/dqie+7O86b1z7aIs1ezRueLoDE4h3Tm/m5NaHEeq4bl8zbiv83EAxxK50j
hpEizEjVNCLrem/KoxFpP5pV+rBGMXNWZah6WdNPwShrQ3UPyjq5jjCj0Dj8K1p8I60IkzL3j9De
yRwOYyJ4f16CMh45buwwIjdzokXj2WAJisEeDKQRAekCMLL4qAxJhx6F6BDX9UqngnDBDCb1ZiQe
TXOzTO0x1X49sqeEOYxLn52EmcPl0twgEmecfeUiHvxoHkBIKvZ37HMmF+Xs6ZCpchs16rzXMASb
1Y6bQBiGFPIAHWBrpDpjcZ2mu6x/x2FQBrV2xm7qW5dfmwgst6t2BEqrWSA58BqFtYMShO6K22GB
EoHxcpTpQAbOc5ptm2X1NM8NfPtMbEkiRcnrl2eTgD3HUOU3JERuGRZDb+2yEzh7fsOQrsi2lFya
aMSNMVEjoAxycn+mhY/HbuAyhm0EACpdgpmCWHODv3eWJTbMMTjpHNslijoX6IMDmlWCzpxHceJS
I65Jzm/r0wZlivjU2g/xtWDHcFIfFtm9abFQQMGAM7zdLr4J49T5wcxPA5GoaC3QWXyV4CszngUb
KpuFOABI+JzPccpvqS4cK8G68YuPgmTLCUjNyjWBCLckHaKD5VXked8SBlwcLKX+VLKstvvh6u1O
kVYyHZhin3NvQC6AiOD+R5LNnq6lekLpHwLO8JijjDCc5N4BOQwMyNTVkqRV+qB3flHlODOa+LzI
ldUPlXrENG6Ol1duTSWX2gB4fJacbHThGqzLR+Wo+ZNbLtjczKGlp3GeT734LOjjro9SFpFYabYg
aDXMUZi1XxC8j1LD1wsKRTZ+Ldtva0bugrDUj4AgJ9PYw6EG6TjiGqhako7utMPxCKsDNnyAKFHp
510u1//NCddmDvjyH2zV/bPkErESi2DZY3hrvWz/rcX2oS8KXi0Y2GQXfS8/Dsjla+7Q4Cqqfr5A
zD8WeDxFLMOJVj/l3XZxUpO418T9ub49KOy1QDJP6qJ8iqW5ZvCqXDYRToSqN2tpWIpxlsP7xtUp
ee50KYS+u81mfOpdjJg9TdZJKxv7GGbCbFQDJYgd4HQZBcVIfBwna4iAnsdVmSXsB0KmVnFj3GDs
3Sw0Qhdz1LzyW5JmemNXQcTvPvzUpKaDnWoMaKpdO7suJQfuRtyDP6Gpfx5Shz+2WyetKdVvKWpQ
OUMp6Buzauf7lEkrusikYq16au3cTWahIu9TNgE8746woiq8DguidNaXyuflRMyIYiPUD0SJcEZh
ISbX9alExE0Px+3mlRs8kNtmwaYQcMVlMgDkU3Pc1/Zua4YvlJV+7hT0v3xDPCc6VWDBrJqTHzt9
SqZUSvEY/LF8JtjXT97elhnoHR3dbFxJnUVnvJIpXn2RXTzdpibNCWNAXeFk59Gd+QPCfN/2AE8T
GYGeEWylG+GFRcWs+3sJolkHHwlPWMyT61UEVf2b7w+Wtyb7Oe/8h/41JJZDCV5v43UCmrgnVbW2
WzPeh/TfPjaXpc+t/8f9Y8gH8HtK/60JaJNj35Km+wFLVnJf/S95R6f5xdoFLe5JlUt1Ui8Zx3D9
8C/M+m/8H9530Pw3NCtT7yZ9522TlY769OofluvYO4z5zcEZcRVM0bQgvwy1znWd3h18dhXwnplu
oCyZ28fQ5t6RuQcmUbDIM6cYiy3PYSfVeWINA53/5/y+5ZBXiyjhCXRCIuPhR1taBb+S/l2qK08Y
JR3TrVKtxt3Hadlt/d85v4UVkW8kZ2XpbJihw9OWZceE97/2+SW88MY48RPDv0IZBBjvOSJxmyd3
5Ulc5klfNIY0wveHuCv6ELWT44vVXaouDjeXwYHTAlkMNW76wtpZTf5PvFi6LnoDeEPlQ4FLbPn3
++r0P24A4d+kIWAPA6Cn89t8v+AmxS11k+WuEzjbIrXcO6TH2m/LHRHYNXjk5VvD62EuORTxVjRp
S/kncTPNwF/6FcO9eLBzEOwSfyQ02qNrsJvKcGt938QCaztd1Yjntm480oz9GUX9Dnyy8uOnGQd8
SsmxfojlBI5hXyL/QvZEisO3DgLfmlIfnCAmjy9JYeR5AoBHEbB79YABVL8dQOVqVk2ejIArH3wE
TA5JxYrstx/qhrpiV+3LKyCTptJrJ2TX1sPWkgfdtadbUE4sVmuEDPX2uqCcL0Jvddiwpo9jbiqn
svkzLTahUtjySYQx3+C5xU4baMhNW0PK7ZPe4HLazd0k76MwcPHkjy8168WJVBrACwEMwWhg9ESe
9/AmBJJj2s6OJHzgEK1qOK0hY9nWnBVnqsYGWJJcVTI+6Tr3XAKy0j6hLnHos4AM6A+R3wNtqIrd
VK3V7CLCBH1HjfP0LNMaRDPoW4pvOUX00JpRim6GYMUbNqZ/ZMkqqYlHU525ojFxVtvgTU/I+WET
oGr1FguVWFnFprV06WKG592dNTGLfhh4BngY69qGIrjnvPh/GfsK2FXtdg7O//BIIkQnifD3JCh8
Qllf27CamEfa0gFxnETv1gHZa3cfRcTViS51io3mv56/u2wrAMeeNbXGMtkGLR8bPp4XoZcth1Ik
EDX+2kn0qjniZA/ylQHdeW/zkU0WX6NVQv0yrxcdSC995veQTaBzBhGTXAjRjM8ywcbbRdeQVLCL
df8rM2JNZcc0BtNRPR5XOZrWcxEFbh5OlXp77M9vBDLIlIJe23WePERyGFNx2UeanU2EcNRvAhYp
jH8ula612ZMgko8SxpW3zVKvLPZOx0XHvfankCAE2rRqZl0em6qEUmQbHxZTyxM0YF6qjUxDZi0X
vEJBTQnjFmw9jDJ0qNSnX3+0QdBdVuNUp+qp3XnmWASQcxWaE8UJv6GY4e/EFp+4uJpJ0GbFGn/I
Ne+YGp4qfnW9undvmUhOItT5LA5liID/v0PmHH2DMC531UdipDNYGLfVSYh0FjQKVij0HjwhYLO2
qyh+sj7LHSOniRaluQeOioMSVvVUt4u603Yz5le3KdfUrWf4fwSdUT67mHcOAM2RYZkIZ/TG6wwT
yexTCO3G/tYgwM4AZIRp7wkRZZmd2eqea6dHHjmkJSdLHYCTofLIvR9VktnPBLIJXf2QPx223g00
CP3u/1eioaEJ+4RroPabr/Dwg6dOnc8Lxz4nDeKvFMLKICNPQGLLNnvK5md5MwfC2z4mokZAI/to
aRRG36BGIgxC960SvwIqGCEKyGadYKLLPNWqfJQFDwSC5WK/wK8rJnD309Z2zEtD5ReFNAm6ejXf
Fi3KIRJGrz6EhJbOskS9b42F6A7KSOXhvy+nX5i6iQfwEY+4vd+/h0ktrkvFx+8W87b10gEAzImv
2Rc13ExpauNyV5Ak343VvayuDemC0/8ECE2geJ9fsH/YqE407ll8CZIoat+yq45xem8QZKPgbLO+
xUfJrq/58mT+FCwY5mV4lfzFZIjFn/8x6hEbFm6eJSAmkTDiQ7IJ4/P16IZm7+RqYP/cSZ2Jifh0
NeBpRdxa6LOeeM/RAOa6B+V7wKjT52R6r7tANn+vPBJYulSy4vOyU6fAQ6gQN14yqpOU/EL14ybE
MynV4PWul9uQtGLZ0TgEkzuEojcjJ5x01ix13/v2ppYNIpifnxMZ8QrTbA9kAkpn1KYdwzWNC+vp
de68f41KbvWy15L99GoMIPcppvHFUZFH6BCM0tF927KrMCg1dmay4EpDKRqmoILCNVuKLul8h3SP
aCmJCdHamPUYRluXhUYPS0t4LsydZ18nwjLcHqatxUYNufsLwvys8XQueXRyoPEOSOXRuaZJ41Dr
Eb5nIWu9gm+HPS/tWhlEM2UN95O3VCLGN8eREzUNuenChfHNPq53SvAO10ziERWC6C2CyVPXEuni
ixV4WDdYr1pwfO0TmGHj60kbuW3/YNZXtfmsDKmmIvbY5/GwHjyI61TR8uw8GALgz8VEz3dyhQ4N
ee0DCigmkFbsQWT+jeuxhaNsYfRMlvgxf24fFHSQSltJvbuaUuwx7ZQuM8AlyRv7u5yMleTMe0w7
0R4x2Mr6nIielbSPhNJYTo+L/BJ5p4jGf+JrGuM8xciwMTblBzhrcQr83JFAFFeX5C3GMdqEPkuX
tBFyZNeEGve2vo7LMwyONbkWoSNY+LB677HoiTzVa1PoiX2iwIIhMpx0TQaSeZvbDF0OqT+clkLW
AaGb+KaZvlh91LQjIIXfFn+h8Rv6fHSAryUNgjljZqXYx7Y5U1BG2p6F2xb/QBJNuw0TsQY35JF8
aIfGEzlgKGVjm+NJoZXeaAkVrm+SljF4N3FxG6tFfggDYoXtMFfrFrHu3V4caVIdJzXh5ioOFtB7
ZoB3tQ6ZEAyDZbkcE1wbljg0kvRw++CV1VIWboTEchr38c4Hl8a1g9UekVFzeCRZGYTd3cLDa5d4
aA45UTE2cSATWISzDwSHmgf5g9wmK2R5HwSpPHO+hNrlS5emciDtFEZ9AGNs1s3zRuWbdqZR1Jhs
VInvJQIWUn/htlO+bzHZ0Yef3zWaQW0ZTOwP0EZGawShWeNRXZG1uiJDC7sKL4IfhhIQ+2NWmw5e
k9RDIBelqOW5A0nHJV2ZmQnI4/hXY3xHPmjmTs3+RJfcPE+NDyJ2prqhtwMVnvrIGVpVWoY8hQRz
j0klxwXSUh/mVPE6VXpImK4zFsG+IziFJ6cKVgmCarECTvbmm7oXtR489EfBDxibZPmmXEK3GG44
piXbnurcdsjmKfzFI4fHrljK4T6E6w5/B+mKE/59GBpgvBc+fdPPxVFu8H6wUNithztCeW/9MWaT
LiE7LJLEMVy9YJpQw8Fro8IwpTiCd0nrcoC6313zEbc1d/Q358jBL+NSlxXZ+dBqy/NAVJi+e7I+
UbI4TV10o3FzWcR0hARHvIBywItF8FnLfofD7ZephcYuVWGMzZmbWl1bxxY1uSIaijYtN/txwl8r
+ocaFVvRjkjjeD+fORR4lDnQTl6v4AmKQwxQo9wvuZhyRURX/I+VZIzO5NvGXZXbWZNpNd6aU34l
itcSe8FrT22szguSXOfmLM5OfvD1xNDIbarRcmltomp8ZAN8989sfBho1dRku60iQubZvBCcSN9R
PUa3HKE6cxGDG3dW8xqbUCNvpsO0acReu401qBM0S9KAm7QeCrNfJ+wYFqlWBEA8AtuFi+JoFFDr
pC9xFHmYJt+0kAlmBD7pHNV7ah+TEWgSf/i78laLsuVyNuM/1O9rR/hnLCc+SW6FRPDIh06xPn3c
+5hUti27bMmUun6LVNoOE7V9ILEqspCVSYWoPW6xTsOAoVVcZOA5AEUuHiRtQozB75Jfj5TSYCHT
oBk6dikhikisL7TAvvP2BmA7PrLVLzEibL13e5BaamsJ50WOV5B7FHct/gfvpcfM09uDrzxzHH5T
tt20gsA7vHOdAiX+uyf585mKgJA8SjxfScZHaCj8d6WNPOMF+OGla5dsnS/I8ZDjhWuTn+51fzPi
6Ee5qQqcAd9y3ab35voKvzEh9aNQe12Qz1XnmTa09cpEP/wIASiYwoxa+Q7CLvLBrsOUadIP9moj
wDU0/k7iSdeJIDWMt5zIkzuCdfYj5a1UlNWZ5MhXTf57XdICpDYj6MO0Tk4AwPzVZhp0s6fnXKsR
iEDgEtYiJj0oWVdHSq+Iq1BQdgNSB0rMAWX/LtaIBfED/FtHBF+9n7H3D/jWM0meWnoWfEO2Z4cr
zO8zjM4C/88Kw+wwqTHSDGu10ppvVehK1c19pMMwWqq5q2b4x/tK7hSi/p68K6tMMB13RYA0TqX3
soKvnHKtsKeQfcfK3XMrsRRWHBoKWP2jrlasNoZ0N0r98cNM8vnmfy9oBs1V9u4DJdkkN1of4bCm
cvM59jsEVU1/cLF+EamfchcSMWwwzOjTLmLA3biL9QasG1SNRuUTtDWHPqyw9wr+qjP0iV7RGXsa
wTlp2CpJCt2YzOM2YLg/T7he+iFHbmtAeZ0BtSihLrnRsoHK2syhFYmEUhrNYukiuqbM8lHftjgE
qhXVsjSCGF463T3w8eMXLMizA0YDbD8VbX9e15sniGAfmw/D/KfDzRRA7qiPZeAF0gs5KNrORvBF
eS9dCeF87uk7NOs0eu87jsHJcw+Cqbv8T8u+SxdO9DztzzKARBC58KlynxcOtvOGOE9DfIeoPDUE
ve/c3hIgw0p7UbngHgLvzdQ5DlcLWlyYSB1PaZ6X6Hy8k1pRFOieHwlKreS74n/3nXMQGpyeCzc+
61n+5gyjS+iVEmuE0cr8CdTWoezTax+bZt2ZY9cu2xi63UiacqMioNR8OBbIyqoVGhyPdK0oHnJH
bkN75N256wsoiNB36YlWXmc76PpcpfUuE1IJM27LiLtarp9LjFX9T837l+EPwofLd7vfVfs6Z+My
8uONDcYYnrGzWlNcOIWR5QwO+TCs98TPkPfhfvNlq8XezME7gn7vlyi9LWOxR8qeRYWJ9tBywTV3
Ri36UGxXW9Wc5HmoXk6/mJV8BK6tJsO81Ig9QHroZ7Wt17kq2s0m5WX5EfsEJOrjxviWnOc91Hne
iJSXBdJwYwCzhJl2y2SlVpeujUZt/SvRBfYzi6jJXqq6UNJZzVjMxfECebLluIr1iaeaORUCf1l/
UKyyh5mtoA0waXziO4WuXgRlC6KRnOF+teaYvULqXR0ifm9V3P1KPea6yiRP0Q2w74RAUsCC1FwC
Ss+98+Ddnt1RRKAj9Z57XsHwjA16dVmrl1yInQUoaIAi2eLx37ftAfW/OO1e7O1BWOSJLLXia3P+
rukT2cXr2BY0h6Vz4JUw2xKNKDOkV2HB9qdJBw1+npMPlWqCu4InRHJ+bhCoKXXrGlQjijW5IDNj
E8PBxdOU4CpI6GZ5kqJcdDrp+QPb7GBu/ZPYO6+l+iKccH0TEWQQ0rPvyLPi9ooyw492w0J+ev5y
ublauIAN2NTAoq5b6vhorRsUhGDPIfQstpUAEZE8UYFYvqFgDgciP5d+KzVMK52A6eMV+9Q/V23x
bdqafiHDUNnE1dzbkf5uCVB9D0/o6z0sK1b/z3zl3j7Fp0FTsyeaqbwITY1rX+bzQCMIAUSPJsj5
Kx54iGBzHuCI9IkAzJupJzlwoAlDlMCvoW+cw+lz4KnYhnunFR0NPd9Xai2jZva6lzExR5dGbNkq
OoiVDWC0Ym1iPg/MCCs1MvW3eQqt5VZISOLSNr78A3+rAjUrcEoIH69Q2+JTvjiOhVGE3v+AUDeN
3w1bkQ5Cn/8aibKbIqE+fWtKQYWXayFpLmFOQdMnuCNwSv3OL+2JidvKb2xs5D7uW0esj9dkIz0s
RPHJTfBEWM9BaJ1u/oGs9XbtqXuTLZXPN1wLsbg6NbjgTmU9kMoJ1Ou1Lmw9pWWAKfBpf7gGsTgJ
2ZiOz76J7s8oxxUjhTC9XcDyzmXyhL8HTKFtbgkZvouuCluCU/ZDex+TRaJLp6TxSQz8BMWJHq0j
S5NimUu2U8Samv4xE9ySUpYl/AeUumI8i3i3g3R+T8g+W2EcI93knru9j+wN16DaA9KBC5o0Bis0
MDzvE357FGJqxBO8CNHcisa7S6X6wl//5JLfjuAhgJRuKS1AxqrGUzDU0u6a2MXTuqEhYTdSdNBy
gL+PRcLj3X1Sx/z0pUekWfzp8gR+Zm8rBRVr8R22kOej+BP9Mx53tennkKYF+ZPWpEJEGZ22D0Us
TpKrgjACQEZB9EI6zwIwM+zd1O49HgQYixhUD+/KpEfK/zJECNtpjRRwbN3sDl6H7Yco9qx43te2
hzs7YQfjsepsfAEkkgTlV/FJ6MUXmnFmSu6cM0pFHpYvox7l2IrxG2lh6CU5UhjazKcnUh28m+NU
0Id+DrIyThRKrWqjlFjs+VnEh5umvHkpHdhOsb0+tz7MPJZLwHigQrfQlZ+U16bxEK3R61HkxEgq
b3ldb7RV1lebrqqpNq+asvlc7aQhP5vEFx2/zkH4XwRk9H+tm3ztGeVPAkc5giv5Ck1P6SANj1DN
SYqn8IDY9ETOMUyMPPRRAHvMXfR4E87dCeKdKBMiz2+oQ00m2fhHbslcKo4IZJdhKPclYFEO5lG+
AN0lJB7A60yK56SZT9tkEyOa8hOlBRTqEJbg5kN5eq9FEjPlSMgEpBXtmNeb56+Dpjni9p6l5bXh
oz1x3WgLchoxDweaoyOB0yG2rXj2lTYoymLHvj3itj5h9D8NCfjtRtVrIk5mspkewN87LezgsapR
pPNBF3L9qBRw8Laooqy7rIvvfip4etpL4FeMGL9gUXPXG/n7yo5Qfu/6XLUU2KIFq61A25x4YQaI
0lMrv2R6RKC34U2wSS4+lJfdkkwkl3IwJMHuq9CXCUR1DYNHOpbwL+Na8NDeeZAK5zA1Y8kCtBxp
pBZEt58bhecv8/q9pn9OiAOqdG1nehHv3Lj7/M2gBZ9Jk4aaWNIbQtOno4uvgeEMt/Yr2+TSA3+j
TYIDR6KIT5vPRt+8c94k4wXzHTKAY6iv9+Sx+A1OaXp7ab0WVZ3PkKmjgQNvbP4zqNeZg0lR03pL
BIQUPx7HENcuM3s+cpprZu91tLkwAjHM+p/8q8B44SNEOMkm/gOc/XtgzTQWbkGwbB8GRTAzo5AD
VfB29viY98nC8mrvSGuRSkswncq3VcjxwTRjqrluga+gu5BN8jTeGbMV88L0hsOUXi/hv/b8SeGL
4sl3vioAvaBbYBKAzcPWeYT+SXCZzEB6lcldurNSv4bJfJNpns4jFg7VyyJKGCQmf3htgUwYt/GG
7sb8JS2Cy9RogN4ojtmcBXsJLCHhVfb1MKSFHjwURaOHJZS/hC2J5JmycR3ZtbslcGSVdpSxTv6x
a7qBT4Wx800+cfGxbIX66TQ0Z7kw9RMPa6bBNsiRKgWBrTSWKQiBgCw4zbQ9rDEvUrd1uxElURV6
TNhElNOYttFqU/CWXFSAsAvIO2+5wAasJldSEuzGpol0lG/ZSjTlXD7xhX/q30sVfRzGHsqpiMmO
fD2Emd6AwQoqpKWPuAmH2MjQGjd2y/61AB38aF2JTq/CoPZt5LW8SUDFbcq/L/Kf2BcMwaZOCkmV
6CTUR4D5dZ4hcegXsdwA1fPXhtCqAJfGDDdlkH4iFtQjTfgwBt4N84WLuQgqhfBrpSR1l3KS55gA
7BBqyaYtOmkNVAdoj/42i66qCPKfsEx8XNCVV5hoVoef4gffry/Q9hbs5rA3dOpkQ3dWGgIFXn93
+vAqiy62CKTeehuLLoiiIs3F1EBVbVASGai/gdAxZ0vPiIXnC/2iO9gys7L1tw9xvrLGy8gxsh5R
V1cFDbluSI5+fXjXuGie0OoJs8hGk3u4DxaWFktFEtskWJk9k1Ds2saPCeTwh7gatRnBiXDCeyvq
JOp6EiXqbMn+sVCweCLQ70zaoyX9mPUEgmaHkQcQ8F9MBTUUiKizz+qXpd7oACIn57IyQDcpC5rN
/k6X79d+Hxxf2BL9NNxzxCiTwh86n2yzPo015E5mQT9rebh81YQE1n8k5f0sL++DJHLeLiIFzHQ3
/Est6vsEyhae1ZjCTTqjwdpgR7Lm5mZ6mrOtII2F0jccWvF45XerSZB9hgyU8j+aEl2yk0mD0O9p
edIZUeHyW5xG7XiZnX3n026nlhbCVvIQenQnbA48v9/B4M3pjxC+KlmbaHFVbtx9G5BfZ0J8PU94
b9K1nMQFJz0CqR4MJ1dfHeGgQB4AHZfJ9xhnadSiC/6ZAN/ewLxQBuIJFaxG+oSST2E4nA9yPopF
58tpoUytz+ZvJdINi+3PLCnyh6zLQyjZeBp6bjVaHrV4ITOSFun68VvJK/Kxxuxes/fH3QcbQPvy
YWd55q11WqIkjidDKBQVF2vvYdGI1mhpBqbOhsdGYS8ZzSfXA643xwDOt7ckDAGeFFh15m1qkOYt
9Cpycmtb5V//DQAKIS5iS88y4W/AVysgwLHPEUP49pJYGI/Z5L7qJooUm4HTggexARyocglrjzyU
+n2l9nl4TmEeL5W/vlXaOhIwHVVBKuYNa+AgVLL5RRqcOifN98T7EAxMGEWI9kbjEjnyJ7yQjnFF
CRaSuPsptljB3Uih23iz6BRVwgtb3kGXJnHddAYXqPdSDZ3LoAvPHGR9w38cQibjIDiX4ReJwjCd
t6UXnCj09dXpcr0Loi3twGuPnwMXuUJv8f+PL++wlaCO6Pg4kTDIOcj5kOCfc7G1VbUuwaeEHNmy
NloeCNG1CbtYf4m7esFKILnGqlTSWuoXjU8fyMNMbHZIQGQlil9cL36gD5cm1YgtZdmyKyvx4nqf
psACa8jRowsUaN3DI1Mv6RpqumaOvrLXjKBHLqEjSwrptNhnQ38PSVTyqKU9rRTc5rzdKdyGznFI
qTfzF04aU7TJulje6NSdy2GcbHqm/jQpPTMaOXs+Q3GlF0iqhVUfIivgcAMRIm8kEGkcPjm7swaT
WaAvR/7QSk0oSMu3biPn0xWoUoaN13bITL2iWPBAZeubLX0Odz3NCCPTml39c73Gfcd2lJwNIvIn
2ol1idXfVoLsJGh1DGsoJYyzznSRNLPGjhibTEY01ma4L+0QrrscJILWP6H5gpugZ1WhN0tAd30g
SX2ndsD0aAy8OSqnx0mm1O1VoL0RjEUsp4PMxOUNE3sNuENMPZLal+FXNMIjWR6nuHmTdZVNsDWZ
lOUk5aYevsWeKLdatjaXmIEsf/q8QyeiKohdwCFZvnOJImP5ugP5So5RF288HhX6Oq8kkrKkRkrv
3MhocZ5LYXc54vOFVxtbH/O9WN2N7dhEopO+pfz0roBpHLqPsLoqWgCw5dAJ3LSWP+vjQn0tYMvW
KSFLo4FpU74k/ZJPdqfDun6YptGUqmZ+n1qof+naAAFkg06hAdn/quc01F1y7xz1Fi5R5Qq+BcYY
TF+nUcbNAUqVLRd39dGXPEDrrOH1FBhHLhcxu135Rh2kgTzPL2aOPqXj6MglR562su4bplSOP6Dc
62+KK+OIU1mVzQBZAzxu5PHalwaMkwkx1NlbEobi5l8U1/AaEcj4pyebfk3NXfCXx4Rn0Lgglg3R
GzYgjf2Yn6sKMKS1ZSdJ5Akv0K7CutyKW0fbEsZoQeQ6DWpv0imjNqyN/bb+XDInGfZ86r7B5/U5
V2eoU4J++Psda9WjVu2RdpMTeebvzT2MMW5f9hIqlsIeMswB/Qw/7mqF+Lwit9kAd4MgQko5DWCx
4mEqMn7saNjIsY/BuaLaiB3bUzFeijN3fjqKH5cPz+G5aqsAcbS+xNmv55qOddxdVoVov+H6eeYU
5RyDXMcAlFi+CBVNGYjKc+xkxD3E/BMP0LZMOqcOCM1fakIK7n8jpkvKNfNyxrEgi5JHOth7UeSp
gPhnXDjzPQASd6FknXiqJK0AcDb5EvwRwtNHNFe1iTJQIhXIKcYP353nRQ3PNAfJQOej1EZhqYhx
CfJRrFHrKcGPkWx4P40xtk4uz79eR3e3+TjVlxWB9fgl+3Z9DC12H4EaURXg2PbdWCIfWd4YR7cU
X04gIuXE1SaYdK+fc4McBkoh3xE2GKsK4chkjAk6C9ZPDWZM9BctctH9yXdP+5m+InpQNmma7CLK
Ho1KaxZhLwLX7Rce//N0ItCxpCjRaBwKfAIqCkTHj9IR2WIFR1JZ2vIf1vV7JhBLXcodKDyx2GYn
kl/rfUiEQrN8H7I5UEZ7IX3r7LdY6749tlvCWe8lDaC0ez9SW4sv3VneCoeprQ8zcWVdZoE45vTr
68LUNMdRVHbuk8WplMWgj5gKJo2suivkQOLitRxDsJ/ODpjiH7A5J00uaYxirS4YsOXg4z3Md3Ze
K5KD55txjqPK5gEQ4qDz8fQG2Mv7hOjMJj7L+TMqB2aKr4a15p8avZcSA4Oi3xrK4KNYD967qyml
ASt39SKzkcRWx1as1LnhXPpHoAs5ta9S7lW+DJGVP2QKH7rqHMKium2TOEjtO0PwXa9VHE4CF2cL
rmub+emYhSaxSYuRlzHaTsyjccs8y6kkgP3e/qxg31pv+Q9MbX/q1Ff8eE4QP1cxOzvPk/XjnYA7
BUVwV2zYH0mQYwd7cg1GJwIoKwbkeyY1JX7t3YotiuVTOXicwyTFcWb0TX0vDy9VHJn+B/MOTUmw
zfNyxJvkAVR3rETvooqVoSCkFN9olHb7XExWtAiLDFEVjjBfssCVTZbaHyIpQemoBOVyZDMQCei7
GWpkrqZhEeMyVe69vif1I9zj4DTtS/lUhdRCKFfDbTpiEcWCeEEIWDvjG84/vDW9B+gWX/wRKL4o
/ffhPvhroGJwI7tDAtzb/yGWPsZMeB1lUKmliNTGMngglB6ENcg4I11htZfu40VFr0NlAJrqREcx
2BDprWcSfR/tK3c7tRcCzUiI5PK6eMSE0jT9LV9YHZ0GLFkSknT9GeVJmf3Y/I7koEvcEwTmaOmE
WWpOyi3GEWoUfi+LMwPyARj8DPyqFoTzfvqkgD48DBeXAh+TPNVhgTynLQ+AkVi4gqDTjfCrtd2Y
qqdjVjCXENpvZQiNZinSXyHlQNIGYmnbPLDyV6vZKp9GinYiAq7Hbmzw0qiL+8gx/YrEDJNpuoM1
iD2dl/KZmQI37VHO2512m43hk1eHD/93ZYIgXQ3rAPx7z3178QgS+O9HYwPcUhyDiwI+q1IDOEkJ
i2UALSbny2VigbTb9tdLqoFiwMtcAoQOWtnqPTr9XIL1+tXWbtn+tnyr9O4ma0GCNIfe2SdI3yvw
FevrP69h4OBXUA5/OETdCCLRlCaC9nbvqN29SJt+yo2SCcfwShz0FI/o3YK8VUHW8mdPa2YgyzeE
lTSvCR69t4CfAI4yOng4G6CYToLT4oNcv4+Wxg7TESxRY2c7UY+qAnpv6c3tFTiDsdExuvTmSw/l
VhcvCRXUlFW3vzDDCIbAwQjIq+w5LlK+S8q+RSDDv/pKVxAJqhHJp4dt2zuE/fqEfG6Xdyf3JPaV
ZlQ4VnFAhO10+LYDhdXXbh+dea8s6woD2zq5BXRhJimlT6O7Atz6ZJF8QX3mpa3/PT7G3+V+Ld11
Vh0k24c1mWf5RKLpYZmpgaWq8BBZwDDaiXaBuxSNM8py73ZnEh4aEIc/LbVdyUh4Yz8SnfBDh5V3
/TCAaAQo3UcyZyx0VVLQLwI5AQ/cDSTUDJ6GEEAXV/5zIy2gT5i+ZvhNANh6w9kTTF+AlWk5S5I+
sddRLBMRSxape8DSMcWWGv1IQ9VzpnyZbFsbS2euGPmlj/00TnS3CAREh6SBOSc0JQU9QWSi0OxO
q0Zw+ehTuWvPxs7OmFmYbye0YQOcd5RWHgdH4c9wKTmFk5XLDd/EyyYqbBZuwlq4K0LLTlQMqclu
VqCm5D0Oax3dyn8u41atNovyHKuRsXGl/B4LxcxwyZT/jIHIUJUgcZ+azhw/AXgZHtFBytmXaoTu
7VOBaHP6GmK4ZdTfo+IplARMzjLXoPc8u5Iw/auZ+kDRZgjn9lUas8qnqU8MUi6IKeWcu9Bh5EPn
RWuK5ybfjACxXxtQneSBVBt92bwYOwKckBRC6GgHe6Qse2LeJZv/edB9tHOftegckAPD0/DuRWe6
0wsDmDOPaCnc5CIxPw4XoFfQkXnGcnOi96xQnf0wUKBQAXfRCiuakVcmWWwuZa88pA/dEOH7KLA2
9vabPfUYqAdhpHSrAFVe++sHc7YULc8JPLqhMj80eXUMM370NhltpCymnY4TJyFi366IkSq8R/Qa
zqGTntyrEHtWcWOxPHAakwhOVw+C6SaImJhA/dVfrccarrsHV+CTZO6SyoN2vdFAhYF3fbZTkP3f
7Go70Ctxr5NuQGrSVF9Y8idalQdFdjTmxLhury2/tFIMESWrGfDa9Jg2xv0hRjwQh8Lzr9TfIGH/
dAkdrR80L8yImVFFsOlcqkYkYbC0I+Le+CE/iDLxPQoB4JQG6DysJxWp/dZ5/l0qg23D/SIhjwZH
+DDu0xMBfvl1e6/AA6WgSL58dw1s+hjsHC4dRhJ16UlEFl6u/d6u4UQ0mdgoLVj/wewkFKV1fqx6
JR9tC5lSjVFgH9ovtzRPLm8vEqg/erCyf125uWR/NdOg6/mlLSvp3yZ9FqEi8Wg7Rys3Em/UAA1T
9YVIV+ikEgZGCoucUs0NnmyAVB0FYDdLiUF0kHCimd6N2rYW72Dw/KNt0hUtT07Cm/MwM3v77Lbt
enon+fQr/b0pwir8nBa4VrAfT9STdKmZcdWe5OhWlDdm5XQNVp4cEG1Ie941uly3MQhgTEozp++8
7tMCWwSVAtLrHnhpxFHIpFXa0W+3E3A8KFisU+WMWBX0l5Of+CnvaOV5XtJ4cfjOJSJpmtcIOf3l
ayjwIHkJtmtk55qDuKGO8EDdHKf+POsJxK2LKqe1QeKJCvgg6nsYNHDxQrCIdCD3ZHyxzRH68Qhc
8vg0WAZVSw17TS4irfFGN2EADdK5ipMfJc3fImZ8dyU13lng/2P+JJrk+e3OsbHjiLRBHg6/l51g
EP8C7iNbf/8k2u5Yr/LJHLErwQJG50T9wX0ix9JniLSzxvOz22CjahheNiXNXDhvniMipGUjPIH6
+UpF1AhLT01GpwP/TrBrMcUomIXuJ9S9jlTteAH/C3Tfe+zEHwCpQxjGlSmmqETe/PN3hP5i9pCc
dBt/7Yahccztv0EoakfUeFKGM/V3A+tbZE06ByHeSDs1ABCluSEtz/qqpJLU0icB7jbcfZJ1li04
s6/XQUPhWmNp2Cg2jU6Cs+ZDse7A7Kk81hz1MmlGn+s/NBLEThrWgGDyJE1G6ppub+Zc5ji28RUY
jHGEy6sQhSJ2hXMAj5hoq+GYQUdDUvwvVtMWItN12g5buJvx62JlLDVCzV63eQWcPNUZ+eLSHBQL
QadNovy6OkpI/zxrZAwiPdP764yay654r722YCkOrne4CWupclI57Cy+v2QqnqmmNobETKQUS0LP
cb9gs8N49rmXmU7/kvW00k8NBchComejM88ZmuHYLKPa31qqvClk/hTRkKRIvLBMUuoryMQh22WE
sproak8lVtYkOxdH1A27Es8yTq2PI8Qdvk+jchg5v4dDFEEc1tXNf4ceD8Q8M0oYbScNbVe5tQSt
qMG8WOQCieGvuhl3bJ7QKYkRytR85BFsh8Pw07BmUv2j/n9sedCXsHXANes/pvv9wNYPuaRkHPzW
/tr1n0V1jkWfOnZkWhyZJpRnIU4mIuASPKgZR6OSWO3W62eO/bkLJ+Helq/AQC1DRldhsxg47GFF
HbbNHumPueGqEeVUhYHDFU73YZTzyy24dWjDB1TfADZfTgckuHjaT5LOWyl4tN1/wEPEr5EK6qXx
vnSAOZa4G4y97ErRNi1Hjp4PKeh6K9N3n3ostNbIgfN7h0umJpfBtihNUwcGhD7IcClI/QQj7+e9
PLPRRJFsOn3RLj+V4amxM44fFhGXuCamz+BtBtR9Rb/JqBhHCSzB3OWabjU8IvDkwlM7ud853qdQ
aPq2ukeuivl7RRP/RFL24uVImwZGx+2VyMlDYzQT8rAod9CBSJxkoZc1pcx2z4aWODrZ2aF8CpZU
sHWdYDLvzMrkzS9c3enm1blo0KtvlKvS/MNdyCkpK+vo2dAyDbX4PjCkEGL5xyqwq5cryiAZlexv
n9To8E+HCeUl+cN9HbgfHC3iF9UjSygnwsf9GiADrNetUrnKvnQNcyu7olA0LYU6QUishekYrVub
LOWa0Pn8xfW6rqjfz4tWreCLBbTvTyKFQgQ9mxIcDTmC6seMyWPy+MoAlJbvxXrdkWRaoRI9THek
Wg1xQk2AB3NxwLcmEyoMiaNWyanx94ZYv0qHC1wFE4Dj+qa7k1MLZjpFfm78mNnTGThInN7+hlLe
fNQ0jtgkikUOfxCKgi9MIJ4MbdnmKmnCspYvB4aNVFb6h+wH8B+b5SuG0txyWvc452ZjPcW8HUlS
UJRs/G8+svoBLbfrcRxRPlboiGFQR8SlxSDSvodkAsi2DdEflNhmpVpI8weSdlPaD4OAhT2ABx0a
Fs3bf3A2v2EftmNaot2j7u0K8ICWzdZEQyupJs/wxYDBrQiiiLFlb0pz3mP6buUU0EiMWVae+Pul
Ss98+7Uiu0khET9/HDpbfDTOzv1ngPoFtuHMbLx1gsXXf9kzAmRl404+QTFAi7F9N2vT8cDE2Kok
siT4kEvyfRHBDZVEoYrBsWuAFg8fUE41Q0915cAJVBus1aAbHuLvMtX7+XJhV1Yia/hxaqoMYLiK
1aUMKt0Z3JCkqn7mmHnspZy8DS1XwohWWY1qfPE4cUoFNtjjFpPfM1gjc/AfYsxuYcw+qJuEnBCx
J+MMiQnLWBy7kI1rD6TRwws+C4bEpIlFY3aBS1ifoq58cORdkqyOhdaS+bcm0tj/qI2d3eBOcKLK
bP9ma2r45SWzW+NiPIgHq58xd0gjFfHGi2Qh6yT8X50rwDX/S0iOOOlS4YonyQ0XSM5KcmoognRn
6b/S2WZX/019OaA/U+oO246KF1TwWrLb9JZawf5u3lEYZY3XHCXdfyEcrm3CtlDTFJBl3jc3lfHF
yg1xRaOPUtZsGeXoNmCz3q6e0OWc1BiaUiHWw9GAK7tgMZkszxgcmpPnUoTyUYsd+3zLPK6ttkhQ
kAWcHcO0flwcTxRNg58zuqVa32uPsXm239yziiUo6kTekbNEG4kZcl++S5uoa+OzFqT2C4/znRRG
/KrdCw//k2IbWoncR5mpidYLXV8vUH8HI1+QEQhTP1cD7GGGiP0vMgu/bwU0WFaudEf4B1Np3O15
OfCHuNH9gKZMEysIIM4ej2xbV7I2/8Z3+F3HvIc8CLfeBdbjzxd8fZHDeNxIu0HEPnOyauCVlqSy
OHq8TEGve9Nx9z8/0N2ANP+bfwVVFvHtIOFCLHjDVcMQZMAjXJ1bEGSGOsDRmo/eKsZ8S6r61ImB
jkR8DKCnU8VwPxa0jki+QB723p/89nMS2Vp54AnPksdtBgRf9+ISjYJw8jOCAdkLAa95RhwaaV5g
NlI0w9+idthcDolojcgJO7OAxZKPndeDoJDI5HKRLyz+eQNTqMxCaZJzP/t1zQcroDE5h3Cvy9qr
EY5S9TNqOSj0OSP4io8dbkdeG8GwxnfrZBSqn7cVhou3w+5Bl3VH6A/ijP9LR10cObZNLLPLYrYe
R1bOMsxGFMXesdRYuVdXCTOboygC1Tbx4pnron0fSN+0hzamMgHIrLSVV+n7xmBTQPUC/v0vZ5qL
s3dxQLP7QC/zsxRy8LjhnciCRzrGgjX6uMR9cxmA1LnTo3eWiyxPwAFlEY0vak+RHJXYKPgGXjFA
RKlCG9wKNMLtFDZvtAEZwvtN64ZQNcH+eY5B5IL7lEIEJMuxGqpB1VbVq/WDeGE5I4P2im2MB4MB
iHRlI+fOuR/oAV3PCZvbie7KQIlHaOPblRRBVyDFh0kTPjyXKcjoIKAtBiBGBqsJrssfQgRSzCmA
GubY4zSUUiWY9dGDiqFs/CtjhBc6Ea3S1/KMXYviSBeoaAV+okZdY8CiGYzKeNNDHOMCATaXe0SO
nFWnwisSEWNEeC2Mr2PWIfCZ62zrleWEYmYC5Ukr65AVBhOrj4lDOxblSiCwtxGlSKlk8zrcA9ot
Hthul9lA2o8L4ZAKXN9arFJsB9yd0LZ+WkBuXAvohhEvfz/laBHBViQsgJGywHJHV/RSuwcSiKNs
Rk8zhEQEDDlalsPRSDfZvIkvuY6Un6tod8NQh80UqOVHT9RSxwv5ujm/vvFZ/Oc679gAaOfSt3Jw
2hiH1++l5bZUsR7qAWiX6NuGvVLoksTcQtlBOy4LawKZ11qTLd7ysjX3NnDPYU7ceYziYWZlYlQj
9EwbYhGjjCtByXLrCxibAYhPGf4jCH8egQG5OdNf9GTYDqfhdismvpT1OMIBtxuV5L+0PdzUAkJ8
QQxkeVIFP8BlOM2jP0JKLsaSgcbJ97EH7tP+Odfy+YQ2ns2QpdLyDjGVMPji0dW0L8DiFIyXj6ia
FPdl6t1xsp/fYkCEopuUlIlAVIH3+H8w+eQyy3KpBU5qy+UDVjAv/W06kH3VjJNZY6KxrZPAb07h
dkQtAJspZH0bYiVEe82RevOlDHtaq+jp63grLUScTLUv+xCiRbFW62GZm6s6OlYXB7WKrmSv5d/3
9AxCwLV4vGq3Yko+N3Q8tN9GLF8O5t+n8LjrD8vLxnMGgG0V4O858G7imt+rvarBS/XGzPPvP4At
x19/mDm4nTLvv1uOW7+SLCglugm/Hmz0qrA+DPv3FRZHsiX1E0w11t8h8V2QY4GgUXBXoLPI/5IT
krTA4ZBnRNDKee/XhKa+yAInmVzLErKKnT+Z4PFgY4pB6PlOtoDB7UE7TNpxpu+heTvc5gsPxPSC
st2lRs4Wn11cHzdYvA8djofVIysqFhLIgggiPO5RfVrX/VoMHONm5v8vC1/o80UHuj3SjSCqNnos
zrwW7kKIRV4lYY4+jqwb1OsPf8b0GleEeyBNv8nA9ay4M1vhdofWpDOFk4JSVfIreUYDeoAh3if1
DnbCIQ5CUs1l1oX4B7qi9YmwjxTjGuzgTW1x6tsxT2yc5sH/P5VekyalvJJcjvylUWuC7GIV1QKD
Kd+kpIyOokuq+3MJYQivJtFZ00iatYI0+Ko+0mUAfx/cZlpxNGIF1F7oJv3QDEQBG9B8ceRNcMhL
mYWp1HK+OOZ7kPSxiRbT4s0JBheRv2ckcpTCX1vjxngn6350/c057MSfed8L2Rx2ptTnG6DK/LBK
1wq+r78C4wvowNBt/f1MB7LCBTgZWctjKL64r+hsCxlK9eupTn+kFxSf5MtbLBvcZFXBSauWaKtf
HMx+uEOIbW6xP8W41N5BJVnPNA+OFjYCnuC+OtJtC4LfvV92onZadya5MMltl96d0MfxClz5lQlV
U2iFP+t1MiMhiNG8Ocv+cm2cmcfe8mlzLae7SetRmVrp93oDO6nMfljE6Zuo8+HRL0VdYIgITtpv
iGtFSD/ML8ffS9lThc2kh2yCGxvSTYA5YfTDeUHKlzFoHFPIifFb7hZ8p3Tuy9iuMQVXBciupgq0
nWv++mdEY0WS6yqpghhAjATxHs/GQEUQpYYZQcpY9imXYAXwJmvYWNUuhIppE80x7d8w04IJRg9k
/eoB4OwJDe/pVfKJYyrrQnhMKqUv3LBAZOJvFwz3YQWC+YRdLTPzDb9YgVTt02ECbHHMozlakW4m
MxQbR8m9vCXklq49SozrUU+rKpJ8rTlFA5E5iw7gcyzMXAc+Lg2IsV1KFFj/ybXf+kqnxSrpBiAF
CDGLymoxPVvQuJXz5ZsD6Z5SQQ4eWBpav52Yrv4cFzFIuQls4nlaelgGfDk34wxRiyf9dV95WAd4
/PcJZOISTn+ML8KovbIpXjQlc9mFyTpx6ICpqB4bOuOo0Qp/K9IeaQ1qG2peo5IqjKpPOTUvH+UM
OwXTcZvDXY1lD/xKbJLgCSn43owDMXLXO5feUQjnCVb0JjgPuGlAJTyoP/sHbQM2Q6in6fMCa6n/
W46QgM2biBC8fBtzpnziM0jXV+lOafEHy4kH5DZArJ+7FY4AlepAW6C04LXlry1akYQxxRcRoZa4
/jo5dneYs+YMIkH4KLEcYW8HgW+kqULti6W7uA8Zz+fVvdVR3cD7YY6XrmQVl76mVGjGZWIHIGzI
JirzunVmBhnb8+EOU5CSzx/emkMnkDP3l4GTGaTcZFDHpOIK8SYsJVFcXoA/J3ENWltDO08Iopnf
8M9NAzCq2qvyphiDvVnoldB9kz7+5KImwXh/RUT/rulN8BQcsaPFiWb01iEaoaRD44wb3VWzmFUY
HintncIRiEYBwgO+1fBU83qepAT7XUi4GoYL2/Dsvwt3FshXk1s1kHXlCfn79vSeov31R7sSbc4J
8m6HSyRszdGFW6gBFzfPqePvSLobt0CNcZ2ijCOWFmAneo0zgY2rqmVkGPgCdhElX8SPCSY3jd2h
Sa/Pu+euspkg5jYNfqYZ9CPP9pi39WsharPTKvF8PeLB9VkYU1JiooIkAxVn3c8YJml4x88AGAMu
K1okbKZ12JR5kfKvmpjhn4JMLZ8ummBy67GC60b1iwu9Eky/i1oHG+WlYqtHnpgUsQHpFsgDLbFK
SZ51zUJG4VgEOInWxv/JWtpomUId3SWf05F3VkBcczdbGO6MmzsnLQmxqxnMlDrIh6wMKpqFm/1H
vgqa+d6vqh0sXA+yddrcUFmaVoxHlD6Xo2VPxJPSW53PVmqAdPOEc93mfo463won5cF94jqzutIB
d0+lkvv9pRcb3j2pAOMX3dThczH943boOYAk6r6q2DTkT/4fPUpL2C5+L8+oE61azXqZDBb+R2Qv
ttJefWd75mWzSDP3HfEFwUHCwp/fjJtYHtFrWNAs1j529krPFJLFLaNF76AkI1/HoEOENTqwtict
A7ehKx9cffMEQ9B34+Tz3aRWUjq63DBLcnjdtE6N3zupMq4xd2O/33FR8iNCWVPfWaOpvPDWAySR
uKEmeNO7U+MsI7QzmOUJLFp/MJnJMi5Cf3hliZjN+LPr9gisuQzRYruf5UO12wXiFfvHNwgLylA3
tCZ/guaSCe7OEK+OcBmqdnr0OkI9ovXepQcsm6q/GaqBzj7yF8jvk2ipGt2k0tI6FLJEdOY6lRyV
AwMxxzsgVU57ZSgOFK0a586Wa8gHDBZ06ckHWaeO4o3FHP9gdyxagLmflSQFsI7uA4BQE0a8pIIb
OyteuEa7UAlR9bzYvLJaDkbdjBwi8lDLxnchqREzl/510j8COtvY1HZlNJFkcSqxEBGFOyoB+Sob
jYYpHo3uC+22DrZAgHXu+YoC5aQIaFSkjSrzioBJvGpNaoX9GO7XU8+pgUFhA1iHwD8QL8FRxGbe
PVeq5bqfEUJyyxQWk/Zuwgue9/HvZMD3kZgN5OeraP9UP+KheK1mOFC40Fhp4fLcKEgBVeYrky2z
mTbN4fuSWwurKOuEucCVAYKAP673rI2mz+YydAJyO/Fx4GM8SH/znd/I5bFOozxcp+jJ0jxYk4o9
eirttmltWYh7sFvfj0fZ48FeToH2BZc5DcByvHNavl4yhLJ688CQXhGTvEM2h6d/3TdFdl0jLldT
LEe+SqDnwndU8gGT8RypXRKuPXkuDmBYE6YPaTxZIuPbvpB7V2pNaSeFotnUuwMgiNg8NmmKbArL
+Nn8+ol4p1w8uQnDrp/jg+kHmDYXB3U79fxDr3LScS4gYs4Vkf5Vm4uOKQJTb3Z4AbxzYbDwE9hV
HgXTAxIlRLTCHWj3K43vNmSCXqt30reiQFcfWF4xFgFdcVwQpxddtxTvsiqRYkLXB0pLWt4MhrVL
UAzeucZFjGrZYCeCmBY+URDcBZsUM2e7HpYZdVbUIzgzzgQkBT4OxDYuaAKKXB8L5RW/Xwb+yV8s
2pOq/WsKSrKe4IS4dqVnM9V7OoZJIPen3OGg8WWXzkjBcJhUiYAWZuycVjL/p1P3SBPmB3juJP0o
xw1tg49EcdQPwKqOnntLV+UviziKdJJGcvTjmeLxXff+AIBQLxVNeWv2lcyHB4EY1TTQH/TsaWjF
BDtsvvTEhcEiyK7AnkhNshzvPGdqb/9Z3LRDBSVXHzBvQWcS99gtwEwYTCrQ9RX9nbAov8Xf1cza
Dn/q7Mt4wEk6zp5Kf/13CXq7cFkCXv2Da0Z69j16vVPzLZdKwJnwK7uamGYxnNLYlZ8sB48G0SUY
DPLgY+TtdLjoWfwW/MTlcwFqMz8M1FSjHQ0RLGy1yloRTOtBIpLdUixZYi8Z6sqRfuQfacna0ybo
/BRQ1wMJgwpJaWlLYs3DLBaGMhkEyfQyNin2ROnKMcObXgeNedQWzOhnGgV7OyXCAv3E4sXKgysV
HyERmMzylJe9uF0bipfTvslQd5lgOReEIF1oNLtrxWROYReBmHCuu4M1jrap5jque+KLu8l8IQYz
PbbJ4fbQLsTxKfS14TlGaGFAGXQ42jRrsFb/h6Q0Hw2ZejQRYToKQqoFM1a/MySOOTzQduG9rnKP
TCFxJ4Ky4LBxmGuTgMZ7BC1JcICYUl3EwgglJvAGvgx74cG/2h/U0261AD6Qn8Pfz6z96pFdEH01
QZys4oCZDbV4ijZXwz1GlGMgNrI/IvpIeWi/YrzbkzRw4j48XmXZhtHfZgDweJvtCwehJbkUixph
BVJ34sY+gYlkMVEFN9aG5+Iv7MejC63OW9qpQWSo8lBP1szt3L4g69U7QqEpCTszjvvQHWmk0yVv
TYMnD8RX86o+pl6yDZ4fQRRIzvnfa38ppetNTXTsiCCrlD8jV9BQ4fCmkmk3KTLhVSj75SaAMRIM
2HxsWU+q8h+jz+w9tuX0KdwzTV4eQLVjx3bUu29TzyixvYHHOWvlysng0ek/PEnFw+cOM9zeOzsQ
CvMgYzcXxGO1iom6nNubdtNKgJNpwT48Fi2IOsF9Ts0pSP2HlZQTzjua1essvtkWZ/a1QbIHA21u
ukprfgqmhrfqmwxWCRJ2xsQvQfYvIf6qloX/gf18/2v4WsFP7N28MFxiGU1hOjRkfPZO5kA/G80j
/X0VuD4Pu3HMZ60IIyeX8R8DF0++bx01tNBu8M9VeiM59lUGdFaRxINkQpggf0XGuHkkPJgvlGk4
yuPp/Xn3zFkFDmeKvLBMS61seMWS476DJenvvWyJNLeU4pQEof82gUqEe3zZ0elROBu7go7YGyzl
JNFDVPzbApoKUIUguahGEyzu8B0yN9OuKrccuGXzj7eyMxpAHmgrV3iu5DSG3glf74y6Li4WvGQ9
BkQPUuCcARn3/+E8hcJlnKwXcJlz4E0Aha9h05tPcptjSGMiW5FmA9V0EEMb0dzmJsyfGjszd4kk
N/O245ThAGV7kWpr0fG+afxAvekVUWblMMna72cdY77vkeSGSfeZkbBSS8HYmPxaiGV/KHIt3t5K
CcgcmoH4w2P9y5tMl7sQrjffqfv7bllwJUQUe97Yq+ET/Cks+EliUqPGZCC53G/gwutyn/adO9dA
C4rpKJAMJONVlsy3VMRROyOtQPpE+NL+PxpLRGUAvabVStPo3qe80SCnpD5/eczGqPa+Dzq6pPBj
d/F4qihN/+O3tQpeFxIIeBuiBfR1GCege49f3L3msgnh8M5M+QMvn0KRFiBkICcADj3q7PFGArdm
qv73euFhn1DBEL1Z9m+4QUyuxbW6nKqSjLyiXY1pgNvc6NYuMX0hh3dM/eqY7BXyhFDkPm08Ojt/
hSsI1Mcx1oObGGcphhVVNspoHrs1YblhNxYw6Xudl7uv6RyFZF2LW2bc5rNHIjQwppd5tM4h/Qit
G7xavzsJZxpx1Yrv60/Q3TwJM0BhVzIIivZKWH1lh4LdfWzPrPxnT7854uyEfnUA0MhKzgf/lIAs
WPlkYu3kL/8dMXmHaknrZA0uudR8BT0W4AAL4ECgHderntaZzf9ZUdky1hjlOTSxqWzlL4icpny1
iOXgAyxLm6KWWCW9y3Mj9xEPX3k8aNrFVQMRwB9txPpgCXShzmbu4wMSwST1mCm4E+TvoUCacNQx
rSgUIH7Uu9zc7kbtOUlCfSDOe/nz1huZ13qv0Z++acWLr9ovJIGSIfbUakx6Vo2P2PmWnqsciFgW
ZOLa+GSfWfThyZrO5JA4+3VRZAw+afw9zM9YenGFsEP37wIhRLeNdTv8peV3xyYXolE9NgSo/iD4
QuWWxDePnxguwigzbKrzzZ67PPtF9yKf2cOgUo9sRRTm1zIB981Uawbti1sLmKyTiK5XyZSI3R71
sau0mAagWovGtUxNkTS7XuLEdcBQpzStsTlfEc3w7qoYzbbWIg20nlE/xLzcUmKNv/MoBplj0yCk
6TE4hX16rVrSGXTUMsN7t8dcEMcRoRpFXNCVYv4yWBsYTB1kR6zxcFqBC+dAJ18LzznUmb1qCjl0
6R0pZ8RMdLbJ6uyo2Oj6676x9UjuinaQNmiGDP1kHY75b0sfoN1x9pb4N+4mqM0XaAc4QHKeQCvD
2iUCBOaOYN2CJIYPMsmLFF7Gl33SWa+8at4TIvuiUiXMPONDck1WsjMyM3ECwzWp2FJKb8WUDrr2
cQJt7ToVdYQzhOQ/T3H5JljqWwuLsnTM8vLy4SBpaVlMVA0LiVZFgsxOK83VAGv1bgUouB1tXpvK
5ALDR54+gSG8QVMLKQ0/i/JhzRixbgEnLazXlayfDh6Ts6S8RuEDc80tBFPVQrOUgXevpS+Y25uX
TdN6wXJk+biYav7G+wm28oqf0Rd10HVen0kH0J2/JI17qWflHJeHDhARp9BaT7LmDWYEm72i/Wru
FAx7+k4aAS6VXqr8dXjrJ7ppkn/Gy5hcfFIDh95XxBraEwyUlDkpzJP1u85WYvPLThnFN1A4Kpsw
k8FtgCiR2xhd6V6x6Zqhi8VKDfvr0Tn54SMryPqpk+EGoC05C3U4OwCJc2evFHC/GYXEhxk8dtq5
bGnTQRFXLVrfP+WaAVOxE+Y+EXDiN86g/ZQnBWLkLW4G0uZb3nYMZwLVQcuwCogi66kc7bMoi0Sd
osNDb+TLuPK1IJ5qHNKvuEOEGabNEh5aQh7D9qXgUOhxe/I5//IMdDywEA/Gu7zeeFtzXFtL8EYm
8aduDtFYuibwNAkRhS8eGiuQZg4KEhBAF7bmWZbPvlzWWIXrIh7K/AN/wIG1WcJEFBn+7kDp8PsF
cDHjKDiK3SQVMK1rK/futo+k6L+xYGV+SLlp5uL0T0Juga0mmyYCcMxrhkl02pkXw3ysZcbuM96Q
Kn+AVVU88wqtidbSy3RTQLtltCTlw1QtJb6S7nUmGWXcWbjGzWzNSrSsCt2c1p1ilmNxuJAt6Glp
CrqSWwPIUMihpwOUid4eI6SRxG9yLZYokVkimwnHtM1XYnl6djUCAKcru2b3C3PxeZNCOjNs/kjA
HDgh62W6IGUli8Y4YqFLnVPN8iXRcfvUQxmMLYEP8puipfNmZBggAXqaoDHM2Fru5sA69QLdQSW3
HEoven86WCdmmJcTeCFaBgszjPbxEKacCq4vlIllNwzxtaf9ci7dTyNFrXfrEkqymQnjcqlAKKRk
jxEXOelxMelVGhinMFGvhcAVwttt+AVwau1+DkYJYKD/JuEdUvQuHmkCXbU3rtBVyuojkcVtOxN6
V1gIydfoQObqC4GWNWeIeUHkTgktPFgouH3PrToA4QVtiZn7q8e2/jcDA1nrhQscdO6YvBTYUm6l
B/YzGlR+Y+vAPnluL30l1oAb0fqwF3wrRgzQ59X0dOAdL4vePLjMqT9KbEn7A3e5DVpAmnN8Fjzf
l5Rjnogjv5DzhAGkAD2EMgprI27cWh7rZRTB1tvP/VBuMTW674PH64HXfchSGyhDcRlRg/vFuuAn
q19MN1WqqhwK5TF3Oz5LaaQAEolBW4I8ptt9gVevM6RuJTbCBkrF3qBt8Z8l6pS6y7eyk5pHMOoH
/HjCLL7oHacG67SJVJHhI6abT/uFQVQ/cf7atF3tyg8WZOlEszpST898USq/ippNhw3i95K2IPBV
TP2pS/RQ2/y+3dEncT4kWuMpaHDDJJA0HoxtjW3y2XVngJWjsY2biLmYVCJUD292ggO4HoIeh8Xd
7/wxAurp0rVYdcG+kJrFO0cvbbwjMWXFKb3fCJZ/3/WXUf+cnoBbzXdfk6IHT9MAMbSlM550dmCF
nLsc6wmSfqXAlN6moWI2tJZ710JEJok0+bcUazfTJPt5N95R9b26ABGLCZnv3cPcwxunhdHq2huZ
SGDDf7bTQw4DsqX3p2zks4VR6TD4j8UORtCDZjC82xBD3kWuCaVB7Kd6hI5am4yzLVEYKmFcxgw7
tAxQPHJ6h4XgtWg/NM1LJmFtemwRtpwt3covpxKsGcEkYZ146PWl3BfRlviasoebu2taXeDSQuU9
A4t/QkEgOkWVunQz0mwb5Nx+ln/SgJIj1GiGh65lc55meX7R5Vy6oGTZ9oVONzL8VTOtPDSwDXGh
nV/jSYyhYW35GUdS7fjeD5EbTSUFtfqsbu5D+Y+KZCtZuxA7CFCAlgOSLisTvVM9YXeNv6g5LRrT
Fii3V1k42ldJifZRAtgKzpvxh63kc7jeMSWNRBruryaKhjY1cp8zVJdWK/GZ/O2ejKhFQAA//5Gc
/dqxoq6qKSMzrPLtBFCCqY4SVluYVhjp4xSWSZ8+jkjlkhxGqOMC9JoRqE+K7vVL4KmIDctmtaxk
v4rvfdol9u5HMA1vXBfBBzuSDAxH2x3KWuMn3YOTifOhq2MzDJxwLM/wXuM2wDQ7aqIF8JR2aITs
osK8JprLnjk9pzYarx4CPLcB8d0SoKDx47oX2QYogLnR3daRR7ZDwGI24P0Ug4GMNu9GLuUSh5mG
ShsvNqoT0wrMNtREcxBRAhaSctlggszbxAJJn/mb2jyy+SxWscOLF3gijfKn0kdx4O8e3DkJDxcF
aBqqct6ZMN3MM+P5Cr53v1TGAiBqQljZChcbLQDMPYG4a31Wm0Q0IrmzouP782vxYwPwsfrWFy1V
hmJRIk5SPlweqD76iONQ8nxFaHicAxV7DSBaNBdMweYgyx2kKA9DEkBYCaO/SALtzKLGVBzt5+WP
TAI1M2Y5NRGDjE/1dLfux5RFDIcP2Pgy/cV5G4HjBVywLxSNR2zQS1QI4eRzga8Jg2UutyyjMK5N
rokOniPTQyaXNg9fFKjOesEp0PVvHUvNCkmkbuBRG1z5KrN8DSsa6jVKXp5cnGfNTEUg3NrEdWK1
OKadxY/HTKB0aNfW1cy5Wxn8pGQ6mJSVnTq+xOR3Pt6BVfvkmCSonCjOclpmzYur287doTnuF9/o
Va8aiGShmZm6JrCoGLMA3cAWHmGLhFiSdt5PdmriOkOGbhuVeG7KDNDp6sqfLlhAAIpX331JEyOm
n0THyM5YwVq5prj+vpPCC/3f0I4lUcgxzUXpVkVoE0rrdzR4xzKt6qTRTtO4RjfGSieMC8ptQHmr
WA+zHQpX4qaOUkvQCEq1zwDBmgi0YynmJwX+8S0mLF8IZbKyzET+Pj1QZ9KKEJWdzl0oHbLdGX6r
sJAyMVlrJuCxlkXzX1j3ZBMh2XqS+OVuuP8tRxDGFGfXkYYNOaFPj1g7kR41sX7Q7q2NTZ70XqyT
xyUkdzzrEwpM4mUxDXE4+cI5TAlhrSo5IM3P6pqkI3L6daVRY77yIguX41q9gHu6jE5GzokxcMkj
pgNmsVf6bPBzAgtr5G9sdwsLEOalPtJRwyO2ryMT1kEAxMFHMzgq/MPqBtEd6sRixqKzdHK7uMcv
vTwNjnZYxISKqdSp7LZRyVv7s6F/X74nXPGIswo7EhenuZxbc/OgBhYosSHMLH41vr05KuSxc7c/
XPYEpnP/k8woupyaijrFHGYrOjI0KcawGXCq1IzUwSQbkOgpz5h5G73RVUhZXdYITnXMqhLNZF1Z
1fqqFV5mwbXwUSAmAxtr6nL8k7Tjw8KWv6ePg7qpVimhCnvq9EwJewgG4ZsfdZMUUCoFLmv+jAhN
e/SLsEXS95xTn4JwbpLX5jnk7Ihov/prkOHWqJj+V9BJS7zhEN+IskU9wNwufAF2f14FU90edZoz
ES6bDd9kQ4hQmZN9Bzd/2rdRz5Kliqik4JX/GT6837cyFSBy+wuG3ZBaUI6ZBwXwM+zIzjhZ8onL
w2W2LRyn6r75uyOubukTtwgrd9/r1pxUqiWDQN5BQxlz6HMrH6qKQgKogUZRowUN2wFQjx4PjLA/
H5M4S+P3edItGdDTzTNj9gzjw4xoPxCfYClkV/42DRJ16q5huAvD1z4XWO48uvMxnkR7gb49tkAW
UbwGSnX4mvWpm02pgU2nj4NZ/mWavALTwEhT3Wod8Cgs+AvOrnLCs1Ham40NJMqjeWLZ1YnhkM/d
PW4cI/p6A6C1VLetNJf2Wuuej4DAnf/qIwsrwPmNLA2cF1fJ0WR2vLTHntFPb1K7fQWC/fwrpRGh
ciRw6Ur7AI3AIckKVUNzBUibqI9vGUhPqvFb3GosAFZjIfdM6WuaQKY/dQF+GgrfqojbwQuZQ5FP
cIZZa35A5WJyye6KHdkC1kBLcSYdDbaOwRVRw+r1f+eylF2f0IFMvgi4+jRF/G2pdxy94pk85AFg
EWMaKW7FYOBzd680XT9L2NOP64Ru2K83sWeEKaII3eck/SkIwXytPfBV6CTcqmCMAyfDElIOpP84
YJ32i3kvajzOw5nIZfURNfphX2bwcRPXMfa5jH8miQCyqvGZCAvDPeIb7K5ve77obQDkiI6QvUzj
lyXEcerTWSPpjY3I6rdVXHn6WSSPwVf3ViKg3jo6V7mUaL1fgGixehzJyXepKgvIrIk5l8pmcmlO
t+gime7JmCvrFJK4Lew0Wd4VSIDyMgJ6dwRPmzKQ16EB3iVaXktSJhYwCpgTPwAwPUgS5MClP49c
Ue0IPjQ+OlAF6M1w+nKtDc3ixPq2VDTYpFaxOIYwtwXVJ28GoYBW82rsiLnKCK6YjzZSaYcF+gnK
SADRyfgivu1wyjGKEW4s+9hcBf38HjRo4KLnZ7FEq/A/BRFlWc5+vYVWgI9V2knaK+cHqnbnnodp
f/zQOcgC9eEoR4ik/GZWWHWIiPmwqdYVjV3S65XGix+FAhbgntLYg+w2J/8+wkhNySsjgDLpJQeb
hcwzKZP5H0bmljJ65M9oO8+zPFhs9T9o7KM0MOAq47Qn2aV600L64z5/AJg6dLrvtMdkxKeA/p5V
yPqi+zutOuqb0Ao1uvGOycTd5aw97bc0FzMgeZjoH2z9cGcliWiHcv9b2HDcqKFAtdVW90dTGW//
fP3XAOhI/q2CKX4mwWBCELlU1IJ83qkM10tRslscrPfiU33ZP+OszPI3F1KXB+T5yy3tlFsnZ7T6
53jbB/kdxyyvxJrblg4+waAWHl9WxdGfuiabsNgc+KDmFnq38O5k7ID58ojo2gMUMc2O1+ECM/FF
T/GIP5mXwQh7SKciK6LWQ8tVeqw5MoQDsTLXMcPatfPcAcaR9lPwsP6oKLD3pd4LMTqwMzvkOzn3
eRUSCH5biTbc+GQqMIPMRz4WfAuB74olRRC4omJ1PtjpnetyTVDW8BNjhSrllXIjYe5xL15L4Dis
UJzG9JiuNT77sNwt8mv7ESGAZAUKqEIQujlukiXq6jKbvZoC+GmYfeX8k12SxjGKnuRgrvwIxx2C
P9byb15dwi335tfSG6Hu/rhvrBgo1QfY/6nDu3Ehw1zxR5F7TClpGm+IqCa6EUpyM3WWCrvXcsZZ
4iu76xlipwG3dGprd12Ee5azWCnbnTB7UvWMv2FvDbBPPRTromL4ibWAxUNKmzUlWRIJNaTJpsj7
gbARVnVX68W1TJYQgw5X+AbDpROCWw0cf1AzWfAGZzZcibVSzxRs8xYVHlyhWE5YZfQjNJmaCDhh
F9Ma7vtGiZpiSgshmZwxzkY38ZN7NNzK+l0gB7Ae9uyT3Maiab8nGHLxKALiMEX2axarWzfoNJlL
MQJsCL7k0Ky4uQyM+T6dSTvz4Vb6utaXTHZqLHGM4DHH0Ezb7DMRXaKVoSBJSvkDV7TUKDrXrBvW
5shLgDFqDsV9bTR1TdVQHARVjsJuDB8IkTCNgssq2EFoMIrCfqRIgaebAaW+Hh47Pmf5n5G+knSk
klWmvnqFUAyrRwo80Xx2cK/rOCus1CEsRfIghb9Nu0Ms1KTAuRnZsP0vqSfnO2jsd4+UrSx9E5tT
uR4A7JcGC/nZGNd0YZHpzM5ufjlVpKwXkSs4VTMZ/V1p0MP8AEUofncjK7TY/vIj3XDt7klOxU7c
12hXFndFSVvZAx72tjXEp/GI/CYVZtPkb9AgCVvcPrv7pUGYfSNSkUgKCLte6WXF6c5fhHhTaUOs
250eAo8Dy6rQYypPu2UMHzS4HaIwAxXPBmjHYPkOiiuk9ONWRIEJQYgCcnY3ez719STtPLcAzyPa
wgnCzoQXFL6KI2O0mqv+Ye2YDHFTnmRWs8Hr9PmShmJv6W2ok4JNQ9v9rRGOAAzyIosapCsREWg7
B8SNp2p5YtiK62GhtXqM14uE/HvsLXchH2SxovnPd1j2wr18CjY8b4Qb+bsXKtU4m4CylYvCz2LR
wVCD/i96RmehWdsjWGPCr+l08KYyeIBfdYb84A23kvii8fLf1cBZHUNsNaVAMtPEl+pePhAcRm28
X2YKkqcERvIrDYRKSSnPlhJ+WkvqZDCXKNVrx+1QeTIoMl7sS301BpYafpO6EpABxrWV26BzDwlf
GyKFFZQv+gdK7yPHWkTFKwH79XrSp4Hr1aOs50jfZLtcK36/8pCcC6cI87LL7o2mV7N9KVMcDuiL
mbultg3PZyfp2oadZeoOO1Pu4g9X3GrB832bANckQVLfWT2ZJG1Cx76OVZ7ey4sI7qvwHYh2diuk
2ZWiLwZwgvg0lkw0C8jKuZRZDN1xZpRBm1kdhZyYdJUHxmkCklIAoiQ0RqzH+XL1axFabaSngsKY
R6RWRjxq6bw5TUTUry9NSI0Kv1WJSnNVSNW0AApG390iSuTSlB8wXIEmnn9Fhehnb4NbXiey9Nlg
vfXazXcWtibyx1iDI301I/HROhRPqynM0lUtqt9FkRJzArqvxaSgCUjOjjUnDbtfaLGNV7C8t3o+
28FlDmhH8Wzo7Epb4Jp9MtvSWhoBmFSfUmw9bhHshV1V8XMP/q3hG8Z5ZBwVxOJ7LhANB2HOanAt
s4ChZqXqWoWHPCDLulun2m4to0G5mBpryAAPvi9aqaQEvx6puO0w9K1VlmwV/yxBdeYj8H2odHNu
FoonbzcdsinTI4702ISNsBkz9FEmw2uaaK30+bHnMEEcYiUxkeJzDhO+cgfHKZS62A3pdqF63wt6
WD6ypmzZNwz8VOBSIgW/xZAagcDnipcs+ewaC55XyAbA6LsjCDPEK4wvjxleas2D0gvb7zv360aR
wi2o/BAVlFPvgFKX0gJyQyScyoB74BmYAcZ4vzb3Fds/k5IP/CrZYaWAWjZ+kW/GN9IA2wtx8U7P
IN4OisO+FjBUIKy4YK/+/DGFv5Ef8mAc+r5l8Wb0D7y9StdmL3agAMLCZJvELSL5mkwg7116W5r2
sTJUl6P7WrToMnNPoB4lzeD6tg964gGHAoKUtSR/v0bKJVquqjuahW6m45vsOyP7oHJPd4P7PFjO
iK3ij+K9GLKoLxyXQqJ+M1JKOy7PARGta6igQMjDwj11Pq1GpvQ7gOoS3XJNqu63BcYWEmQ8Y9Fq
6MKPP5BPKF+oUQijHr5x0LydLpBu0yhc3W4nZ152sMf/1M/oVB60NqLIMmePP6UKIrFm8TrdwKMD
Kqg/6ZGV0Aj4GVzxrBM6ptQgOCgYgkxJKmgZLg/qWgW9GL7jBVflqSKKxrPDaLYC7ocSUmxiTSMT
JNWTT3FVB+w//mae0jM/75Y5R+V6SSAO7BStQw7g0+RbTVEYFOjnZFLuFkxswRb/BFX7sVcJ53i9
8KS0HCm1S9WsLwdUhuzghAspMAEUZvI3YUFqH/8KmBC/1kyn2uaCZd012WUy19K3h+46Y6xfuYTE
i2t4T4KWdcvVQczSzsTcPmxfi5qgsDTMO4AopaYmI8+5UZ12X+uQI0FjVuW46lBbXqf8NnnIiRE8
N8ZMAguBRkPtFFmJ8CpXnufK/SBuVzkahJJVX1l4OJ8wMTr0zFDG223OVCVNoKK5qqFfoeP+u6T7
/8iC+KIGNHmTZZev89DkgFGSG+nP/ZP0gr5lHND+HFNQyaE22LR/noW0nBYViGFplj/jzD1oSTIL
TTjmcwrza8s1nDEv7LY05dcjtRAMBtpALEKrdYfP25Dq76F6kzTcXcR7LJhixOXNmY22KLuElTmD
AHdVAEkF36meIfzLiHcJnpBtmKKePDea86bJyV0r4Ir4qQBlVjxpyOOCqUYfhR/TnplC9qrictey
art645dDLAEobrjiZFKAzHi23dcCjVG9KwEuvWG9DjTQmQGnLwPV/F9sYbFlrZZorKKoHJXnU5HE
xqkQAzJ/brmGimZKLVvXDeDYZ+aLZL39s4xbkBOUAJLWxHU4oQgmBk2ADbYOAYGD28X/9Tc0I/SI
MJhOQEPaety8U52NefahflI7RHEaA9IjQaxUn7aX4IBJ4CXBkFxZakqlt4hb3vU7xLlncM8gGjJh
iamFoIgcUdM9WbnMtUTQ6FfjXMxCM0FsrBDen9sKeD2CZeBIeskrKO189IvbGBG+XTwm2YUthYuR
c6pwm0pXHwL7+1gZ4FKRIlpw1OLfqpAiLvdH1aj+2w+yR+Sa7RNauEwja/QiB7Ut++9PKQZwG9oP
P6he6ftIzyGnVnzVYr2DXE7d36ddXogzD1fWXo/FnQ3XN309K82j8/gL/Upk1w/xAMu6EiaDb5nT
dy5tx+h3W7N+/SmIRiyqsDAOLSDj1B3dQfKxmVIuYcW6x/OAyh2pIeW1QS2l7vbkZT37Ef86k4QH
3hYqRExG+cU8KIl1IXycRnzksj2BLIod8HHcs+DYhrem/bJqzqW64BdDS+DooZA6DpVru5kg/i9t
np5xsmmYEWo1raHZowJFd3vVqqc92dt8QHskE8PIPSkuts7RNTcCgiYc3g2jFGmurVCmQL22Rjgy
4Jh0BdeoTpa8PRv7PjnKhP6nm7FAJ9ht+zE4oaw3X4OVBMtaWDQ7kM7Z6Cif3dfbsQHhgArNmVeb
Rr5PrBHiZA0egTZPqZlUcEvELYEv+vLzd18LhHxIeMzMdWEjp/xKlmqy3/NOjz8QyXB1dCNylata
gb1Di/O4ViTLdS01aow37oJUK1aq3d7cGiRdT6LyCgplF6/iRaIhiXAd5GLzmX0eNHnoOn1N0+wv
kFifgfU/JKE+EYm8Jj2HxO0o5rkYxFNiL1kZ8l4EYHBN/gaMVpipbcjXcgQyE2ClIppS9XQ+Mzjq
4reZ9oMyfqXyZvZAPEiGqB8bcg5MhDKNs6mg5ee5vCSvB+rNACKXMHn59GcjmOyX0jggyM4x42Gh
6AEU3+ZwqVi1DMUYxQlEyer+TtNrVapvMB7HZ/kIZXMd9gCKyflEySynoD2fqDW3Naio5aXl+aR7
64QH+q3fwHqrhNGcXDh6g4TVOEScfKNjQFzjH4ebwSah7sQ/4wzO4bDTMHu7e8xpkXxBmCJkr6ZE
MYU+402mEWresNa14vG2Pu7wFOEPOu5eUW2O+HPTyWpywMz0HNKVk8wT+tHi3UYmISNf6lYtOP7e
mHwphkXL+kFMkZVoTm+ReAqAg0HADf8EV/m4mLYpo4WaNhhKjXaJwgoWQtbhr91smHCx+LDBvIu1
12J17t6RfdOU/scEYTcIlqgoD/8+YWDs17VOXzrDXZTb7uj8BUEloTELv6oxaSRy/DVs1EbGE0tK
suebAwvivMBH+Vv19cpDGhulelz16xg/IxwmbNzhOkONfGXZ7UzGzu5mzaE5oKTZMgEN9YCSsZuw
VZObH6pxg5PNvTXfF3K+JwncCBleu10YkxiC4OZxxVM+W9cXWZeotTXBQgmBpz19wPsQYN6YYLNt
ixNZlriZHctIM7bg9dA4H8XT1GRXyczKZaDqdoxx77wZ74YJ4yYamXdJpL/VWU4tPpzjwLw9l4m7
ny/ZuCKTYsoS4RUdlTdEGdacl4PQ2fibLLHtIWefZzHjfE5hfeJBJgeJKyspfDS90zDWqhrq4LhW
8yR9JPyZnzmGvZi7pM/om2wW5xW/y1wKU2TRvAbUUQIo0AweHVUtTgpbYkR5dlO/Dg3Ig31FPBQ9
WOEpJ9j/NT2BfBenbE8bYl99TVYqy87bGRCD3r9RvD+JUAJTU4WQFjHY/LIBYgN2GBMXJkK5Flga
gHG/QTo7mq2Bxvjch/c8Ncndo8tr9ibvtifUN3/ZftBxPn7rKJWuhNDWIiAFqtlz4tFMlXDqes97
nVj6j++oU00gWqiitmsAg4IAKDToJMrWjjyxHM1wwkkC9QBQf6CCci3xArGM45UJTew8tBQixPMQ
ibOLnRCO2umkOsh9n1UGNU8ga7mdld0zLiS9Hs/lHuVMo6ge8qjq8zZXnfH+bM1ZHZGJKt87ub2q
df905PF0tZKo4FXXN91w2yjRR4HseZj0trgYdrOv03JMKY7KeTriynHPd1tyu6fN2OhgUPAL4+tW
7V9W8vItlgQzrLl8/Adw4rAS5ETjxPX2ac8vvkPM+sakvu3Bb19ugAKkcDOw4H6vfVRYgEFtqpGA
HpMPdVflMBVhI37SvDzJ6jZX8Rv8+gEKLzX/fI3sANa0xYNyhx1vCl5lSI22cwlgAD0CqNqKyUGj
b7DCi3Yj6v66k37C+yDhaBBaJdGV8jELT0cXd68cltJNdc2yC5kX9NglLAhqmx0OBE2B4qe/vxf9
IeckwGMQAaE46+CPsk5AUNlW5W3WskXSw4yH2MbeCGgHCmhX3IXp8fgKHd1sDoTuv79Q+sSumKgV
cKpKNzI+ODTOlpPiOTQPHyekbDRqNwCrcOf+icikh2GlTj87spQNvlcA4mjwfIoE+SxDerOVIOM0
6WnQMeViPmq2ABH+XlXjRFD0Ny7YKMAutpZbbyJwjwaKmsq3mcMI13fra5ArCegYBJlpnX9O82+C
JcaZCWCPhArY9os7Y0yLEFWNVgAmQiV/IMSiUBImLCtXi8WJw6+Fb1QHrlPzQZQPDbYqfYAYWfhf
iiu/qdlGW8/mUOvOZ992/61aV3PYxkfJl6l3YVsvIaEM6RBu26gCcNyuhhZT92dVyrLWn8HNaiDb
MEwpuVkN1FkWknxOf4NsNyj9aR6K6L1PtrnX5Tpf6clN/EwYeda+0CncCeH4P6s0WQDVk/VGJDt9
Tp979cyW00yV+9Hy4AQk98Qum5uXJ+RfeyLvu/qW4hds9DprhjJ+3t0zX8dzItlO8X6+/OgPodLL
aTo5SH7Lr45/eW+4dP70erUyIYbT/Tgkg47TS6eY9gnQsLaVLr72mTF+r/xEgPgyXSZmI60P9bTU
IsYiAbpsTotqHnXJPSsir7B4/PxPQo3BShnyTZUrwc0ucmUvxjU+qIJ0/Fx2ilOWhSlDRY6xsv+0
SdaVbNfhG9OI48JCe9WS6RRuKPsQtfMIy5gu6LAkV0gWUYHZpPDMJcMD9jOLN+NL+b8xcz6+SlB+
+pW0Otal76X34ru+y6kAwHFyRNOWNWFZ5Li4il+JfU/AieH4JfBQ3tkbKzjVOdysiC0BFM2cOg+y
i6bhii8eIongj09uaarjg5M1tJA1TLtLeMwRcI+cCd/2m3zAgHHN7gNaCmwJ9BSl1FLcNjdOPk8s
GoUpmmfs8xJ8VMcDIMcD1EPIOBplwXw3wC1FD5Vrhn1hF6hMqdo7iXAweq4MpfFblvKL4Q55674w
uA8qCoxEwF4DFdZQRw2AE6coBYV8Qiz0aK6yQusjt5Va72fshmvjOfx4R0rZE6hnbk7qck/v5+hQ
q5sjynmgzYGlbND8A9W9HR8COvnB62lAhv9D2KGrRsd+HlzmhAKgY6hrFW9Ou7oSP/2DDLSldvj4
BcD1SGcswv3KqvgYpmm7hr4rzvaQZ2BdYumT4KkTawizhepdeIYr65Ghrdo97Qwq5diYu5oDiXsb
mhDA9IHcCegSNgRLX9WUePo77jtDrV1h1cA8YNeK/Ap70BWoW7OIUj16Rm/coa2VLiD3vDcIUEL1
C2NWB16+8Kalu7F44+ewGJ51S0/CcMQmmqsitPncWR7TcHXl0a2NU2Zs+YAEjYd5MzaIR0+1KWWt
nUHt51bMAShVV+vwCUtyVM0DYbl8fH5CYx+AwOUQ1lpbNTGZ9NNuQBROiy5UXGKrRkIRk1r/thmu
7RrAzcfFOu4vRhloiWHxo5MVJ6ouKlufdKR1Vd6en0xCm6auRPmuzb42tbMVN+T6YJ7uEGGjZGKD
VI46SleO8XJK5NOSY3dPa42qhbPRtjyThUwICsGy6FXb8alCzimMnMup02SBpwgP92Gl6sEk11iv
msgc0xIkc/OapyF1p9/gJDzjIXdBhUh42uR1xYGD7wqq2wKI8UjXE5FD1WAD/fpKu/RlK9SHA+fH
lNR5DbLPQNdzfNNL92oADKEw3h4CvCm2DEvLGmQpBzCfS3WMg9PdwVa9wsXpWAVss6NMFLlpJWkb
P/ULhJzOvSt167HHh/bTyteSrQg5GBoum0GJ37LVbaq5IT+T4oMK78CbJ6QiZO+/T5rFtYyCf1vc
s60O8R3FaeH2xqdXHsphn0q//+BYHRPv3kJJehgWs0vBXME+PjR2onEAna5OKBKWTqLtEbqK/agl
JsJ/94TCqOmsjDDDgiMA/HZ/4708uDHMvlflx7DWbf36J3xtyRA+1APpI/dU6k9/OaCtQk9JXvmz
Mqax96dnD8JhEPTX2z/hpg8Rzcv4fJE3t9ZhbpQtl9MXyHq8JTXqx6xSZ6wpsY9LWRlW+9tAwlta
UTsa9wdzphVCwdV8+ceR6gxelIDQZRGduCcCwyaPbB+1u1EUTYOYUDIo9ubFHz9OqtvzhPIwQ1IX
DZqTXPvNATgCFgYoq3uxLvPFkYt5v7BRIlAK90Sn7HvUTAkzcSM9t7dbfXtbguLnXBAvACbc0+l5
zz6zv53tdGDcgnXvh5R12Qdu4Qz+LJVe5YGeWXYkS4KDYnt6plwU0V5yQCrnNtRvliDdfE8tb0ys
ui7x+Vj9x0MsKeJzR3mnY+FDMzHPXq7yHinzmphl78ThbUyT2ZUmtVHI+ER0yEnKpGWjtf4L7edr
XzK33RpdWhlREc6k3XhmWedZJjXleuphVYSKhVRqOXAyoi6Zjk64KxGWKnDL+xdQOVGEet3TwJXH
SYosOd45iIW6zmE158eN0BdoRRUTzvTgYnCW2LOGWEYVGKadEDKW20XZgYrtXxxAXKeMUu0Suxiv
UJVwDQsVo0UPCLgwr1jDC86J3wmaSZjaCT/wY/t/XV4Q+CIfAUZAxKchOQ5eyzHKdXJpLd6JyGCP
RyMeOiZwCUGuOUQpnnWvjwtW14ovNJw8N3GXzYlw1YjSydViv/LTTIhHrJsTH79HeoHkYPyrdFNX
aO0UZ0zuBTsXPS3Al0TNrmWcLCv3uk/gGQT32TC1qhEjeSo/KLKO4wTibymlpXxKrL0MbHqfYiHw
mBdalNTpR/yzxeOOXuG2M7VMKEZ55w97k/zT6scBxpWJya5E4lp3F8HFL3DmI+02E2W2tvnKZhPr
fqX/8vw08xQ7qY4ZNG6KAUk3REaBjyKVfo2rNDFkz45wnLsBiF/oiK4i00gWBZ9icfO7t/fPsl7E
zdTvFf4nwztLS74hFTejFWH9zgOk8dy6Sq47mXXerf/C0hi5ZZNAES9707V+EN5WytkiByLqeT0o
eV6YjUY1VRoDpi6MjZ6jJNiHxmW4Bd17FNRaRN36qxFQVe1BGU5vXrr27rHCkpSMfJuEGx97n+JF
sS7dXXsqzlDthWB6ieaKZ8F4D7IOMOTot8KyW97m76BspkTNHhgj/N6qRdceUywDU0KZVn74+hVc
hW6OVI3rvIbXeN/AoS/D1TlusVS1yxrn9irB+G6JRL4LO11hy1MDGc/jma9HOg+GnnLavpSCDFNC
sys/9g5zkWV/RXWbnNEXz6Ity6ODXEdFmjhT1BCqRVP02/q1B9TJrz9t2+GwcTuQ+X44dWXKg7Ri
jsAPyXpCi+5hm/ohV6G/gdyRu2zTTvnHkKBAdn1+NieheMShTREEnDFjeI6zza4RiLbznEZ1Zbn1
p3FBxKjueTS5Urf7bP31SEPlTc6NxzkIqgx1WpkFiMZvzIQsAVzprHtOcxddim5cGWF3CNGZ4c0U
sPCIoyKeLq3RALY1Yp6J+Rb6RDnTRwD1X7XsSemVV6/BD9nqkN1DOgD1THkC5ITxxhyOVYgdlrZ3
qGsG5tKlrUfoAbXlSiW2LVyLY5bIaegDa/cpoehv8i0bQgsaRNw5QE12KaxcJrHu46esZ3MoFgTL
WoKeBd7EUfSQtwBlQjTz/R0t8qJt/soZMHIV3X03eH7lFcr0Ubu4dnC674gnZ2TibgrrT/kGA4Qe
EA/0kUmN+5LXKpUiIpy3hynKYYAe7sXj8324kNE1xnfo7CcJWwjxl67jczJ52nOfHGysmA2Xfwq1
aiVYXwRGgAnr1G4E7JBFUyvZ8+FXuRCwaJB7k+NeHW3vMR1EhaTVCxxwAtDOLzaNjeJoQDm71nXh
wqaikqACFysaqVzGtbmJjm5hmVPMfOfYih34A5yohl75r3eTMQ9zfr1EouxcAkyftE4XtvvqbI4k
Bt+axy6W+b+j3RALfWAayPiJ0AgmSpcvJk8ZjpHirOnNG7SYCvIYbU180bYJEnb2gF7v09Gcpf0P
roINKzvg29j6zzFDsiI6VCg9yxvAg+yZLfLdGWh2fQdPH2MYLpnc6NuF+RVsCYTFu/PFP9OlEe40
uIiPA9lQb7cHsxXvfgmQKEi+W8lMZTGNQ02rbPIGNjKWBHSVilG+QJNc26uwjKCOEBYBdWiqa22z
p7e6UUK23EI091dWHfIV/9J3T3Jt3e2fLPXSQ9smJ1Ty9t7sMYTXIFcS8k1t9viFYpNNoWY8TsTd
PsqRn5dZhGgEy4ZprrMfnzXYG2aLSFplGgRwOW7JlJsFC6I2/inclPLNaOA25HgEsu0fV3wA6L01
SH9HwnUkSMr6qD7QZhOw3MLa5aVBpSaIsVPCvAExhYC2PqxZzxW+BuZw4jNNlInBE7P+LUQuomWa
pnmYNI35EBgFjAt3r72nhovSr8OeZflCoy0nA93L6SzRJyR2G8hS3B14baSUGUjsSyhdEsY6yEIN
KxjVe+wWFaT26G3skKu3XxAv+y7UhHd7npu+rVoGaUKrvhGfqQ2RujCpeS6TK3X+J74OzyT58BOs
mJHGrA1w5HiV9yPIEfj8c+QibzGuSSsvGqOuTmIxI0yoEHNdc7LVBZdv7YhIg9PnOvpgsiLcbkPs
iZkCOrEZVfzdFfzXkfMf8qGSSC9YCrTou0nqKSBZk/wQovjMvkV5cnQURdFK0QpLpJOIxaam99WX
9qHAYrms0Rpk32KXXaLfQ1VDyXObqChoASY/1HsvIMJFyVPRfI07di7nd1nco6CwQo3TB4h8GSQ4
S8yk/HmNtLdlKOOXRrlwmnzkfMSp7Lzf8+kbMVSFfsCFb3NVxHtnH+J0lt2lAd5bHRgXOgfqx7hM
XNJeuKEo7jxZ2qMjGlSTIgy+mI/6/0LXGMwqMxwNhoiY4B/WHvq5WB5fbt28a0cYimaagIO3Ud8p
QcN9qHrV7TSkdnEflxjvXAxFLW7wvNqQ/P6MI/mVw6+95lLPt93O4CAbJvFXjIOuIIColYcGg4eA
9XweM/ZMunnKOXUOgJ1ALePWnqt0a9806zB3t5ZFssdQTwHWntUvMInMN8pol+FJ26mOCZ7E/7Jk
SS9vN24G97W/qrZYdv69q4MRFLLKrrLendTxU5Hq/wcN/7ItmF42t12PQN+DSQdO1vQGREAF3Dkf
+1OkC5p2CZOjiFfJEnM3i6VKc81r9aILIKO2kHvvgOWD8EA4Zo4kCSirpJwCXvLBiRSBGdyNpGXv
jXaIpolKeOGz4biFK+NXtmFBQgduAl3X20fKdoORWcub5gP0LSVualWaBxvfVq1oS5ch9ju90aTs
sbeiTgKYDcJl+adz2R2qAFGP71FRghIFGoGwA9BVdlfq4kECHnzM/XPqKj+kiuBJGivhSkK7G41H
9z82m9HjXe9DmLNhnXbaRZhwTnM9aWqw3L930SIRcM8O1J3hvKcPUxAlgE3SMBxQXgecUnoI6oDf
clxxhcfvODuLzFX3ZRtXKhmmWkhMBf45XW9kA/NBw08ipwKGazChe/8F661Dr+2YCjOqq0li9/NH
c6qezO4WqDTODlegPbN0oQvexNLGdN8PxSALaYLk6oL5xwLFyUKrc9q6FagjXDjwv+D1j55exLVR
btgWptCbpAC4SaSSDXLZaoVlPdrODimV11OG8ewYj0K8jhSe7OXwLvP9kHcq3WnreiaML5I1wmcm
CHLepcCBLQaxjurRHDxN/Ujev7kuCA7AwtZ/KEXP9e+zQ2fRxxaxhJ1mX2Z8Q4t/rqOIQZFihjdE
7OlqqOXLg1+UquaVx7KoNhjSNA/NyeHXrMRK2l/a9w7hG0b/yVYI0jbtZpRWbd/fWS//ew1hQFyB
7ptNqSQxX2K4fl4tcYWIehjZVyppHjPw/zL5ttlnm+c0Jo4N9lhOGlo2qv8MPJVMW4175TECl/rW
yl/oe/MNYw328TJDrhxw9ZkRbvhIew/kxTF4A+2oJLQ/UyjuNq4joydNaPFWkk64dx8LaUDefGlj
h2gOu7ifxZ9+9KP3axrDb2jT02iGTIbUy+wphxrQFXUJCbhHCJS4yFLQ8a8lDAA+CuhTD748Jz+O
+NXQGVIjc7rksVzYNp9tI/XKZJ7mRRKXE08cf8ji4NLS7+rbMJt1BCWHUiigWPIyfqh73NwVPg0K
93aP4DutKz1RpKl5VRJa0mUHzf+I/gj1cEGbH4XMj2JZfoWn/InZzpG++G05El4Gkf7BkZALRb00
EfNg6TQ1gVNz++q8YTMujf2WmL2zgGA/Zu+a0wmrXQCHyMWszrtMVRQq0jkyk/eHB9StqCR8guF/
aWbI0oHqFjY0KGXc40ZXr6LNzRznB9xMBQ3DeUSgwTMdZhAPV6utHXyUoVQW1shieuE5LSo4Ns2A
O6kYrtUCo0TVU00+DU4+x3WZT8X1VJi8bwSVwP93IDvfD65mb/wOHQH8fRP6s5cNr2fM3ZzQdi3O
AxrU9Pf3fUrk4fGUv751CbfKByjXDeH3hPFUDa0pDTbHZ31dwv3PeOwtMZpHWiimXI6njIvN+wh9
kmzRNiwO6yOkQ+gyCYDBwCHXLrTW4pgXo5+SHsJMxDyRS8Wr5bsKOhzDcqvGf6PLsLQ+6KrzbJA2
gDypOuGu3c6uJlegmXlLKBRDKZ32lTLoxaRnxZzPvaiKr7Jzr23g+K9uRUOegcU3NK6SzSS/Hkvf
ylFrbh+8xAg2fNjphhR6yJHk9uIjaEP2WZRqV9DiK6XWUzAsYJ9GdmH9Bg1NdkLZKNRq+gWtGmhu
bWhH6cuPRYqiNcRkpaK+Po6ULwLRBoTtenxpdQv/BnN42GG9o0cg6S7CUYKUNoVXo0KKsMSdF0Uw
ppc8MgwhTwER3c+A9IIgxyIgagHNxH1wrgboAWXRFr/IPZyNXrUcCqSAGsuR+AxkdtEjSi8CsTGa
raUWrlnhGsuBqeS6grhHIDRns7kju6FawdOtB/s0BKlU9lLxwMFONlVUQMXXNLoypuwY3TKbX1kz
pcnT9ALGY3ZmgNZoz2+HrZPmR6q3TlObmYnFwLjiwdHLZmeefg9qA161yreUhlhfnQsujBMiyGfW
nnqzs4gdsb9v4+C4LHKondcbcUSw5j4+jnrI/5FHP98D0w4UfuOsGvr1aubyh9PaSfhUq+jc4WeA
YpqB22sVY2zyYcqSX68LVgxa8LKZBTIRQ2HNi7MG/Rp8MpwUdG+N8fR8DnNLq8iE3JBM1+bBHGyN
XlOVzq7mJddupb/UJebMYXY0hzQp+JF++3PpGUUZMmYO/K218CWqOBRC65pCwK85c93s6O2EgASr
FPCbxn6N0NmAsNcQgXjv8KSQbNpbz33m4+7ZlgScRuHpw497QK5J8H9m9Ix2b/4wcg4ULOmmSwqg
rz2THd0vh0VDySNL90qRCqruJWaQdLCciqzy5WrPF0flBqCg8uU2jDn7hQRunihT8EZJF3kzKLQC
aHmsDz+csC2kQPzecLVKm4S9VG5v37NikQOtAg92T2SCWDptiyQfhnfyvkE6yQyVNT6vJJWxBOgm
ylFXaqUNobwXSeI/sZM91fGHCJL459IVoUbpaKlhB7K+ksho8uN+aduvAUpbYzmNFgbk6P53kkuH
FYHKHQrDDOookEksgZcgUH3laearlp4z9uS2dnO2/lTJ9kIb1McvgEYh1yB1Qf+E1YcktLft+Qp8
0KeMPbXTnujvKy4TK2W4OMR10sy7CsFZ97vpg2XF7tcqvQdoIfbSw6QKpTZQdgaHHQFzYras8Mjv
T+k0i5Y7MtFGHLmLuEDGgaBShvkaYGEqUxQgTN4MEEtmE90T2xdpumTmO5Hr65rykYZDgJJIf3ue
nWKZhU9UoAtYzqFXGsvWvrkWAcYS13JYcQXJalC8Ers9DbENdBs7nqDd83jIL8TolEfPl3TcR6Mg
IpDBBqem936ROrk0N6OIeVCdATwL0PlENKpz6XyJAnmrBJHfb4bT4ctVEFn6dWB5r6FFDS8K5FYV
51Y89EdrIVCzotgUkaAX74+KgKbn/OWmIbf9SXgm9P7V5TSUrDC5TS6asaSCmY84eVJ6Mg8WGePi
WKRrDE9/IGdtm9+8CbuNAwD9DdDOUZqJdG9mHrhxmSOfoFoPzAM+cSyW8vca+G6JqZ7OLWs/uKl5
srFoBuEb7HB5QYYIP1Ey+I8T031811ICe0VHBBbGiVnlFnQOK5Z3I1hs9p8zM/UmShrzBofmlPQI
lGSZyOTTaAb7mE3iFiFJz57tifv6f9s3ah3y5UqjtFnmvNtZF+faQhbgdeb2qnK2j8LmqD3GUKA4
a5FoiZIHIN6rUkN+xYKvCFOCXreZuOfUibO6Y6bY0QncjlFVtewt4rQCtN0XZIJUP0yA75db6GHE
H6Cdx6vXvpirih2Sjsi61SF3wrCbwnJX3p0eVyD2r77X/Sc2157Gzf9wgRKhczDvdmPNsmmqNtVH
pPZ8agjxJcCqOqY16HGHH8xmHgwut/GobpAlH+GDyPpaNWxw6dhd8KcSEmyITwi3rq6RYSBkBNXJ
w3NyMpmjrrfS4Ez8vuTIuKHrk56uFqiXVdAfp0didbC1QTVZSxtyP30bkztBmH0j8ddZy8C7buKU
TNpCiBirtGUmZG3WTENUxksAzLLv1Jvq9rXG10Tu9WhK7g9JJ8ZNnfhGhwhd6Hi560OhNicmd83o
ehmTRspcvyAlj5vdVUc+NgttFlI+HxI+xdwHjT8oXxAeXe8XhBdaaR91WH8GKOhR0+7MFa9y5jiu
HORqiKMgk15e4O44/AZ3VdhZuHJYSc7Hfy35LwrqRpvenfuOFvHmjCF2aQC1p9OkZh6+FIdqxB9I
GrwGSb+jOxUgVeHIRyZx3TKcPKNAKBehv4DxBsrhVqgcAQSaHx2n+0XtBluFYoPd9/BkMnJWssVK
xe7+GOfyMo2pMHUDgkdgETyj5V216O7om44tRxCo3S7b9hPFtHbtXsaQ+OHyrQ0aOs5DGjmdgaG1
TvmdIETyG6g0O9f5pjuBGouF++tsiDThL+YvpnFOwWZuTrCeP+gEAQAobjB5mxjS6+zdHwcyhBWU
QRmkJNXt2E+uEGI3X1Has19+JCe5FvqsyfKLI48n0orLRlLf+BRqj3Gm9uF5amsfoynChSlI771S
q2OHzyCTLLopcLTgqHZGGnlLJEO5/lumNQ/PfRC1IN2kd/I0iwh2Bp5FwYKI1LQw2acD+hrepdK5
/HeJKACFvZCPbu6R+irwOOw3j7VBnrfwXwKk4yPRUlyKmq+L2wlFI6BCgCA/VcN8MCt6zlTSr2xD
NLeo1/QV+ALfD151pWDQxBJ2qpdugXirrG+IS+JNqKAsFTns3mmWk5juKq40NvrvE+F73mTmKffl
B4hgusmY4T86QCUVEjRuIj3avrRWmfuu91Tv6dDWXNmhULw574ey5SnzwcntXsIfaZqIBrjz+F77
nGo+ehSNiuN8hKlVIq5rYtijsNGP2kled1xBNNvgAuXvhzkJFlwm0NdYKrJSKqKZlnLzEwOckaEW
9xFF/2tG7tpbXHizRrE7whPtNcPyzOujmOj47lIjbn34Has3FE/lfhUD/pXcxgMLU0J5rykLsgE+
jmf/NHpyja+HC7h66uqdGo0uA4e7ZFZqHxI5PYKvkIoouAR/4rF6IP+EpQ19qVY6lWskrRWQI0Ic
6LYfZTu+MsfkpSc62G3KF2f438CeWipv4JwgtUpquFn2fKUHpAdP4xAqoBsm9vjg1lorss7678RN
Cq2+dXTn0KrC1+oWMqU/VqHXorPRxFbDCo8//MB85HLC06Lr9bzWNu4w1rhzvNDDCONoki5jdupv
3vmXl2HFU2jOaJHN9t6sFAjAK8hx+2qKTPWsde0rSO+Xsw2racXrkU+RBSa1hwzZGZXqg+XFXJnn
92p7W7rrujJJBcAriXBiXlDGj4eUOOP4SoFTYXNIJH/VnYYOwjcOfAFQxavx96zTSTJs5syRm0iU
YqIuf2XMmiSCTtpwrsxPAutHUxozU5xc16iIz/6eSbuiRjKpEG/udAZ3ANo50Ip70idirzKj1XeZ
0jdn/EigbL2YVzEtFC8tTEz33W6hW5LKK7/7wH+OFOAfe+h/shFiZnAfE3HaSlKMdqZtbKRUcmSI
XeWy07MtPbG1X1TPlHbNl3PQgwSyF/3aJHuAqbsnP99j9uk8+H77r1whsBfuzufQenJddMbabW2m
bGxc2GYqkLPRvX5pSJVLoCehfubjEVR9Ynmzht4MxV0xFBoSwZprLg5EmM7FH6LLaaG1LueGH1ZW
v9oeGCmsCsIcfKTikltCDM+C/3gXsQK9uznJsNcULrwvsxjec2MEBu+kVAw3Yaocco7Ma79NtLXu
WVqqFnlhB6W0q0nOHJmy6C6gh393A6dGyqxB5b5gNhIaE0qEBdWtVd4Q+HEAGDz7vHbvQ40H/LJV
7CWdAiklkwcocWk5wwvqnG1lHIc5IX5vsUqlcUvZwou9thWaEq/vYc0jrgCaCQRXxWalFEG0wJRW
1U2cMSXO3V3Yf2K/KToEKmV6EhDGfWqrptSqOOlVJ4DMqkkg8Z0ldL3XU2eaIck/yH3T+1CyWZau
RDmj0VJsH1cZyt8zzOm6xGLqyXIizeHH4RhBxOlwBVmwaMIb8X54LXWnf4bUw553tr8trFodE+Rk
K2psHZGh0Bxen5ydyEn/8XoG9MgeAimCQ1s9iXq/UqrEU2sDKcayWYCMO5La34EvKyJbEqX9HddD
/5nMpaCgwO6jkfAu1wug3IqIDqQL2fqFNQvxLBRwTEx0f+zlxK9uKbO7KsQf2soA3X9fjeHX9euT
xvJvnBYJ9uVJSIMKLccgim4qKFLbVFVsFyDvTweKKDOXVuM/tBtUzpygSavtGj4hKpGzJJ/XCHQ+
rRLEuDLHlcTIcUlE8XhnksM7U4sAjMh+7Fb1UXFrD4a3nU0kchb+xyB3xQA9Ou4LliZ0GfzdDjwV
XJTCB2U48nOEpgSDKPw4HVqbFUX/XD0g2OJHtaG4ayCS2kQ5fKbK+ncAxey3l8EgOofvWoBoGYTg
IoClD8pv/jX7R36d7Ehf6LiJ1nQqsOgZGSBJ0Iuv7icR67SHx8Sbtij1fhx+nzz/6FzIjlwtadwb
Z3RW83H1hRy5H0grirPYlnYM7rPqPfh00pKzfKqydm1OXLlQfPob+taQPLoWgDRFVoztXKh3Ceu2
vvF3QyY93wOBj4WDuHwSm1hY0w64sELRhxj/tlKRI0mQXB71inZfK1dHbbgHNM86tJDPDmq955F3
5x+9MU2gNfWc4kqENjs5qGdi5y3C1aqQ0jYqaEFx5ehY8O8ipukWSNu4PA2JbpGDpUjLDGBtevf+
ufaYT/vpytqUs0UO9LYCOGZgldvpLtBLpH10XDNHn+Qtj8Aa3lqxzE786U3gjpjjVr00Fqojinvc
1jko19V6/aPbBex9dzOpaofcdy/N5VcLjTRQ18T6PlWs6+o51TzZuegTeKUWS9NwDzgld//OiLJf
fwCyvz9ySyV3qB0xbYzi+jmia2QFPC/COCjocJVy9tA5StO9AZLKgbfl6m0d3Ixa0fi7mgf/1Ivm
r6OoZRDcMXwMnis+Jvs+hlXz4d4clZUmK1xLVdLmAGGOT8fsTlPOcJjO1cMFMvxb/8RzbniHNioi
U4REgxKf7A7IQ9nUaLHC51FPrDiwgUcMPe1rcJRlGA8wWd0u/5XO5XpMkq9Nuxb5qmAh/dtbntnp
X20Y+ZscOGJzFXFK7R/MwDxGitu9+VVngFs4LoODAVg1t5o29sdxlRn6z3EwAxtKswk2h/81hTUk
UTTQpddB0p3QurGZxQSRhgeJjrV1iHYouzz/Lr6vqeC+eRqGgBpISpqLSJJuDOvz3LsFlLoee3lp
OilobzHeU980HGHCPgkmhDQIDCsEOAzyzvuk6GNSb8269U3jRAO8eOmLy5uLXKCEw+YTNmlwuMcS
jPcWcf3+1yBPKUyC8ZRO/plu2CfJ9ODtekHmlXi8Hltll/CUCyE5Ldp1Wbcn6Waw9TicgpQ7QJR7
fz5ikZDOZjW3S16zYKHph3+wP7Slou8HhTqWmsegLB3I7jP5QzqM9zsLPe8jHt3ZldsCSiOoWM9q
UOkYvPkH5WldmTbuxq8Kd3WWf/d5bNj5Lwxo2qAJh/DhvYSUbed8EndOaPVBt43GqMi0PTtHXOU2
g4q2PA2QqmhAxOx5nOO+yxkWzxtpJAiTfgfTFDu+vsKMQ5VBst6FTbDksF/FCzve/83ol8vLNh3j
OZAjaDTb6hGdWpifLV54yfBCKDmX/A9sSfe6E4j13zhKcw2PlbLIaXk2nqCEuUsJIY3piTTu581G
RrD+4E+TMzXnsk0r3/kHW5JazKltBc6teOCW6JOrcgWMU2xXUVvMOLmUojKMHbUmwrB003qM2JR3
xXkqYp37YTsvkT5bFoCqfwWrA3vo+lKkoauHecuwBJ9SI/TrVqypV38Qv/mPck23VwONFEdDx4mT
FudJMo53eGPwUe2g7U38DZO9r6OMAGP9B/jY1xO2BetKdMlr3cMdlkwntirICyeW7/gY+7HMNkvv
waxlV3qgXHvE6V4bqZNR9HnQ+tNWkXnTg6/EzOKwAyzZhKQbG0/UhaCx2WTZUqvf+qrDMeH3aH7E
MEBLap2JTDz64/RJIt1Z2018zT+TvuOL/SgC1lk5HZ2EfpU6HOmq5G4qbVxlgFCPJJomCRmcX8pZ
RF2xawq0yiXKnepnUP5PnxbAo2HmQkzh1l8XNnh8hnhw9L5F0PprD5Sj6qm35X175O7YyROn6n7y
EcTkDahZ1Y0wrU5MFX+jEiywPOMLWzRxBrtQFZQSUz3EPBQwDeiiccOz0m7ZoEPrvsK1RqmF0+/P
4zbPwwNKfR5chIzTr9ovvU3uwAY+j/OvXT4aHF4D5/LbR+JhM4nYtI/lAwi7ahVFEOHY3ZLSt4SR
7n9QicvsGSzNDNqGQMbIgXo0wsQw+AwBfnuR8Xq1nHd8BWpkKIbE+gqfcNlwvNCQ0Mb7MsR8a3p8
wZQwUPvgove2sF+RrpmRaJ4i6P5X9BIAjLKayiMwivShY2+hzObiL3j7YUSQ+mfOLfzUhm5tvDME
9uIfdPdWS4LuHGOQnZLPmAP1n9uPqRlMmb+mw5V0It3bFZsFqGOP7tyutuCeb9bYlkZ3f/wzO70S
HWQ8AxvLVJnPrN/9ZWQWmTv7GUWnHW6hG6QpZ7gn7VUU3+c3QrJ3BjwjjWv8WB6UzLl39HwHPjVQ
8BDPATsDwUBF+fNdi3qP2bsGTiT0+UsQ7zg51tXXkPgnAV1MfCyoToYIHKSwdbKm6bOxX7X5PMJC
QSgWG2LlF5sY8ueXw4jt2+WeL7Ponm7f8X0mul65gNSA/RFootM3x96818Hvb1vZZkx04tpGuM4t
AAEgBovMgD4m1L4cna+XHpRqvaBM+QSsbqBwgxYYx4f1pu1r/IL5ElafmsI5whDItV5cKu4sKzUK
SLBbY1zgqSPFl0fham71Lu2YPH9JIjdTeSMD40i2c/6jmPLpBtjIfGwEmuVe79hiWFEsS61ks1tP
Jn5nXeAo3a8jUkc8PBmW1AAu+s33asWy2kR2KfdhOb0e7RCPYaZh7BVmTHaiw/LGcFv0lFJuiTEo
9r6Xn1lZBc3Pq/Oz9uN5vm9q+F6VPeQs7Aq99Dstxn2To75KJwLYHVM6nlagmPDtWnrrKHBw7uik
Mxx9/+a5k5Nr9sHhOX1urQfID1k/yhctDR2hok1+He3XMXWtzSFWWoUP4Bnv1F62Nxa+fLN/vjXi
7wkz/1TaICk5mLialRw4vQiY+IoVHvXlJjlojfaGDtPYeu85re2r1L1mW5+Co01ZdRXemqTiDBi2
cGBvmOBufjnmjZ6o/D1LbxbYs1EQrIvtZ/tEHdNVod1NFmuki4RRQO6to0l1/hOCMp30AwXM+6y8
Vo9tr+uaRiGvQyj/LafZ+pUGEVQPDp6JwcE87LOakbkO+tilxVKHd4oOSEF6zNxMDxOqdAdGPV0E
t6on90ejed/ylsnRsbr4v/7kWkz9J/sPel2DKAFBAzJl8gh1T0IzmCNsmKptLB4rtugglaMdcRJd
w2tcUZwy4p2FzPSLt8zz9DzMCGOnDD5gkfk3vF1MPMvpwUdCfl1pRZmpuI82ah10eDu+aegq2DHy
ja2i/zDA9AK5vgVdZXIvci9wwzLkb9QBjdzAhidFmAQLL9DHhEMRwTYJspB1yDJBOkg5AmW/6szB
AFZwSOL3QovPI8VeAT7D2ZAbO+iNkzgNSqXf9AyeTfo/ytUBoilKqmDMz2g5b3TanGJBZv2PitJi
ImeIq9J7DEkkiSZHKuhsUX/muD67PsrQVLfCO5d6jTHnwFAANvdJafGbfNfKDjvDk3/rGuwXcvuY
ldygp7cONxO4U7NnQMlUIVQo0MUyYE0hd/QZjyca6HoceMF0Ner02f1iKvCfeAds5T1hSA8Dren+
DjsJS/C8KRiigoVbggmrIyLmZ+80uWBd12zGdPrd5ILXAQEYlu9HQySPmxaToPpk+S1RbvLPTsnv
IOWTa826RKQiywhkrAhsZ2LVie/hJe7IdAPZ28t6PyMnA5/3fT/OGV1M1JMPt/UBxxxLXLhgALVO
fbPFMKq27D91R/Sj7i2hqrHWvO36NhR7LBl5kNC77vgmdLdDyW49ui4Mbi8dm6ixdQk75q3S+AQx
W+2DX6MUGOGRjwFZBoAQaCiJb3khuIR+bJj+1ZDiqxLfALawA4MrLdtYaiNwjxcxPUpdqc2K8NoT
i0LbmXxUx9gITK4v4miZLRA/7qC9FKAtkgIIARTTK09zpfA+5/t6YXR9mt9cq9PtjaOXaVHCgzNk
frpA0yW4r0H5aLw2JH/EZX/LQoMOvbG1MUFF7XX9edzbP4bxAjoYqUMZ2Fcfr6a48r6Y6qBrTtUK
nI4TtQb3w8CMBRpl6sZZir/lSeDqURCDX5/1XNq2RfjB5h/JorAu/FcNOWJHbVJgHAHDa99Exmvj
Zpsc2eSQ93bhbCv09MjCSE5LitGh+t5U8P4josprIufdpBz2Ck9u6K7WecfXajlgnKJlThsAcOme
2cmhle14wYgqjIAuIFDAB//ACXawjkhdttTTSUrM0mwrsl4pMiWvqq0wfLFYAkMi7WaOzv3xWobT
w7h5RPf4zMASMUyqsCGUfWertRBeCq2n/pfqy1zC49lVENWQEoLP40xsAeL+Gs4qNYsdPXq52Hfr
inrYCubC8sPEMomfyUtrVPoAhtT2sHlk7mWnHsoOfrIT3kD2C7BckKjOOfnCnNRjBkCSDVoQRXXI
w9Va10DN2wX8kw41+Xm1Llk/dYFmQqUuS37Q+6NbyjKlAuxl5PLlha0r5VCU9fVPt+HOWjqOuZHe
4iARe1c5m0cSbaqNLwbuCCnvcub/g47AtybGiFdhsBDxPL42Gun8SPVzWwzg6sjBQmmidpPoZVIx
GXlPoBMI1iydhep0bHow4XdkyOh6bQ0yuTE+RuO8Vkv6EldQM+UfSMhR3Z+pfDWC/DOSvBasGRep
y+W0xHspLYhclUlkwsgHG4bkZWEjYOHOuVzwyV0VJgJfX1/Tcw8nl8zLyWGMQ95eiZHxi747pSqP
l4J5H4ImiKHGihqy949iy3f6Iz+iC8Y3mDVR4O8hEnuX1+dUCXKDL36bowBwPSQ2FpAqNCb6s1+Z
4yw35lccKjQTmeeK7H/OkPkMbq1In09QloANXUcCDM3B+I5czzrUxFGX9yZABtx7mWykTScTybZc
Ci6nKYblT1ysW3xoYBrlcl/12UqPpNzRXWSEi6EEFHsOtAZTLGjG0KHrZcCYm718qkCkKpacjvme
Ms923L3ACFGBmc3MnCpb/U15u/tEhNKeNGXniCsqq3wLq8iHDAaSfa6mYlFQVZRJBpPPsCgOt74w
4utXRzHkw2rLvlCcS2zYuFn6mbMOjO5UFHQYqUvhkKcXJkWfc5w0kLiGSDdDbJSzik67Sn+62Z01
Ekmf5UwGHQCAACfjwRl1JnYsPRHj2OVES6+fENJ3YRL8wgPgfOf55sCKfpIyMIJ0+/0BA+Rtj6XT
sCoJt3QAGw2T9ZFFpj5JNTfcwakS+ip1xT4GjmJ/C5WIZufk7sIaofloe8YGVDO3ji3yrQub18I+
wMgbWsRSNr7r7PSY5Tlzy2ASM5W7v+DNniZfEYR5QY/nsI+9Ezze4rm0p5QI68l8TCXENBTAU+7S
724xC6APCeiGcIXB0egdj/obtKwwzR0Vod15hqsQX8zoiE07agi3HLsotenPL/xvDYGvTo4Vu++1
8w/RymDwwsndKssNnKkByeCm+F4cIkfHDQbKTk26hjY7pphmwOpkFDyMcRFbCg6CqNhQzuU+KofN
lLZY3tTV1wzTDS3XS8Lcw8Y+SBmwgL2v4tPu7u0AKkU95CZit6ol1i9PmAx14CRy+X68pf0aGV+6
WPEGLbrxgJZupYH0qj2eYq2AcTfKrUKFA7VO2ogX07Ut23jyrxOvykmOqWwsiq/61QaI28YGEccW
fwPBlCf+/W1BR2Tydw+juYbWs0d/8+rYWG8BN3rfDNt4mZp2nOf3UzH99DPAOdsX2OFa8HdSOdhH
WGKTWXfA5DIajvoH/J4B4d8vZB3a+R2xIp2GXWrshByesfjAkXC2uIJptls1xBaZVxyTq/NhGEk6
r13/+naS/8gLqnHWJvGtWOfaR0of8TBhbYO9AYE8QUyt4v47hffCZ8rfP8JWcpuDMIrZfAzOBCrP
WvsJD3lN6rDPVbD8m1XwVngqn7fgyzAG7u6IrqEoH/vzP1Gr93HLt7ipwayEGA61bLlHpK1bsbbO
88RP3TA+vZ9nh5Hz6WhvkCYMBfIQXhohmTn2wp626pqmOB1MEAvHpI8Nwkb0RUArwRrmuPmTQcnK
QIxa55UPhQtqAMkFxbfVs3+ytOdYurD+pCrVpLE5ec7Y6gjgUUpFVjOiKwWS8mSFzKGAfzAfYP9+
Zg7rwYtBXi69nypDQlLTHgW8KS5bOYS04fYg0EPhIJvTp9Ndd5PZy/zgRFG0TsbyLuJKlIylJ1zt
+08YgXcQp0HQBeqf7ajmppjWA2CMm25k0Mn2hF9C9g6ei2B42j0qXqrP3fGP6j+YFVue0RdCZJHA
e9Mvg2YR3xbbr7ATwMMxTcZQYDAmE60IfUn7vW6RUjRH40tYfWUzwGp9H4myclT6ewlIbWkRe9Yg
IvjCOhDM5W3J+jNCbdVmShkInK5C/eTUHAEAS//1mwlnubWHm1E87EPKIZJ5jAUljSwZ/1LTcEeJ
ceyxgxtz7KzgXz2cV5M8F6LjiniobLgpEDabAM2qPdJlQdrxlCZ5FbB2585kB1fxlZ7MNE5/Efxn
ckaeMlHEmJxsvnD/57c4SQbJg6/jHMwIJfH9oqmZHZHflMv9LoxkUzqoASsePD3dMdDn7Sl690IQ
U2mhd8172ButFEFffqfqN7jZq9Uf5wtFkFN/hVYKZTFdxSRoEdQY51EclQR0JxeGf/RI098gUBe6
7MEkN3J0iIMvTF5Rggb5hu8eX75kqcUm8BSeevA+o9PsjUN7QurHxPotBH5+8m3+A4FuiDxR58pf
RBIfH9+6X9Q2/CFgMNCQP/EhGGoPbD986faaH0B7H8m8rzrL27yo/oPNyXeZHg4RY7VyibU5bkrk
1lWwIVbmMWdnBVR0MNG9J7bZuzXdScLlsi2jJxA+nIOaec+7wbBTcWbNrVQ0L832J6KyuyDBnxsQ
QgdfBLHbSSMi8y8BQ63/sOdi3c9GnJEKXCPGEFahQ5oceez0xD44lYqM13rsWHLvCjDekKxm//wu
qBFy+JOm2IUObjif9+wmudAPebNyrvv0xN5RD9g938DCQ2uZOAHCk2KX8MIcvoWrk0+yvZr3S2QD
V0am+oMxJygjXCMAQXGA0JKgnrbAb0snJy9Ty5RotVDUd1m/byHYXpbFXJxZoxHzxX1NVN3ZVCTY
B8WoR1f19Csa7x0PndzpltT81ou19pwnakEy97LaM8dg/S1Lym315O+o+E4C91EZKnJIsM8zGStw
cmo+JL4YNgMB46coHpppPGwoWVCBh6fUa5Yhc7GiUZ/2/KOpAsuTu6r45iXJ9i5r/kCjBVBjNSjY
oA/lzW8zGeSYIFx3tINVADGFfuoBSQPAObXuXZGFlMU/aVTat28YDzl2GVf/4Jtp3Wrfk48qZ0bs
Lv5nLrlWeViG1bXgogKOP7P/aTZ2V0x351hYP8ORPMOcbvYnP2ta+6KQsTItMxHZ4KYfcVVpChLt
5cM7HmQluWpGRLLKQY0Eno8rQBIPNeo7b+Q36MwW+G3GEbJNYnOLCialiOH/p25kB/svmrtxbW3W
H7taYmaiGg4fHJR/5autTQLVssiN4UJfjfg7qN5YOA1SEGbywGXnDQsx1STw17MSJHH0R2ljFOID
hMjByADW7UBrB6CC09/7ErCGdjOURIFJmWEF12fI4TpZ9clUXv2rY50y0MYO/g5v61ceOyJdiy1e
B/6jkpH17PTBTUMg6ywpueS9/ZjJ3fbDgMqahodv/oHU1RiAez+b31Ciua896ApGBH24+waethIq
d3Yo1IIV2uwhtzRL7/K6oy7A1JFkKCXmIwqfEkC0/zn7hyDNS3G3ZxKLacEGLERud3AG+dZNDlFe
jrfzwrqJOYsdHM4F7gIzht0wqrTiO7UIExHQSUOG/9MgqIbgRCzlu3qV0XzW2QZUV5PGnD1zbFre
xN08aRn5FsHsU2DnHsR7xtHxYeoX2tvTSdqnWU9/qeGjCHVehyYYB0on0q1L/kdQgIdRD2HIJwop
mDiBXmxZXSXdQoECXvSbg7MXllaXQbdV1tHZogmtHn5f2Tgcl6qgoQj+YfHjter0trAWLR7/nZdc
+tD/voH1pBsNwL6utGYlvh42H4Jv+mPRbRJZvrUy4ZueVWMxueXU0fiHttZY3lTDP6SnkoI/v6Co
DrrIRvifiHY6EWgYVYFoc+/fzdRxmmUmrWy5BTp4NFK7ubXWVvQv/VC4w21AJKiBX54vPBe1vQkq
MfQ+mRqAkT+Q5NcQuJJsMuP2Qqi7KrYi5Y837W6S5/U5xgPRxpeMst6KoSgApjpabBuFzQySUzJC
FSlmjOqIIMYW0f02BC8yqy17AYoiqiFehIzenwtLHZ5B6pXzo8qEL2/KqpbjNpU/oqTQkJQiCH7Z
YOWbSMdAmi6PRbrBfwb4Crm5GLFgJRj42iCy9vgncGPk8vtcDh3XiiWyzq5KyGen5ZxAWxhzWKtI
OkE/VvuSsQh0E8HOZhJ657RrQ6pCJFB0zrD79PpOWmyk2uaYLR8wQwEHHSHn9xPMYYfvA36dgbdM
igfleYzAV5NLuXDVGIBP4rsMnWLJtJANA/q5OpMKbtgx+bEWx4FC/JprZxrPyZp/lJtTysOZG70X
F0YqGv3l9F6t7uxOZUGDXwUvpBPxWhzko148DYVm/6qyjnj70oAg/zm6V6KiJCjXhVUo4YXDBvec
MhJg9bxkCh0AHRUiiTiea9xbXAn/dsaWAeOW//yEGWQhF9TWmwHySJeW0unyAA7lyN1hh3/4XuqS
B2zZdU3I6OQcsJpT14MzQU0r8S6JcXVMWdEPQFo7kwMzJU043XVhsln94YIo9+XmQyI2z/V8Ei33
TDRs/LnL7ingy0kc81xkCeM0nDYfXmcs1UDw/g/f7JvOB18rS19iLv6RrBCaBFnp3KSeQA+Yz/L4
nmD9xGiemCJVMI6SWcnWjv7xZ6AmZ+i5Xqd4hjybIW6BTmH8DqCSLrqbkYoz9mhkcxWNC83rERug
y+4GQgOLqREw268WsNnCpK2SDHFlUdMFNoxJTLwptlDDKzGdJwiPxuIGEWHvzGG+Xa+yJm2f4X6w
TZ9GBDJyEa9s7LPRsiFQEM01hXpjzj1qjnb3gLroSlRGTNZFfOlOP+qGzdqYFCnIDQJk/UbrPCQt
h76O8VmMibnRqwUCrWxxKv+VF5OX6YREecQOhz22CDEA0jHvMolKW7X/UWgY9IHoNsyg2EKPVtiz
imYElYgAs/81IfhMcbdqvG2hv+uPMPs/xhR/q8xMBEtoTraKwxtj4EcnIyiq6zZx0gdnHozFem9i
h4r1W1BG6mAP1EQrEDLInl9NbHC3PMn+0QRASqgJygy9HYMt7P2NS0PNjtpnAW3yx3mY8fqsa+7x
9h2NbGS1TlZ3hn/Y9cQd2ShMO/E9SCyxi7EhE9Ksx23lKXWHqILU/emHzEzBTNNyDXT/w5Erl1SE
JoJZnXQZfMNeHDNsWZ2i69PiIebebKRepYHevbHwUeyuA/fh/AJlqCtzlioQ8tI48E1CBXjb63aq
/HYM8FXyVrZZlh8cLzONGv2WFGV01Fo41zjrXmwLtjo2zkVnjUXZ5rtq0ibwLeerzR7BpHF7mM17
Cy8OaV7f9ZqSt54uXbhdlhb6+I1rWfmlP8MixccH62Om4u9Htos45+O73pqmKcU8ptTfrpRpHdJy
CM/DgmvO3dbV+/PD62alAuvCqc7tlVeCIenjeN0z2vjruG9LHUc7nvWSvIPWJBS3VMNXPg5t4jKV
oXtnsVAvPTROTdcT0Ss5SV65HkDFLZzxSThE7aRTy5PWLKRV1OJllY8I1t/zpzqyGw3yPgGBEDKk
ejllWbd4Gzv37n5otJJj1wes1wU1MtYkh8UpG7ek0C+3GULCNQLPcMecKJAiIj4ZWmxxiRIPi4oG
GtAuwQDHvUJostvX8htKT5PHYllTkztdMKP+ad94N7RvfczE+GqV8dX3LZeNQlcJn2kTRuLqdpkQ
AtHr/3f5KSX/9SjaI5kev0zyj0Lpf6+CYRpTl7QNx3qcUKlDFgy7M1cqqxllBb1uRFnuSUGRzZvb
g7URUPMrFshro3Cc7fG+Uk79/pdVgzW7KSJrg2wczcLlCfVtq0WUwr6gFeqNkH6+OyFD35ihKni2
tLv5XF3pPWXNvkpmu1/8W9hx+aDfIBiG8v6SGW5pE1UZ6jz2t4LbJvW1PAHkMNsSUHFGx4dWCkHG
0teitDLxi1IfSz4uAf1YJna2YoFsTAYhK3X8ImqaeHNk0h6xDvS/vYaaFck2gXmxdkHj9XVgn8X2
NoRUptd5nmkvGrhgF3dtJsuNXYuYHXcV0fuDnDLFeS1jq9Mjy0L0HGUFniU+j2d0CcFF08PViWCQ
m9/hZ8K6yDLMFiDLVuAGZqx3fD6HDE3XVGZPlOBFTnoAlGTTpIVsJt8dH/QBt/FoYr3kh+bx41iz
RGz4Co2vXdAEOSvF9gQUtrCOzgNRM6HKIiWf+aIIhO4FQxtYMaHmhmob+6XeJuwdoe7sCNR3PxlX
N84t7BqlzJ2YcVjZ+LdkLNzaVLT2L7kBK7y8WafnrKZm3lRb5w+r/Za9zbexArdnigqiwDAaYFOQ
SXk6FogylQyEc3nLlejXeM5YbAgi1DVHOU50fLcyUZImI8WzP7KInbhQEXg8RQYwgvThz4QSFyF9
HkPw4JEh+f7Q9m2ZVpnrl+SEJgtHpcyG3uKHWN3GzTSHLLi1XUgrHJxENGqrvAtNcvv49MKr+4oN
C8+WM5Jpio69ieCoVtu1JXPs7GICp+uXOQQulrT2h5FfXzHkGmYBQvse7jz2hZ2nnRGYjThASEnL
kLkt79s/rFdHTGiTHYXMB8RLm7hGlbzZk6JPF5g6q44L4X8EvFEwlV40cjrZvhaDUU0CjbFWlMNv
Aa22NCMozf/22ELYqiC/x/SavmANfOsDtxTAChszGngbGT/ed/8zrNRDip5x8xbqlddTky/awPxW
7HX/JbHvnCpcYmcpmOGR9mSoFV1H2PCSqdcNmXPAmjfTZL7qjmfvVT3xzUWysAs058q3Zjc7YL42
8R/eeBQSCMr807e6mP5ZPm8fPGKc6iIsLu6/nPG4hgD8kiv5VaJf2s1OcywWgc5vYadjfewsqzM1
UV4vH5MC8poNvpykAbXCatK0PR4s0SPzhhrsbQZFeQpSD/ZmP1llCBvoO+aCze+f0OqGJrl1dLkF
TpGLDFa3cAHxpr3iwudG9PpoFRuwWe6uWfebgcUP7nK581nlU3lEaqDFFFE4VUi6rGso7xFEmter
xYPV16y1eahg25cwah/Mp8C7stV/HmQ8RkCHuigesi8ePYc6ZkDT7TEvAdII+XpbH34fw+QpSUFt
x9WQxVbjomDGFKwc//woTCZQYXrpcF34sjcOtEsA9Rq1Cv5tchzkUj7+1iQiLqJqTc6H8ALJiV1A
x5h0Tb8Dht2oJc93otb91b/tcdHzi7T7ri4zatioiNIM8bC/kcBB1RoPNB/Y2o07K8kvomKrM/vk
nVaXXV1KcZToyvA9yV8w2Y8/v7W4LiR/f4zrdD3t153Dbk2ADaeYa9n4cELD0DZFcF91eIFGRVQJ
Jl6tgp+Hudi2jpv0DOFcMHnV1cg0pbO8kuZ++OxTuShxYbZrd8/L8WdwSvVvIIiqJ/L7EpGaL77K
QC27xZgTTYVqB5dnwLWhXymc6sGEXqWLiz26Fn7PZs23hQaTsVjtIVyocdfV/AKjiSjczSElk5PK
iJ0m7dERdJyqkfdF0YGtgzPwDkAP7npDpIO2bnueY9IvnfE5zSazmqXqIfZCTcB4AJCud8bt61oi
gWTsHF41j0wmyREzZHPf0Dv+TETcJ2c/PPPTdw3ToOtkt8GuxDbUbrGFZdH43px8dMYTqpG0qp/V
js/2khINtdedFCq4Ef0W6IPE1TvVMvGada9tBxN3FBJm2G8pcfe0dofsvCDnnRsBduIqHf2PaiSY
atbTD2UTTrb0ddilp3jGeUblr+GgqivbZE6k1jT4OhjBCUak4Ff6xhmkbxcqEOPeqPNJW/hxIF8y
fxqPeKyFfrvxHy50gMyNv57TEWEMHu+nUPXblVtITBNbaiC2jeFMxK9BKSoZizlb0pWJFmm8MrT9
oYCidOOq31Bx49TaGKGLinAcO4mcittNFuorzsvw65qFlDBoh6ClZ/3YFGoefehcw4E78r/N1cwo
R+F1yL5qLFXryjks1LOBUCWeAV2AfThG4bXeCLhcwsyneF4Yd+BQpwZhbMCerAgBLvyO3f95rFD5
wftzwa45U8PfGz9KrJ5byxsTnX4WZOFQspJ6zPTaHDkUgtb3FVDMf/2otfvn5pDetXdvB6uOkSPE
hJQHMVqof4DLRcfeRFiOzi/rqEwBl6Q5AzG+K1LyEcWt6ubDgssSWLHsWvIwP0bv2af1autBcyTi
Wffip34r2BkUVB6jQv3pPVFwE+oQY5wSZ2LJulIRfjldO7VcvR2N6WjWcmnt4IU4KGBocM0eYJZM
T3qk6DiKTBbwn1rZJWANXIVZO7Y3U5pNRYhgnDsJPVgqrEeT+LylsP74EMd2mRUGnVL7DPFgyvfX
EaOW/GFUnTZYlIjI4JNtCn5yQIlyeVh/tXVhRj1rR+Zr/QOmo2e8mlNN6H4ru0hSFjirFCiz+6lB
xbVx0qkO9jCP2GAzHYctnnhACgrR7oGRF+nh+hzP1tG/n4bMRaeaoY/dOisdnxdLWUqFftiThNYQ
wKLZmWnSqHFc5QraI20SI9OTQ1XuToiJW+mKBkxJxFS1d2rCET6jV8ztci4fwmlv4j6GCs0yWe3/
ZyKPQxw9dPesunqBUjfGMQOm3gw9VIWClH1Ul08apZsf6afflsZP7tCU6S9KHB7FauYZXMapkvX/
5vZVBJHpaL8FaeOrljwpq4TTx0n2xVc5uhFlPHQpq1T+KIAFAmTotpQ0BJnG8JTt1KVci0yaAF/b
slbl67u9iIlzguhrKOX2uOiMK1F7uYwJnOsGzH1Bbxi5qfMBGr3iCuvGSZLPOnfWf5fc6Bg+4tFj
jQCP+q9ueV5SLipqenUtLe+DkEC39HUviAf2G8SDNWMSgfYkh3eVjdUJwX/p8W9tFjGfsWFD2zYB
VGkKkkKdNRbOJX6TKyZdZHFBdKWoV9ytVR8cAAW4trZ5QGLk14HSDN5xYMuHfAsd5VI+kFQLKwUC
erzTEebrBHo4ktith/sCq5X8UYKUO0C26cOyx4Xg/pSUVXvrMMmQOhlkbZ9dFTOBFkS46ncw4VYY
WW2uJj2w6FZPNAh/VqcrbY4u32zg4eBlUQiJakkHYH5fzQgxT8YppIz2J7yiJL6I2RbJCrhnjrKT
7BO9Zr/FANhe9Osb8jvPkRxzoCO+vkRFAtUBwhd7lcyzisOzL0TKuazqMm/yZj/RCw6adHBHwGa/
H5wHxjfgla9Wp0jrqaO5TsmAh0emBYdMlJAbV0iTcnLJjWrpVePUmi/LCeN4bbwi6F0VhC2dCLYq
Jk+N5HfeqR4RcPo8BI71k8TMJU14pJBkQ5jMkwgQwLjEgpsX9zB0wCsBdr+X0GSWQkGtBx/BbKbf
9mZb75MxvgcxVEwt/PzGEabqom8xm3SOm4N0jxv36AKcYhEdYipvLbA0tPEP1khExAeo+cLVaa7e
8QxxIcapycvyKJ0L5RD6zG2F1KuvUCeFt2sdBVyv7owo+ZP8OIMpvGT66xHhFH+P24iiTvwFVDyR
5XlLUw2lOA8TATpznFB+UT5Ghlb771Uy+XttTe8YryUd9cEh1nuwFZ3XITNda53FDg0WIXy4qnAd
yw3mBXTA0Fa0JNKIdQDXGVUDSQ8t1CYqxteqctq4wpUyhP//tG5PwOt5X6/uub+Y4LhLkECceXDV
tll5jX7P61Ydae2ElxRL4fMy6WhCu5vukPFCAYGHqyiT70iPGRjrKjeqhA+4khzqJ0sd4m/xqbY0
RNpTaxIUwNZJ8jl+4x4Hv6YROiBXf/O3teFD8FmRTcbQXqyiiJx5CwZHxaamfh71ZSKT8pqROgkR
YwhsQN4P6lv0qUzmQy2q1rkgS1R1GMwGb3wOpgyrrJtQ4sSFrGvmgljVuZwSx67eIzfKlI8PZI3N
GPn9y6LWx2//PAx6g9yqwqMfK72Q9YyqHt+UHYVBcmn7vbcpN/AbUoZJCwhrwZtQ+h6dmD5q7BOe
xn3ValpSvsLxBfjIV9E3W0hWarMtEvoTNPb3oA5qB6znPdBdUddCxKd39+VCNzSxTKepPydASqTQ
02nGkWkcCoRaDYSj+No9/Rwk/S5DHH7Um/Q+iAUJdMF+2ORTL+RFjBSbEb1RL2IdnQ0shsONEvJj
u4l53CZfoNz0B4RDXQP66oM6Am512rEv3/HwYSlFh/cNXCcg4aCLZA2Vy2zqjY/4f9R239cph73d
LKNMFIWcCyCqlLPTz3Oqu+GyrMBRf9R2t0szhB1rkVQaFn+hXoDY0D29h7T6EUpfjywK8IBh6g+e
CduIaDmPXKZQqDM+ec+n46HjEZd1GEntf2vKrTL+bujRKUMKtUCckoJ/5KRCPlV5QOsLfa2oHubU
eHNZbp9rAOr8g4kqBZxS2yvczCC2ZCt2FQj16Lc+0gCnXnvg58o4yJcHFt9ebI7HmZDJSCzfvSn+
6Wqec2OdNhR1yUblDsw82xH7bj8zltcYXBSz7PxD4guwK3NeQsmJUUjKBe9llsEVbqHvZTtShDvj
iLzQ0S0HDPK640/jDg4gfLIr2cC9MGi3G9+hDYMNGt2SwvpRAUDvb0nF8hUM0omb/o8E3M2ggm/P
A1nih1t/VnsRZLgn25noqQjhl0oEUyPNyPCrl4PQOtpX0dK+9qdXKKBK8+RD2lzaUI7qkYufBL55
aEGMLr/y+Z9wZ3uX0y2TXPDqTCiDs3geYVV2hi3rvqhWm8ONEzLXVffzNCDPsYKgM/uB4ThHL330
/CpvjRlHn74KF/spcTo3kMfq4DLQRlKtgPoT32wyP5HfSqkwJF35bsDoYj4OUEImD0TGQs7oZBSK
trfHtbsk+mcG/nvW0OHxsWWg8lWqjGAzyiPpuZAsAHDQ+kwQ4mbcxajEx04l4xmPvxbKylVTcLJ9
4HpVqMl2dMmZJK6n2LW6w9gWipbYOdPt7QKdYN9oe4K2BFAYNS0WNnZJxR7HZmQlPDK0pX0LdNcb
C6q0flI4GCimrzRSxbzuaqunGjevxEEgMCbtIeGqjV450l4i2JenFVqw9G3qC3/ovZSDXym2ikC6
0wKgjcZBb9joeKFTUWvwUx9rxdeu96FyU9fcqQQXDj5IVpnJ7KyReTKK/nk8GjoB7idIwO0JmqOs
LvGpIbtJnorg6BWuMfza3IjC/pfvJBa5wt83VVHonh9/1tuBDdeRvOx3SEzyehZinjfWgccNxJW7
Uz8euTTPizzfdO+AcIJ7lqnmgHtVhhfjZ2hoIFU7Dg619qEPfe8VI+p+7SSkJdPwaAa0NZ5qHTCm
vsfgor9VS5qEeWmfPh0wvyvyRv6NnWpRhn4IBlh4h8wRN/zODvpwtpBJb6wNzxs+ECKyxBuxQO1k
iNinISeYg87R6/pZ+wQxC6ZGWXLPQ1FvYfL3n5Yz+SLp4qXnc7vM8/93GgO0XuVdoVzlSrEaHSXO
v94qMXfgiyen44iw5DQkOj0rkZaRrQt5usnGZkD5tS0i9gAtHUCE8gQXf/C3niq8qhweCahz+MB+
vA9JmiEAxb8iQpDy+Gdc6yTGO7Tz0F9SGzTC+WUEwABBWdP8vnfQ3AsN7wROpSkny4/TI3OKxLq6
SS9QhibDxAI75Tj9vk0YQIyBx7sX72f1hCSmnPHtMbrcX2AuMen1TysV52H53liU0qosIS2gDtgO
N/AhKSnoTzPE2WXefRN3H6DzNRa0GAst0vRkAyeOK94vV1ucsO68ZtMihX8tRo/LO2qvA9kx8B1e
dFvig33rsFz+6qc+KfsajZ4XVWizj0PXKbqxzVMMdoVQ3S54+xMCts3RZ84YAv9lGsCQZBDwBsZE
wgeKoTlYlPvT/qPGDAXa840AN0W8+YkxzalPJavj/pnXUy1AOJ0obgqK/k38FlL4RHhEsz6YY0xp
k3iNJGvFuhiUoEhq0I2NRNVbd9FEmCy6b+3NuIEH0pUkTxP3YPzHuHmEOtbUlBnzGmJxT/O8r4OM
v95WFwYcuFAGPfrb70zFbl0Mx2m8ylmSkoISnLoemj49reLKHPFOI0/+UrdzTNIRyFr09IOBlslP
pHAnjWktOEzV5umt31nBAOLOW6gcuXhv1IK6rLZrt8tSCHBq+QQFrxAJq/YmKLmd4tKE8zikd9dY
l59Os+02wwVX5X88YMW7/vf2auxEFE2OB/blQFewEDb+m5O0hN0GC4J7ZDrGjqmu/xNG7ms8MwnL
YTtyW9606tyVS1pndfIIvEDawjXOWwvg81j4Wd2gIzPa1cy6dhxolqQEd9eEMOEkXDE1o2VWMZgS
cf3JRaUBNeGS10bX7NS70V09gSqy0fnh2RxGHcnQZmrZeiQcACeug26LGPpOjaQqNvFzIgwQu3v5
KA1mKCtD1sTfa6McmiTUsx78zFbAClkhu+HPRQA2wNXqKSnKjavPwE9o1BowCHvU9L1CE3RpvDGj
0tC3IMmuI8bl/Y7C8KctHRbGLBMUQd3XXbgzJokJrd/zAXbnNFabYj+oUv1AkYptmCkSdFxykNNb
7e+ECXS8QzP5+9mjltKfxgWBUrmFZn2hnDGy3MYNXerm8NlmnZdhZWUj83LmZ1Nc8gTaRpVhSI9T
6C9qOZCypUnubxmpuyOWD0Jv5O1F8Q3OoU5fkC3gXQpr66SBRYXIdJKxgJQy31QA6JEumM8Yx8K/
NAhLxrPg3RLXshrJvyM/uCkhqA7CxF90Pv+2IZe4isBObLvMeJTclgOgCIQ8S7cQffQbUQBHoBVP
s8teJ+szmNZR9uZPL6c6o12qNKv4zMIqYhdVgi3+ou0spXlORsLlPkNoAsCIfHNBxVgm+UYllBNh
QEnmryEl5wRuBe+w5K6Fwad3t7GJ/o6Jy7qK7Vgmk/cRzcwJLI5P+kp/2iaCpBqc+WaOXwRhuh/K
Rb3LL/4ma6hkBOLRjcNe93jJW4q/Xeb97J82TdjLwWEZtKxGkhZr10QRuN5eKLtbZNqueYQRJUzt
Bqth8s1rvpYeOYtetVnIeYYNQy9p8PklxgpYAmp+43FizDFiJg0eRgUEoSNAD1WhQ6oxAj9jVggu
jjAShNQVstY/LY04By3V/fHtZIC5icsyvueBcgV56AqRtpWwOgJKpFoCL5s7Y2czS7wR80olVPnH
Qkfb6rxbgJV8n4mo5WRNJhSv6EYabP4pCXgJKWdSny+5EIrGzUpU2WUxij0CfYTH2CbJ7vcVVG2s
4Ng2/u1SZFtCeewN+zanAaKLeZivrQoqeYN7JRuaC9kZ1TytSz0ja39DAlceeX0r5PGS1J2QxgD/
ikT//iK/nRCYKPmfY2w//XFoRgvFQTzeuq5V7TKUF7Lec+5tVQMKFLxNbz4lTPHx1kXG+3J2qfPW
Pfu3I3t5foev70CvzHEJILYEiOEV8C204iSJB1fhMGMy8hy8faI/JQNKl8BJFhZwhvmY73W5v0RU
LjsP3O1L5j60Sb64B+ms01q524HWAUZGhyMh4TD2BLn635EGjR/zgfxlh4iNSWN+w3AP+rRuMYf2
KTaaF4IcjL+4d9naoh/fX+DQbAUu9DxYVg0Swun8SlvY2zRDi5SmHoj6hEuJN9SqptRx659Z6SUx
ROWTCyORUjrDfTM2I6fL0x9KJkW/lwnwmomT/g8e+VYyJ7uQCV2uverxzcUS+Ylfm2psEgPf0GQx
/CVxpH8bmy8e1WooDk2akL+RIEIK5eycsTvUgRIptHFFE6ppe5zVBSRz5vwc7YFrf7LHCXnZloBI
aMh9X/hUJ29eF2aAcYe5dqp+1pkH6kNzTPanRUOVk/Q3Hpc6F6vgRBHvBRFJaGVxrOumbiBT+NvJ
hUfjU2xTqSO01nQzqB6g+Dju9P5trENs94J2dBGYT0SYUQMlNNMxLCDTVvJAJMvUo60rX5glnN7x
Fbg52CmezdAEE8h14IxjsNkhgGZDSgPF4KsTqsMTZTJSu55xn3hgIFaSwe3Ym66Ac7WBhRgZ1ddI
E0tsJtAch+sKqe3wMj4QFX69Ami79d1yvUc4tcKIEnwE4lOOvwFf9NN7jJdADZmQdKSKCIjkkGtY
1gCGGLg1zvb63nShzJmjbcXyHs5aIBPQ891ic/Z8uiFrqQMxFwinPVcUz21XIlsWvIES56RwJk9f
97FGYhCyKCC7fQfgOmr7JLyEiaUH7dXaNtWOmLmNK2+QDK+xO3SkFnwijfUQy2ec8vCxsEm8Ua4Z
SsbU0CbGbDoeF2CLdrIijzBh3pHLJxXHVtKvTWQ0F1XV0Noh1HNfi7QyBYPCjYxqreuCZ60R59Vm
1kmpMqwRqiMjrLmLgbPRu4hNX3+k0r/OOsn7Y6zdBV9dpdJ/63C6K9OttQcU6luINcke/GqwXWCJ
mgnrYU7fGQy9uOF9xXcgbgdpFCT3WeskAzoKDLkwb2O6JTvX5geDM8FNMjMI2iQWMgEZPPFzI3of
3JiScOorZFEK4jSiDCwvhDizwb5MM+BfGTdQpq4KDpM5NGKf+Hsy66qEgw6NNowvumPwKVxznrEe
SGeuRaEZHYLhOtCqP4tnfT/SeA3zIwKJmW2HNC+jNWz4XoIuTbyqkmwkZQ8RBmfDMhxQ1GEjV/3W
pOet2pWQVLmywJKJUGtxshL/PVb8uZV/XJZgecGQHegQ0HDI164B2Z4HcIGc0E/8Ww4ScSM31+ez
wO5Dv9PxieMDtRzC7TpAwpewoMNxDzyQvWWWtAG/DPciVAXH1e2eKShoXgDVaBIPw1uVAfeH2MHx
K9yrfWAv7mYrfGVVSBTihlB9UuVZSkZmgIEhsSVi0rKCTrL/ZV0QYosBc8vjFqulllSrOc81TExg
UwC48n9GXkYz8qstHc+pQ2Xdgw+JrbiaFCwraoMXEWXuo4zFP+5QWK5K/HrLluUEu8MKcIRWxWWm
ZjDynxO2scumJdB6+gnrqm1aV/9Ao1accaVMCjWFO7ZT9y+lVNIL/6q2BMz+T6io1IoC22JE8tFx
32/+WzhDmRFilUydIfdnyjg55pu9ZcH46VE3XHk65SRjC88tgchgkdrAPBpuWo7wF8kbm4ynP8T3
25pw3QnOhKg9YVdo+/LXZKXKF5S/a2oUyzyyQ8D9lHO94CbgC+pMamVNdCIFn0VEe3RMjD1QbZl6
iQLdrU53caa2wIj7IiGSR7jmhHEXqZNd6rj1Gs2XvlS2j0gMLE2Nyw38jZuOGs3h1xLtxWG3efN5
9WvLAIhX5W8UM0YOSBebp8evv71dz0208hNnKAvQTXlud0GqPmXqgEOPTf4yVQ8WDUN1zOLORaKu
C8343XYLCmMiL9gt4ktWbymlBFys9jnv0blBZQtZyNaf6DGIrpnf29hgOGMZv4wAaiOqIEscm674
iftD/fnE9KCn6wlA/+kUsE1X4nZo4H/nqltb+aci+IO8786apUBrshPVPBSlofhwsn8KGEdGB0F3
TehAV5Da5IuypScaacczpdQuhXMp74LUTkAI4DJkJ6nkmktLEHlNi/GIQzn+oqRF2esGjq62iyW6
y2w9VyyqHHaX548bXhS+olPlZqkFj5XIavfI/+JNLqQtoguxlcjlC+yhX18c8P143Q7WTqLXdmyK
qXZXrcnf9jr/kJKFN2Cvq9q55cvdO4cGnPTgyGg+4V/GsrZ3/yrisOpTj3v1xoj+zjQijA0plTFy
690cPdwLPEcEMYJUPCkXy5hxTDa9yHbMld30g5MHKIn59XXIiH8/+hoC6sHbHzSUj7Et1YlM9ulu
bnGu2yxbm+PVL+K3ySYaWvlpb8JKCSuAjH+Hirh3SZmslMG2yracSOuAo+YGVOx4sL28GpcnzEA0
014cY+MS0/HoeX31hcNVLiKUKDnmhwceOZXYzjZ8TGg729mqabEnUm2pLa8xNDz+NRhW7sSjns29
l9jfS/6mHFSRhkB0hOa9vwZQ+BgphgdwDViYby6ge7ZUDoCLv/0XXboMzPMH8dvJRQ3BhTQTuMfd
JRJ9et1IOU5f9MdhDZMz42F5DTGIh+EUda5RJK2YDbTlC6To/lGyiHoWp/LxrDgT2a4y05a8vDQc
Y5psobVhTLUJtVULhY11kd5zi5d1QiH2spA9G8U/ly8LhSRYcP30D2Kg7gGZrPj4RXOl5fT5FfuS
5Wq1h4QXuO+VdI9GGDm50rbGqfd81GKX+nSsBZjoBNX+2VHRDSUVRmnywmKUotDu/F2l0xVFUONr
xTDFhRprme9lfnTPKSrdtqTl1sFhD8K40JRPFFwmpigLLPbJS1Ae2ipII8IOVBp4Vr8UEz0dqXUH
As5FSzXdM7CUP8jteEB3zr8ltncf0bWoCF5WFz+bnKWBckwCZV0B0OXnrR149YCJGQJ4BUzXFAy7
aPCxW75rsw+o0C79iIkBKtrT9J3E+KF+zL+GbpfxJ1DESjVrUs8xCV2tYzFFER4ylf4XysvHLYgY
luTBQzCos1WM6PlYiZ9fBSvHKfVgqqCYnh8NyY1VSjgVTdPB/2qIDA3lT56wXJobJbZansu9zATP
uw1DLfdwTXiz4cUFHeAKQUpsjDMZKWDrJ2+UKNkM/phRx4tDzSrI/zTsWDgzzw8+R9YLvM5ja6Ac
rgCUG5noW5BnNkqmuplmkRyFG2YTfx/fOyvyVGcrvHoHSMLhQP92oT7fRAeXzp/x6jgmA1zVvMqf
gHjV71bKCvizGjVc7Kt5i0BFVEZc2SHV1Jyn6fRqxb61I7Gyo3H0osWBXfXBTx0k7Ungk0ovcZnH
QFHoFdyYCjpKSvSPSi83PJcJcUG4bNWSRSflmjIopx9Ts5ZniaSa4UNWqbjOR+r0fnKxOFeQ+PvV
pggeTV/ft1q80QvAvv1Ck2iN2gC4S9LEDgz6iq97M8UW2ze6NRHkYnnOMnEtpnLsb6Hv612CgFez
1B29iJW0nyVqnL6prGTvSvDfFtIBlsVMcFOH+gPluy0vwcoySHziwmwwLZCQkoq3EVafVATqTypw
LFxlc316I1g3egv9C6BlNKvvJ3I66H+JoEJDCMjx/isfcPPl4Hkj0rA+5bqKxWII/akIPQcX5S2C
4Wj1F+sxzRseqtfv95J3FWGZoI9JRBhnSMFIG2QKBuEzdlBhMyJYDwmqG7mX4hw+H1y496Bf3UQp
SV6LTTTU8qRK1DyRTaFM/5MsENCsH5nL9JV3VLBRMU3JqmCkmDJch5RD2ZMmQeBTEj/GwkdmwOrQ
4DGIwIveXzNp1axUtgKhm8Dec65xPX09tvmIVvhsEBOI8/oyhGc4VJl+ZCPdCQA5NS5i9Kmw1Mjo
H3iuQvyiqz3tcoV0DwF3YLdZ219ja/xyonmYpEE6hrt43bRWqSMb7sV/Nv75jdP7/sb12SLoShJy
lpv0QSMFL0NQgjy2k84OcCdH3VOpbr37jinw+V30UpVMISTliFlnhQbq/TMKILs4sPjyDjkEaavy
sAhPZukwFkaDTNk85rnzfM3PWGMfyYyAq5MDppsFTK440wn8qBJSWhNzyVim3g1eWQIUo1heqXQw
Y8dDgzB0T23AKuRJ9rEggR78a0yoygNR0mIQTyOXnIGFx5Bn5nBzNPkytiWHNU6KALDIF+3aijA3
mCfFsrGzTolXg9Qk3jzDGZHo1WQSIEvsUiqbuc40HIsKSjgkd7L4Rb69P6cbbVd5BswvwfcfZQo3
Y4jy7EVWxPG1yRqu4eaSxycuuLNtdfgun3BL7gAc6q0LzTThmryTVaKonL8MHp8v8PoD8tl6rpfJ
mQmfl0AeDtyrQbclvXgSC1X75v05SLyZqcm4NUSTNOsNI2PQt+suhA4oSbGQvj+RgyAkwWfdKxPK
xveXgMiQ3Heg9k37r4QEYPFJXzwtSfAAMzY6qXtkoii9KOzm0UYrqbOx716F6MKdh0dkY7LGtB7w
LDZjw4hYsfR7vLek3hoDiNHMY1QiCYJyUsKfWVpkFOz5HOH0yTF8Mw2EJlfgbvmWoRqO6uw2G8bk
zoAc5iRWN6sBuz+OtUM28IViQIL3W3qWi5k+kM9M7VtGz6P8hd1Q+0zhhf/0ag9fUzLHGAgvrWJv
u2AkmU+geQb7IGnTR8fKGA7He4qXws4WGH2FjetZKuoxOUF5Uj/zadbIzIjFyKSt6r0Nvkw0GP/p
pCdsYDdd8NdXFTVgOh9cTQSYBhZdJJV+m76mCWEa9l6/f/4z2xhlZ4UpxhdphxD1PLMjV0K2imCH
pdSoMQc8ET+IuHlvyZzabFgLGr1IT9AKYB7NSue3vG0UyQWLLquv+9VLtJm9NLI2S9Vq3b1i1HRs
KQP5IDJT4HyUeUWHuEWeUKJkZUswnYXYCp78MfCZTmK7lTi91NR/ogIipuGcyGQwORCXifRpQSFZ
k7ac9E8IUqS5Bn19thjce5OJffJbmBssPWRzA7ERurXsliP3DL3A2tW3wXNWXPc4Qo58G1qracO3
f+qdH2jIMBsqNy9TBls2Wo4TeIkhtzL9al0p/M+phrLH0/6RBhBnyBt7RvQuz9/uqkLMLwyRjmvm
bQQoT08U9/mpK/AFRJkvFz4kEACJlui/sU8wITES+baxpsfBWP3hTybsCy7PPIgd/JdI3HLRhhEi
XNjT2zpAj1jVsKESfawkOkrraojb2pF9MCNQAYuXQr6Wa1gqOE6mx744cVdyRhak7Z5pv4Qm2IhG
/lBQn2MeMooZx0uLTFK+sHfZ+OB74Iu4rhrMHH/WRd1kRtAPzL+PwoPG1UAuia6h8aqjqVmuMFto
mz5qSa5kwBLu+Kb3/5RIyj/VhPrClDqZ+AYYj1a1SWS8gqhDNWipC8w5kVI8yMwt0FyhX4GT/+tf
WO51uy0kSG1tpQwZ+33fD/jz41zSoQATq0y0C4FmYqzR3DFQcM5yOmUQNZTNB9slkwpC0O+m3+rJ
M9zXKnSMcdPwfmqa4mTotCGFISEUbXZAt/3H38HjZ8Fol2T23ZDaS7iAxPjUiYUhjnxnNO5JIqu5
i5Xu4bAvg0XgrZw+dRx0mnUmI+Wtg/XOs9KkBVHcDiiSmM7TMopahyzCx1PwzNol72aWq0eBCmO2
HamMxCTbI2gzH3eOmRkhNR85/QXgoj06EZpiVr22I96mdsBOYONGsxxaWOJaY3IBFkzJA2ZugdKg
shLk2tSIM3j/wrc/8KYy+LMsaQSOfJuRHFmh6uNr1d1Qjz4EkfZlD1Y8gh6yoKOEfbFY9NETEDOq
TSF5hAjnHfj1PBkFbOHl+HPzqjygtnf/sGokhkW8NLNea5/krh62gDfXButPWP4dnwKreWKWQpSy
dp67p/tvWBbddvthDTtMfLbf6MR1stFI1Kk6kcw2bu2wiSMC7w/mNm6nGSdVOgkTsIccg+XcAVl/
wFvaMvRxU12IMd/LHG9Jiycy+ZmD6itHtq4+OI2/qXuUL2CP9KIA6PeHVVNfZ6EbxGsjKw/Z7m2I
cU8K/tryjUddem+z23Vn7teU+03A4o61n//44p32n9RXv12Z1I120TcEBrJdQgImv2W10GvHm8WL
Cw8SvXtB9u/1j4v5rjaph9FAKR0V13s0GSbvPdu7HI63LdqBj7OjWUpEa9iA7qv4ZgRqsjZDxuMq
WCiT9DsFUp2kcicdKb9e+nXaiP/5ZlFryuk6Au2GcqG7hvfppk5LjcNciI0WQPpE0Olo5uDcqw8W
aAL7TYhCKkGaJ0gU5npC9CBBJ8nuMN8T8qaHet/3g6MnBMiXGceSnbDI/sDj4oJcAkXb0w6ZTXiP
4rSAToLwssvIVU0ZvlMkDHZPIgTx3NlAQgAENQQeGxPF32xHqyRgq6cfCa7VgzDjFV66rpmdgUa2
muDh+aLokRvyDKbiHtnbNoIGPoBXq6CWtrgLCYfcGmhgO/4gP3EUjuaAqZio9gZXU80BdizYh6AE
6HkJANFIijNZB363emZ73UJ8KKQjZescl9vFEsYpgekNlSd2pD+SmhzQd38qFPFUfz/hemJeuqKj
Eklr9HXavHK02CIknrUnCv2Ip3bSQtzpZHUJKKH0NLiGEz4DYN4H8mikxs6ctA7FtAPO450JUPnf
LFCbP4xxpjFi2DRO4iKYawk9QbNAgIxYEpe7LGKenov8RYECCSfWDj3e/6RR2G/uyQ7bQRkVavl/
aQq3KJoMARMwPi9KVjsrsmm50hVEQPRte6JKadCTyM6/0A5hG2DUXGm22/tHFM0rNsGSTEqxU58K
1sXLlPmV7J/b4G46KG4STdQoBBZP0uJ9cmhiRNPNXGCMCApXfUj5SvDk94YX1sX+YkqDTNBfVPCU
+wEZpqHaWuc/vcNzD7gfYhSJkNPj62lhHw2CEMV7NaxZ+hCPgTdr8gFvv5TvaVONjLjpWiqWw9R7
zUh/KUaKydQ8sPxmfQmd8o+sOPB8katZyZzkrLt/+ox3Zo1qoqzwgX8yUmR+N4fisxuvvyIwMkm7
mZATSYIOatDBxKplC1TzKHHh0/v9ZHmcX2qP9cIvZ/nUg7v2f7KzBKrEln2oFfbT3A6AkLFULAog
yNGm6Ilb1eL1xjgMOj4BjiLybM2vdDqUNx8cCgJVuNlxlUiFBBwhR7KHKM0EB2wYdhkeLtzGzRd9
vJ+c1FhmL2Ao6Lc/kdgasRgPJWZcGCVBCS/MP1zrajqaRZvnyz64YOKHQFuTmFy32mk3hP7QrA+O
8Hc/MS0uY904c8lmTUMkYReDTyDhuST83/mJ30PJXLY7ZOOqFsvaG/mmcW1rKBWIvBw897QiyAiq
RqESm9ImuaPFHIil+wgenmT97lyqZK3DCqR3eQdp0zFDgx1yGxOtQVbFKnyHmJdbzTIY5sb+bzn4
yUsZXoMTzavkmfAbinvmCexE9vvgGu3+6O+j8irvwmcR5bS9W880AXvueaKEKnhtEkqkNqzj5qRN
Y2b4061fUH3soN32p3s2mWuzSSvlJwnih3/nan6Qj7VbHciEcpgt+umy4QBPUMB+hKCjQE2DL5cS
f6NRD3nwZHORaNtInFCJC5eT4o6OJxCQvld3wlHbdbgAjIzdM7Hp9wBIMoluztZYOUdAq0zuo+ZD
nrsceg8nc9xRQOzeZLlNmN8sHN3jzJt1fwgSwTfHkKwpezbmamQ2E1rsNdYZUz7bSwbk3AWzguam
/gC9i8VRq/jtb96bznP1Y3ptSR5yeZ+egvHTihDy0bByyVPALhQJIvip9wkVMxBlVA4vqOqwuAeY
rqs3GQMtOTqce1RHk+bZvJSjVvDsP4essz9pgyNIp1nXjP9vNhCe/hUpHXegBTHuSqaJgxsRCvtN
RqkTvHwIgaifI3vJ15oS04X1auvvvl9QH1PUGEVVG9bK6zrVVzdqYWkOfwkUMTFL6XUSN00LdyVY
WsaVzO+lzubYSy+s0yxufFWM8hW+BpcIdXx4vp4+0BUPtxoSIs8dd7Uni6Xbz/jw+GLeZMbPLvmh
RX7kbr8EL8lbaL/sQYc2u5w6Kcx+KkzyoNyf+P+dfyvk8ADSyGU8ne0AOP69jOp4jBSukbDQLfmv
gtTeZCqvRoDvW/WSPnJxFwl4shn9UvZUfMipDChuDyMDjESRkBa9kbhplI2liYHdTOHSs58l1Fj6
2Yv3sXY7Ogcdwnwl9SNJFkwktY/8GObqL2RZlhvRFJCo65y5/MFm229TSgw4sd64VnPNR/VccMGj
tVYCAHe5BL+0FYJ5QVft3HqdZbpcv/kFjTH32BRDVaXI1zsV5i3wn6Jne7mh/XdBivwnZ7F17kYm
DpvURob21oJpvv6U3SK0ZBZ21P2mAy0RZypQFpQiQtVRHrKSrJAVXZMVjDI9lJ/S/pCZqMSl2/bl
NhAbtdnM+NAjikmWfYOQaGzwSTvy/2AbRmDZlJXmXxVTCmbpLuqVN4RRoc4Fb2UoiEwunP4yCW4k
bSazPIMHld+CynRl0FUfcMFotnYeVjI4Llnh3kf/ecih+k/9Yr550DP3m9S7p9ZCj+Zcvw4YFL1r
nSX/7rqeU97X6zW6VJSYqEMSu6RJAPro/9Zxb3GPfP79zzpum+8b3rY/DF2lnv8z+LF9B20vDXba
msm4oZc/TrV2t0zzEigEEXKfwivmCXDu3a8UsD7L756+OjmLhB8Z0MjW7f+zuHr8GjDXKALVMiSs
wSFaSdDO9vfWOrlqKWAS9NYb5N9YU740lT6O4pXEkdmfXWUaeaypSUKGn9YdijLf7UNZuMZ/KMyL
kRVCSRgEKInOsd0Ua1yZ7cwIYy7jnnXkqOrSjZVDOquBMeW5uAXT8LFjJIi/EI3gC/MWvaolOOpn
v0HeDSfoYWtVB++UC0Xm7YVttTexBJ+FksORbIxr8xX0T6zgcf5q2F6wDXarH+wmvCCggU5B+zZk
ZsC/uVWw0tYOV/yvWilbHgXrJ7iapE+SXM3umuAVQRdXYg9sdwrhRTfulYkkdYSXLrY5gxryx27t
NwahRuSFC54GDM1wkHrgXwrk7D2Gey/lCL/30hQf2wOZs4XpwnRR5sO12zyZw4DbICAI1VONpGhb
WkRjH+Vp/xE3hnHtGAkMI7yDyoJTkVhiCB11WM/eg4a2vIvzryW8hiIhDQsVgOURhjvig615QVx7
w9gSTNQyOYhIZnXI/f69IXbUWPIqzap39sPeuJTZef8e1z3MsPvhGoE1M+750ZBq277cdNFCPDy4
ZcsYapUnw7qQ2FU9P8KhZMLFzqboZGcQSePcausZEoKD7ORudtnHO6lF8BIqfQ4uIomiWpbGbK88
+NzyyXliZ5ItOvSI0auxoIyxem2s3I3KVmk8WiswAvHW8pi/66pMVMRkrLD7yTngcm6TGD9+T95X
nrpiQTsFrUn//ot/NUqRGDFIQ8ykDDFqs8yElpDwGNcDlgso182m5tTkYECH1JaHyf6buwoBAG51
MZdUQkbwmVrW9cxIsuGjsrIbTkRjASspizmlrkfliRxzUPztE/Qn61NZsi4cT9fi5GdynNZCJle3
HLlCQOmCXEkew987Pu++J2Bo72UEM7fpTAnQlgEssFBRlTqp/laerSY69eKUv22rLEAI+eMf6E8M
JTsI6j0LbwLTL2vC+FO1m3OBflnVP7RmSnRMe2pPP/NyrNAaaUpeIuM9uauSPu0DEiuV0FpnvuYc
spcYGpFMtAabtW2bzKl2QCmvDonN51SFR69CT+LSEFOMbImA+9w+j2YYI0KTFkwiPuY5aW5kzmRd
1DzUrJdTrB6hi+ySQOh+8jLIBupZyvNJ691eH7hxcLwKRuDX0sEUtfkwcq9MMo05bP16exXJmnMA
09kGXLR0M9/RXdXjbgdpv4LzVkLhpcM36wq6BzUF13PlZIK813syZuK6ULx+3thMeXoF5XsvSKyR
bfuRAmhVcXhjmx1WtNDDuHQQN+b6ydzS61WZBbP2pdsIR0q1PfCROe8ZHTQ5jVnAosgZT8AjPfQp
P2q2FY3V95VonCsl0u5+O8qDZitolQTJn1Yss+vMRqqcryOG4R83B467uBg1/VXIOXp5w7a6loW2
ERcpEwQ1vLqABFueVxzepLJ+NvIMuZn2iGilPTK/hpqTRr0O0EXI3ni0kvITtYvvHXkH8oBVRkqM
2klTljUCoUqy5aCu2jl3K6Pusze2X2DRGf+N+CyK6hYcMBgOU5Z5G+xKw+RYR5yRehe7+Pw5/ciU
lEOhyOME7MmjhlSqdRm/G/CBAn4IkDm2DRgGuVO2JgxtzsFiu0+koDHY4TB7AiNMTlHBw6kcAeXY
/10JjgXgdPJj4/YkVFBqR+MrJ3upguiGKEEirlb3XOXsFepdFEjIQMkbEGgA/1qwZPO6Qaimjt8N
rYA0X5Zok3zVG9gAxE6TLS4/ggOweEGLgo2G81DVDMG28wsgyrqy7sTdZbycEnCqIfQKHBftM8hJ
MW7sssmLD1ed0HmAgPIEOgGPlwfHlNRP5wyf4+kQUkm3PgbuE2fuPo7S3ow+HMBio5mn8BNi/FqP
JX6s4EAkt20HFMwNE5tEQCdDi/alYVBdjMMOQcHrcKg4ojA9XRxLglxlUnkpfGmxWA/tt3ErEHag
lMDo707jY2T7faErTL9t+8mjVTCUAfWV2q2SWJD55p0HRto0C5uf3KETBtDmCOtKiJuhegQutFu0
D7uMSCWZ3g9MFSRCQvdEfVSMD/l+j0KyRiLNjTbbkSgliuDmRxASqh2MubRHu2vOr3zKUSu+aDl/
hoMc4iO9wwC+C4Pm+9XFFIkYW50f4yww+w5zHvOsaYYUssyplUfqvXGJQUvvyKZnHVt5wNWPVcYp
X9x4d2bjPQSfyGl6wAczZk9ZUzHAaF7V2oWpj3U5YcPS3tYNEnioimXSgYqzJleDk2Ui28eQk5Dr
oqCIjHSqSxYX0LHG5qVtSoHQAaaQYc46ZiPa9BXyovSAqDLnznlXkagwmeUeXKHiqt+D3IwS2HCt
+isY+8vmiVEH/OuD7GJgkHK+SVozqSjXmBnJ3jOPuYzq8mWjI2VUUtEKt92aSCdqHoZJVP/toGsC
P7V1P7FNv/Ia1kLjLsW9kiMa0+/fUJcYQOscmQ2B7u65Mue3L46FrQqvsVoi0XkmhQgzxuqj42Pf
8B5B8NJR5G8UyeOodgyrutq1pMo7+Haf8sgKkxNKOzl25haKfypJkeiUitLoSO2VpRktjco1ZZdA
AwkmGMIW9gT1mBeh1TZPR+o3t/NKvnLF7ocdQApfllOswDyGOE0QtpyEbPDEEEVJh2FnUpi/i4sw
XMrMEJWoKdBVZxF/+mw/shyKF5EM27d3dEq7HWqQV3eBxHLmO4sfixSBGZgDp8EjNo0xPlSlWZSP
rEa/ia+XD9H5Mln8FR6yL8TS3x89gEqfQuvcJ91De5jRG4xpa7kD0TqPQT1bWziOtlKStI77OcWD
y5ALD8pjMVdX5T+90lDYa7ch0Em7SwXH5T0kcrRFvS0SEHXZzVJZnJ/dXm/NzqAChsto4FTsU9wA
xnGSUTLlxAca2yTQTmxc8oz94my1c4PboPt4vQomwXy/uUGwEI0U33ekNVKcqnTu/QD6Uj6UkiB6
EowUi8kdy2cCTcKOrC7uKFw+xrR/BJ0Lw5jqLEeVgqYPej3tj/2sXsEG6a/BxkMJ1SUVfF4oSOmX
RhTiHYQYuoy3TLYibhXlt5mdPCm53ZGVfVihMvyk3P3L8VmePwJ9roxk3g/F3TyUNQR4Fg/x4tK9
ghXLjoPIVAp4ha5OaBYJqz5AoRyybGEDdQ5b2pcCjjKJ2gPDVC2AKcIb6g7ocJ+zC/nlz4gHQRF8
MU2nOFbLu+1/i5X85AzADhFOZnG/FITlBJlk+6xwPjTWpGHqgPBTKN1E2Jp1/o99ALn5K+S/VG5z
thMyXt/Z+pv+AboInbDjHpvAkLU+CiJby7/cqeVPEezS6Xaa+h/nnyWXKAs5bjTaYIMlnz/iQrRk
iulSO+EGSuzw0+u/80Lt3yv3ca8QJPNa/SoTSZtI6eHR3M0gS/BXpDT969ZAeg5ytiBNICc+1SWI
JN6eZ2BR2l9CQiiss3dfIPGdQr/a6JHmiSbQRaPTnTf+tVnQ6s2FSczpbPcMtOX3L7QJOWgUSaUO
wQWLEJ1FKKPWoq53L2OgC02GjczFcxZhtI01qoH/HlBl7XziCH0DxklSPJAdMpmwqOtfveX8zaWr
jq0140tW7iyuvzAyksdl7QcsubIqP0zlsETn3gGvCZN9wUfxQDB3Qn+iJsDPI0BSPDV59uF8hW7L
x0dTmQAjxlNJwrJ8LdiI4qJZMUvk3x4V46wfVokFv5UlWJZPyFIIJ7CXRAxrTq3CFSrDCFaCK+i4
RN0yAMI0bfb+afsz6cMyKcWN75xAoPl02t+r3c/sudjibFz82lJsXzvh4Qow4w2oWHpCKRCslRg6
VFJN5ZSlfQPjLz34oW2SD+hkWlz/qGqL2uYzoZXxL+7s+/lN5sRpyvTgVWJrCcpWMN0nnJoaBeHy
dL70jIydpbW6Lx4XlHiQhZPBeT1P6poL0ocW7WzdFlBzaR2vdLFCoTr2/IS40J/WGX/doxoVRrPT
oENXHB54LKHnSdn/hFVFnqalmQm7QiFbtfI71HrjHe/yGNrLKr8hM5XEbV6iOgKVNqoVQThdPgBm
wlTVGGcbi9RuHKvK14GWryYDcU3ZJ8kTYPuKfOzahjVHFewe41CgMJj8c9DV+n3wo29sbHVEBHjY
/9hkA//0SUUbm1CF0pCY784cdtgNly78C/FeyPA1WW91w6S3+++4LSh1O5BmOkFWfPPi4w/sGWuH
PPPgrzgMu6qycHzW++0zqxd1zREnxUgnRlsbQYD8mRUtc5ukzCK/1UODyvICXys0V/908rTPI526
phcdYLg9GP2x7b5hiRla2dF+jH5aHMIOYkZygN/21AbvxBQdzuQUuXNs9rHe6vbf5dUufjcqdqNL
q6BFCk4CmfMz8W4y2CvR02F2X9ZRqnSi40C3dnrpWaY24AkhwH+O0wBKlUIIgt01ik6ShgHFEprQ
E77Kmv7mweakL+fIzoTkbPwyASITnv2BGL4N733u9lcuzIjd7wClFFxRql+MPlz1Cr1HdLLghkgo
95yt54ysx2dZLIuLfjTAd57Xf/SuuhSIbAQzAuEv+fbfmJ7uO+Vk4n3x5dDyar3I6kcmd6u2l1Ga
xLg1KxhllLBVQxTUeNkxJjiNAkM444uAtKfcNY0dGyFNohxxOJtQdOi3aKrZHG/wlZLmtCAT4CyK
Mww+KPEGVUko0VvZf3U5S625ZdkmCEqF+2Uy8UUlozCBQkiL4Qm943R7Lvg628o+oeAFAjrbLtBQ
L0/vodD5OgV25j1JbiOAv6zO7pdVNxHJqqcxcFv8RBO8HdUvWPalVeQfVuWUILSVQjXawzTUPyP0
3m9UmCZTdRlr4BgFZRfOMoUpGbwPbXehjmtdyjxnCtGfiFGztmOJauXEbOviczm1oLtHiSkyzDTZ
xY2WQMPZk6fYZPi9rfaftNm446nxeVS/R8AHdoKKA2f/NxUsx2cALqgWHbaaTQf5CRgyRjIDEz1+
cWRCjRFxZ+UCihfXGRCv+mANg3a48CxJQpS0IMtPA7G0Qe+yMeHvEQmKKN9hDHYHI3PRChN2WXD3
8nxNfFZiMetrelZZxEMmJDIUrtDURjqNmo9gCfQ/oyjYTqTXJ7L0H1pir9NKxs1jvueL/glIRgaB
+1/a23RoQxB5BRwfJtdu9366OZNn3hK2tbAlZQMV6bcc1SCB2VPWFv5AW8H+NK4oiLtCW0KG7Q74
vBK8zxgAuVybf2CUKVHhtYx+pP9obbiLEXWsKJrKYFWXM5t2s24hK4QbtDAFl+lzgtEsIhoo3EA+
w35UFueVcq5XuDsDXjKIzgyK0TM4l1MCGsSbq5stNmEtgCAUYGSY9UXrYtI/uhlltfT0LQDexKE9
Qhnn4IX3BCOEqnZleKCkPKBAn8lOlI3nDWjonOdQ9JOEFyPAWCjikpGitEjGxTSi7Smhbnl7NyNp
EvbEY04Pt3FMe1yF7KhZwxso+uq0XsliKF/20up19wtAFxLJAz3jvWPjHPNVwuZvcsfjYpAjRg94
DMsnQ0s/m9DumKXL6Zk7vhcu1Hn+Yxgus2W2LFW2gSAao0YCfWD3vqJQ4KLin3+N2utnX5/gbIuA
q4VPDE4pRN5PSggLS0aNOsfa0AdNlJlttVa4DRkbkVvTukgVeTW582ByPtFt90s5oDnIE3yWa9gV
oQ1HqHpizvcaxpjBkI1/DLugdO3CZz0t79rYWy10EFRqcc+1PqbXtV1mBOuTsLmeeprC1jsTyoUU
sFTD0dD4Y3srISNBUatBb3rDMtAT1Rdmxk/mzZ9XVhPsjPkQpbEOgeNlNsDIQqy7nRAywPE3RCaT
gM03laJoB/xhPn2PzM2U3HHgSNPUCtyqmuL3NdZriWyoueG27O/vLISp8juqaU0EHkQkLSpt6m38
wN6lb5D2cnCIHJUS3SrqW2qurrDZ+rMozmaF2ZIkaI2Q9ZE9nB6a7Zoiq9Nv+aKu1cEb2umRatu1
8FIdbTVVKuUM9AXQ2mjMS/jprxyafE0DHI4LVFYVtnfo0Ped7mlqJBIdUaM3SthNzLyhSvDLddRp
VI68DKAhjkVP3V2YenDkweezd39qOhPtif3ERW5d58tsompaoKzLeDPg06yU1Rrj2mknj7J+e9g7
HUQr5QnQE6C8EsD+QY5KhpKMmi1ujaKIbX60pSc3qHd9XgkYF2vrnPzIZeUZrNAOrcpfPCUJKYJW
PyN+EkIhlVOpzQ00smGvqjC6xF79e3Q459j75Upqwaf85Dnjp89wel6/7/X0rgdqKNaLznY/9zgO
WZ5vyy76YjOXnhFJRLH6tcY5sU4Nh+4Vo5fFBG+4T4KYsmzrRqXSXSXByhzw77VavaBuYtRGQ7tQ
UTCIkL/mLWegnq8P8w6RrsRpndLxyZP2PMLIIpKjUx4dpqjiyONJPNthy+KKu4iSeyKUigeW0LVK
MVoKRZt6G12RccFeKkLSbNLl9epxOg3QJXF4qbgy+in8hwWb5YsSIXvc4ReIXDVqaR9MdNnXnpPO
fUy7ws+LwwVMhni1n/ZuXGG40wVzX8DO6BqFZ1pqj/R9d/W95k3oiyAD+rUWGWgTZSVHTB71F7/9
GB88EoaXCXahjqSnYcJIUbuW/QCMKZASKjKt1aPp74RYqIol2M2J8npBQExCsbukD0Uhmg8Ld+hx
lnc0FUA+ea471615sg4WWDc8tL9LmH65uiO9pvY/9anC/e3htNZGIWadlNm2hKJBbR9exYZsESyP
y1PwrIe3swaiqJES9OS8WZXHmlpMR8+Hjnam0N9AtMxJBwDaPJxAQE+lIcj6fyLSaW52+zHdHigh
iZ/+05W4/IG6k+8Dp5D3pUeinLOgRVDurY7EE7t73DOkDdNwnj4lN1NNTgo0D76guaCN38aw21Ey
UryZ7jzrVTbFvuj0uqJgCWPAawbDnwNtN08jtgtGnXa9pSHJrU0LgAu/e1tPP8blCYdO5cq26gnD
To/0Rz133m2ZQSWWp7yljCuii6JnKqAigjNkMpaVCNZe+OfxLUFB9Q1Hn0jzzGF11bPKi533kAqo
iHzuez76zj2HL9WAoCNNWHwy9qIJGcPjik/ruHp3ObXwbu3QZInzpXGYhDewlnl4ROPsIKVN6ZwV
07kIiPRXamsu2Do+DOLhRoseEA8A+4l3eI69J5GYj/zvmNFQKbGwYjBW7+L1CIi8sQGnNMUsgsRW
xC10fE8xIeUnJ5gO/iiNqxeT0NLdZL0l/IvsO3L7szLO79OGePP9/VGVzBwd6cFQs5ptddgxBrCo
Jva8Xc325GQl18BSF3hQV2pL03du/SXq6m2qUGmIT8s+bHuKd9B8T9mn25XT2tctHka6QD3p2z2T
GJmSkLWhoLgL7FpV3zhfqFaindwB7B1JCNbm9YsMbSil+X2LVmj+VYFsVuXicQs+EB7AJ1i+30bH
iuB7C4Pk/+H2HhDjD2Tu+Fji8fio9jTBc5CxEyf7FeT9Pj2kAZ5kLARy+SXUac810YiykKD1Wqci
S96+QL9aSAmaQPJRdodIHzzjNhWi2l9hKAApYToNwv3VezLGeRxY8JJUBvhPVvg4Bafg2qC5C8IY
UZCoEmAeQB4ziSm7dKzqmWMORq165ef7ude54nfp4CMLb3dTM9DbglqshWRX4naV4cNNOQKx1iaY
EFMZKK9b3CoruBYCHAeirPDW/LvrQHcesbSipgAHWNjWQ0SqYT8/7HcvsIULG6Z8GIWeobyc83x2
K/iojllGWwtZr7Dg5tbmrkKTKDQzcX1kYkZix264QdY3BgO3kELMa7sSxQ/l9oX83gJxSD4hSfYk
ZaHkun8+jacYYASvNqvVu1j6PSKxcuaKJww8g5E5p9AdwbnlcaZJOIvXGUqsSZLeoxmaJaYa98WN
BFWwxUq6jEUYbVWtJH11ITbjk6o8HrqRRodDM7onot57dDM7auaJv28qu9oMXoE44y/v2w/YGvgq
DyXIUEBSxudC8/4XwZ61vKiguTAbP7WLsqJNHyFFESFJkJJ8XU1mY12i2FK8sRTdawOPxTAS7hKB
1gYWkfm/jIhEAqwI/vAqV3KWx8/nErHVJAZh8A3LDpxJDFaAHUAM0Ah06ovk8Zo8Vn4CnQjvN4Py
rnQygx7zUHozsOwr39fHKwU0Tdx4mJkBlwDSsTk1uDbNuJXDqHLQ7VVOMAd5cpYSdnE3gjf1iCIj
1nL/Dax/SMMKYbSexTh4oRktmhKzYOphskVD0d3U4EAttXHgz/Tr8JH0OOvyvVgLh7tC7+kiBamB
Bn5qJyhbtc9xgBuEXqXGiZUMX8wBe+4e1SJMhkjQG2TrP4rpPrSRgkvCOBjMzkUYRPK5j5z0/OFI
Mo1Xl8qkStnLSMY6yWMHEKmNK+vBjVk0BiYhnthaNCLV9+8bqnErPrCCAR8yfl2ibaoraFtYt8B6
OPCbBzjK713MLcxIvvbrwFNxE3saJv7LV5pWB4X+zOWfjoF9ajBLWTXt84N13wOaXqqIdj3jO6Lu
DbdQGYRTmoqvGUNuvz+u8bnJjAPbd5FYOknlV8W5nylhlT0rO3MwNfkunE7qP0T7UTIVc/A0Dk/f
UA2iFs3+F9EK+SpSKqAp6+781Q0ckjkeTdqtl4b/l7xx44RqUDOl4Tcd40gim2LLX0j0Jj+4GnUQ
nkgTEFLGQSTJvkRO15FII3L60DbuVVRafC1Fgh6/epgkhI/k2HRNyfpDu7lHwrWfH7BXBYd8P/Kx
92F9YG6qMg66Bh6VIEjLSMblwDukt8btEf73Y5awTc0I3FYj5S2+JtJY5zP4Koecw7sOL+eanBUe
rl6y5zW3RaygGE5HanTtAPdYnJVpygUc5o26zCnRAlOKsBX8YLgfYTL9o4YENrWGeua6ry4TxnT7
GMF0vDzxQ54U1pVlMQSfnCYrr+HBpXFwkXVhyQth6ehF8mRC+sHdAg9qcZYvS4J0iy62eKWd0h/g
VpnuXkc8hwObrnufh23sGgXHQ7FoFQ0R3GnPCSop1ji9WHcKWtNdIK+cgQePcemsxXC4LFtL2Emh
pmYxwBl+sZbFHmuzdx3zIMztfm0kBdD++BfS3TCtYcU83XzOsIncGI1s+eQwvIRMVCusOip5WHHt
lgS/GCRY0a6a4P8FUPfnuaMEKn8U/rzWj/iYmFfgSox2feEBVMaSyAVHBGDw+3LJXp4MPTQUSODH
F7Rv23dD+bHCU+A/4aXzTkSP87HD4GVaHgT1DQMPP8uc2g0Hd/GHAK1LfqX64gUNVp9mEIgByv9i
KmvaGLwTfXOXS++7dqd6jEbxGowRu+6Gbn8N9ByjNH/ECZEVwhZlehekF7XfOqtSC2JlqO5RT9i1
J0FbMfNGVY9HVVUtAtHo6EoDvOVQmEDdY5IpthTJmYH0+UvBHL2ml7s09cTTUBvwQCoxBw0amsqC
+to3NJeaAEJRZxtou9tPSBgZJzYh9Kr32Bcynevl3TcKY30A2OJSNE2i0RnHtxWdoyO3+ozf3BAg
J3FFAH3OQOA1Dp30O/JyvidygKnkXq/cosOPrN2Gff/uAeXj5qzz3rsn5uk/Ze58CrnvwdFY56Op
W/Fex1A75e4EcCUxOiecJz4trADS32eV7XY7uGBOaXCshQlt8Dy7rxTWMtZcFBvx+oAcg8M9XgPm
BovoljQFAzb3WLZbTGbJcUVuOrUNYW4ePX5Lv7lglN/SKKnUQ6kwaInGQwwLEDToDAUtjPmUV1N9
Bmt/GD0NIhRnHZWcoce7podKWNJT7K3QRxI7wdUcHsTXJQlMLSh/nkcQ1ajMLjvkjs9CfNHxWkfH
8gJIvaBA5UgbXjnf+8vJKEWHqur4qSuMlY4ciohW2aJ2lX7bmaBr/uyJrQCoubzbETZPWGjmeH/r
NHu0YO6Uw05KGzLWu8e1wOCwJRKKp7zXcfw7GwDIABYI0hlIqaWhuIPvdu6xt+vuxCIZm5+dIf7I
wEVUQ7J2dSbB0sgIGh8diSZ2UlNxq2bqRqdSQjny5YBSxsiA6HY5dl1Ogkc6TumvTqtu6sUAwNmQ
feaD0X4e8GYPV2ngcqywXiZargKaEnkfFxG7Wapym917f3vavf4bJohjUAsMGwMHZCmP+hsjMNYP
6dYHDFqDiDFFIVf0GL5wRrCpPY8o7I2TroE4UomjqSzmwW0NW33y6nldIUZRI/uh89gvlCH4v1zo
KVmPsyETPYfBgq2tFM4zagSx0Bwv+rqIyhOQm4KMoawrteCzJjC2CI17EjDjkvgCqBYKhOk7Nem4
17+f6G46YctxRGvYZBmb/zDw3uPVN9BVg1p2A/zudZOG1YA6zv+PRhWdH2BtJSws1hL0Ncc9Pcle
NIF/ps27gsZp0lP4ZjsnbH37qO4CRlRpD86wOrnp8fhm9AkqLxjbQxhkqLAh6Dmz4zGhJU7cXr84
MlTgr8sXabmtNdilbYLBYn/gLxFTVKygVpkRoEPv5T1o/bYgxCuR3+udP5wigmnM//SiAqg6VBBk
jTxst2CNaxakipDIAEImaFVZljb3TbClIvQCGKa3nvzEjcTUwYi83OMd7Oquk9x4eKD3HtZZ7Dnt
tyEyUB2wLCeIhQXyZogtWbLA4n+/2CKr3j8fGZsMM5iT0CAHHgczZpSg6zzZ8YE48HhqFwC/sIlO
JRPusDmiVjcSTFfxpznHdZuflX5A0ByIhN9UbsdELOBYGmkCeqdoFCWD2kbYFMqtUxMmbRyRc0HF
0HkVTUkgyXwuVpX5vnGHfwXu99BN1KVoDIIbTvNejFZZgrrpUYBC6m26HXA+jlY7wEtIPtEgXyab
YCdD9ZZKKmBHQp1xf0SSJDGxNBoiEXSI8HLAETicAJKDASDhSMJi4il1R4dMhQ9exy+fBgMjOvcD
CEhBVeCbOSeDwpLhpRIQn7NEVRojitGNpGeNb0DDw1I/X0i0zxXGl6JoIq9RsNw+SMM9O1CsrTUX
MboJaFDp8YPFQYLigu7+kH38De5wBUolIqUdimafWPx50PDdQHeyR2YRsPAXWQRM+t1FB1yV+BjK
5sKdWD4YIbHeUPiOFDPMfiVGcDtxxcubrJqo5jdYncPRQyV4gnfSBahDGT/D5U0Z2UL524OuWqnG
xfMcr1Kkv3Uo3do+gT52dhV9qkJG6UosYNj8L9jurC14krUlqGYH8uD3+ERqQe5r5DEf9MLiblcS
mdi58cvnv1RSPX/bYss+FNkRepBM7+9AMAYfI6LXUMHavgOQR2mEtVyluDMqu7T2qDJ+2IcFFQej
w/Q7BxJPcokz72NMVyhYtLVxEV1gnf/L/b0IwVwrKkNVfxHG3wcSqVR7uaNvIXe3QbhxYWD/c28A
kukzjes+QHByxJmTXBYLvR7X0hj/61so06vK4j6luu4SE4zWGyTH/hDALBYjb1HtkGEjobT9u0GZ
Qz849hiTtHKt4VQDA+BwcDBM0hDP/NCQ+9X2FcyGsx4cv25RueEUD2Q3/mNNalT/vNxWNFGGrxqo
GaikGVszIG2HGoo9mrEWd7gfJYGWj9qerxAa6n2CM4Vkl9v9MXSBEJrJKEyGPHa51O72TSVeBPdw
JfqsC8EbDZYxaw67ZNbA1GU/GDTy5toWn1dl7svD8qj7UjyiKlZeDb4Kxbv1RweG5mq95t9iALYZ
6vRHlbTzEsrv0Az2GT368bSidb3grpvKPCAQs8OC51h39PjE4/mvJNnW/NepNNeLrfVJXSZDVeut
znGZuHDNqG77TrSFJa7TKkR9hoTmOflDVdi2axn7mmRo/zXa+54S8pgzAH9CesdvGFyYAY5A6Z9x
Un1nRpuy45osrniAqFAQNSCg3YMwu3UY7F+OsWBwHXFQVk98u/ARU/TqucinNB6DRjv3jHZPxXUJ
JcioIIXuwPSy+d/YafJ9hOvo7AE0XYnMMnsRSaIyRDuxCSm9LX4XBuuFx+FWONpT1+sn074J2/oS
mJQz5GHaR6pLMuKIu7R1pW6G8TtFgHtdIQ/Yk3JGIA4KpgXoq7ZIxJbXYqmZPId1oYJSvSt4myVh
L0Cpg9uoNOD8HvO+2MPMJXy8L0DgCWrPMnl+H/q9oFa+5+RaQ9ziIXFzIqriWt5zKMpelSvEiNVB
1zXfaF3s8aT8DNnHi8UpZAv+lJ04p49pMb671g/6AW/ylJhFel+NOJNtieFqIryWxXHGCcZkjMaQ
jdKFgvTqIBDfqxE+Vwbdlgn/jyTxi5/X0/RYbT4LSGiNxIE2EEnusGeVa+xFVBvUaLpEdwoc3ds6
Kn9zQQCeMBwbm6IIHeH+k9YXY635hx8l2AEZVNmnxABMu3DVO7Cv2RMgeeVzt3dmFe0PmtBUBARB
0P/TvLJTLwIhLT/HJ1unScOT0WyidMg5Jl79LhjuHCR45PUP0kQ1qWylaRpacpd+/9/JsZ19Dto4
wlsIkMMjc7jpwi3vSNnvOpBdA0OCC2neIJmw4+XgNxX2EcojUef3oMmhGeLaBrxcAqudagLoDaPC
MB6MylUuJ0ap6tFmSX53shwjnmZg9HOm8l6JHYW3bspKLPIXTgxz6CYrxyIlpkXwfPfmEohXC2ue
tBVmdtENLIz+HWf7lBKiUqBfx/uAqmCflU+1iVeKfnvnjHoVYK1Rq3hriBFZCevRviYvNWyW68CR
AKEFN9IFqbkERRRerxXnE5A9+MdzfFP4ZQnCiX8PszoVZDKx/kHxPGozDTEmIvaOTZx9O8HqX0fk
IvAWAdh6cUSbNmdrq4vVT4XyhIf3Qa4nocRLlUzn3cd7dchWFsEjd5F20jTfBKhqFp/jOTCzmg+B
ZAEo46yiRZkpzdtbWbjhYyxXuqcqUyntgDUNTm8udMotd4L9G+4SzVsKjTO9mxzw4PwlmT7gJmMp
gMEopkMwbQY4otxOIwiSOBT3wUc/eE+BDVu+tQxuhQ3CxuhJ+lfB5PrT3aQN9FcNeJO10xKxi2Kx
QZB1kGZN0GfH9TUHKaF2XI6evBlJgKz6MhbErjyesrDLHFdHUnKxSeGCPHZNnfsTsDwfdrMOagUn
UMlwrhSvTvnHrkVjv7O1KLcd+x45Tq022ldYdx70KRPLsSpCeAgOFyoQp1v0nNzBghwCbkUki1XA
whp0swv8+FWJuMgEp+9Yv6OuK/CP9Ha4YmtoU8RfalauQOp8e5IhJgowyeLcoju9DDMgE+oxSkFa
u9/tL3wyM9CUzuY3mGu0jIzq+sTSrky3xjepu0zNRsiuk77IfHpm/T12ky7wK3I7mHCDKEvj5ZPi
FtUf9hSzszVHLDIHiWcWEPGuPk71V2Md1s9LJqp1mHB/Scj1n4LbjtrboqIQbqoeM8/8FnbVTsOk
I5qzjrzQVQ5tQJV1tQaLHlCB+Oqcle8SuF4MMoTR7R65numcZSdBmOG+0Lugq7LWo+skJ9l59VFg
za/ntWuzt14eN7gjP9vjMEVrbLm8m/JetEMVZ0Mi6ksjX0KqsRaYeCA9MNr7IyqC8Q/8PdJVQs6S
OXsb32kk0570uOQ4tS5T2lhNRUDLEh3nvZcqhhWZRY9tQC4r4WpugW51p4XJ2LQx270OpnCNLKks
G0MQU5L1zxkzuUV3+y6i5w0zZT/PVY/dhpnQnJkMIF0dm3sYlp/UYFBf+NqmUFG8er1v1XcNUKfh
aARMcTYC/MAEj9nJYqHGb/tMRInsXD2KqlHd4x0j2IE5V/JIbrjpD9fPMB5RNG4zAbZxdGSJdL0t
6WgwSbQ2TT0ga9kg4ltDaH3v+0yvISXJ0PFoEQbjxvhI8euejIpZVdzWC5/5tJkB+cNTohQg/xig
SgY70/fXHcGtFsic4Gskra1gh1wys8k1yT+XO78C3a1P0pVy8FKR3FhoydXRql+Bv21DUS9b8hHQ
AXuyGMdgiDEdIYEm7/C2ZDp3BuGuEj8G8FZFZ5a4zLLtEjZlKfsRXnqMc0MRxnH3vPR8xv/6aLej
a32QDg7nzrTFX/KBAAWtQZG9L/wkm+lnTqlke6sXjCL4VcxeJSay0PmgG1RIKVFR7tlQCKW7p3dt
llqqYnGPxa1NpIkAt4/6h9xlWIM5U06/3D+db1pwIIf9f1VSdJ7fNOkK+4GGjJz+Bhyb627HBmjj
z2siXhVUF1IRaBCKqGcIZzC5tGs+uNF7faZffLrxKhegkctnAAo8BU00aLBKp0TSLLnqdl2cN+9Y
KUnWlhZWYlGSnbVfzVGCHbjayxtrQ/7hbsSFluljopBTyO+31/+sF0HoexemLVQnrEarbQ9ZiVM5
vVuCjZlDSaJXiLipf4flhhvTte4tDFA+ccU5T+fuFLibnPyBZuzxrPkQO9yqLntHt23TStDe9LKO
izGk+5lVirGCJynv99VPo4o7gHltSDY146sjzk9h4upTm7Fp/InUPvb6BpYHxmy4ZPDmVC+gZh0S
xy7yQbwTOI2rt1hvnKN0tu3YwXvxVHS1B8r4oTfVCSkLHOIWygKgJZNa9pyfWmheWvhE0IeaVpkh
QSU4LxhjP+PIJxvPkhjyHjlJ8gBm5WzPQ/7/ljhswe1hsI59MpzZMakxd2LabMr6yZIDVDnV3n9Y
ouQC2MBLXNCb9VadKxE0CH15ih4xjy4En7MD6b3enNOSZDyBhjM0iQA4UFymtK6d0xShN9mV/tM1
Xt5h4vT6tHirMtTXns2WdFoNZjwV2DT6hKUpy7QLak0KnssismyMipdFt9XFSqGLuFWsxqICmxkR
fYNJT8YpNW3GNc8sN5X8jt+NmPD3ltmlLhBwwBuGUqkGDV9917FWHM/CopFh8qujmTutknFwNuMZ
HshWL7GJokM+aD3dfWbtpffxZ/PTvPL36jkxftBRpffemWkD4objbxBw3EFKNSe1glygS1R2/bu7
hTbjmo0BGNUA2/oFgQvossj0y+5EVmEtGFJMwFJTmDy8mAHSedBPLVaeoWkSHP8ucFwaqKEc1iAc
OJf8gyKQoG5N7ZHyMGDBcrNbzLyxs2GeyChww2hogd9uq4VR4G/oYN5XGlPH9S3Sl7s7y7vNUDmT
R8QkZjFPxCxbo//pYXlg4WzMm2oTCUmAuF5e5s7SB6JEikeDntGp+PcHnu2qpu2wQIMq1bjdUdXj
+g3QQq3YHcKioJ6AtjsZYdFWnI+RPJkdnH/VDpc6qCYmrdnnOp1JaeYzjI42Z+Tor79d25KCUb5D
WV1VfqgkZpojM6Jp3Khk8q2lgbaxf5SXqnTrq2FBh1TDYp0ySbiNb2K8lslHAJN38CGwTv4SOak/
dpZrkx3mdvKdQM9kZmzKfXZcgELsJR8gj6WszoIT1LRjDrp/WTDUObYO4rzS+4AUBmFiKar9t+si
7VdN3U32dCaNZLzlvQlHWn4F5eolGiNB2QF20hihyvaWTQO0HZr6XKCEfZMLK+X32J4jLVGnKvtr
jBrm3Zo8iDBOWXT1V1/in3SAkpOPyFEFcWc2WsiOqkbwHeSSc+VOejsjm5wAsStWbsWZZjcGNgtu
Sy5r3Y5DoFJzhCriRLIRoFPm5cEzcHC9+H5nsnVrR14orNvgDLPw6W7x2I+dzaP5NSTo1covFhqs
I/KbDeBjY8nE028XSkC4kyxD+98f53TSf+1/yhRWO2ysjnfsBpZz0RuWrSjemJBY/SVzK7NCius5
qKYMx2MeaJD26sxUep76zYuHVZjBDGuOP3aCutLiXyK2cIp5KzTX9NMHamrs5htQwB94x2EfNKH9
UrONQ1eDqt1PKHmJ+dxY6ffGMvux7j/msL6WE/04iS/PkX8ET8LASNrK2fhS8FIUCmJPe/So9nlh
Tom8puIYcvUVEhtbL9fT7LV1F2tXFcHMC3qZNwUaG+0qhnIYdlsspHU89r7L3rO41N5JmIFMJJY1
JScOi1JQSafuyHyxCthgdE1YFlVR+tHgMDyxdIkI/S1006vgE7rzuSvhJPZ8l2Qv8NdEq3wyKhlF
EWQAJS/4NOSgs3jJ3hgcrH5AEH5qJ5T0aRsn4g6MndQD0okUbEQB2ns4g09UhEEMz6XwewA3f66a
GT7PqghQ8tNKxwYe6uBcpAmUbiYRkspjRskUd97ddGM1NLxJP/xuq+Udf4d+eudZLEEDKOwp5aWf
LkvBLHLuqafeYCysUq6RhYn7SZ5w3s7ltOVqr8sqK3L7tFQqKaOHxoZIhCsiD3QyUMaDDGwodxYA
U9qaC0hQ1E4gBKb1TjPaDww5xTFuWc5EbtXQKLL2IRGehjMQIY4g5nwPoQvYAyEeFfW4HPVzYkr8
5OURGaKURq8PtfvRZhwpSs0vXjZHUa6q/DBoPFZRt89Ag88n2HVp1Psu/HSa6OPJO54pW9xAHLxC
vfdoswfq9cBUcfXroi1i0Le2/svRJ4ba73sTVuMIAIO7GVSEDHuTxe1WqgBloiol9m+1mmEzcXyc
ciuo+wqYu4TX3MWgT8GcKsjtr07t0qHI4kU7VMs8vONOerWgsN+Gb2/6LpPXyPnJQ66K0ue6LepX
0/SQWmWIiFf6UqIsGDkJi+RMX2nrgw2N4MQh2nB2lQx8vhfvQD7oCw7s4QsLLft9iETKHeAKENP3
+tzK1P+mBTMfYRiYTHAtuPytrZFkRsD6x80wpMoQ6RgTk7BS3eXTjED66DV0ee+PhnYymiDimEUn
maB7kEkkz9t/Oq4WwIF6ckoRApB7zm0XFK6O7nF0yIANCtSLJVRwQLd/+HEjG3XOKTOdg+t3wqmt
0ntIfzbBgFY1y4VfvTiRfi2cFJnB+GGMy5iyJv8q2coFt+TUIvUjmOKimwGZNp/sHZi1N9KbLuxT
WsF9tJB1KLUTYasRIeF/970mUKLucdcTRj1YUfcfem3T3abC2m5MFRbTAjtGkEOreG+vYD3pG8NK
jcLdgq2G7uVQlIDQGEKmdFcX0C6MbTQXX0zeeeD+sfTuF4HR/0mlrDfaZPooNf571XOAJynmVIKv
XcnAuGI4Y3N4sG8kNsa1nJjaZHg17vtEfIS9R/YEFizIOJxt4Yy83xiBcMIRBHPsvnQtVhhO0ZKh
qvCf1wcXtmtQXDLqbF5RFB45DF/914WR9Bksc5MgcuYtaaUwaZWG27NV2/ngS5wH1BZlL8E4c0nu
wAvO32AItBw3wE5pXwnFe7L1Kgd6wshdhceNFli5EaFkGym14PfpeaZzBmc+Ll9h9E7CM0Etxm3Z
AZrlSZ93E+YSBU3f009v4swSOOQHjZBorwsbl/hjCQesK6IhPN83yS/xren+raCLdUZEuDFbjElI
e3wxHBXIaZucZ4ZRch9UVexD29mcX5+KmewAmLvxlqo4MCXhZI+HR3QWI+ifN0ggrCbg3kLNdcSC
01lfN2iB7g1L/bbN2WjEV7EuDxIvEInmIoFohG5iW6tUp7oNmstlzJvxqBEDT2GIW9xGqEbeS9XB
WMDEbaMgRVQPi862a0NTpJWSgWpLML1FraW0s9strDzTcw7Pr9aHhfJKoqrnmq5Vl5JHC2iqoPm+
mAXNIReF3+FxS6dp/qilm3Jk5SPYqDUuMAF1InXrhpznWrTtJv0pzWWeRr3gisw8YK2ATzrm5M7a
0algHqO28MC7BxGT0j4hVQcDJZpYZX3KcploOsdojZrIJutvlVekMXCORPMZLn+ZZktHIsUF6QUG
5IUSTRsPdlrHyvSfc42RzEEomKhZYJuniP8ZHellOsPiwwrHEwXBFShOj49cWI9Irxg6AT7K5PUv
9U+W8NK9nnafGk3UAiHdADJ03Mx2ZwGx6D3IVHUhWtfBqnzW1Tru05GxiZSY0nCzB6wMCK5xWzTI
GWUQd0qccWvzh+zfQDyXbSCVeNocXCVmIMy0o9Gf93ntczGiHpfMDR2wailUVw0qgcL0S0+4Ircq
+KDMd7zWn+Q9AmHIrC54uqCKLKW2ZklBVDbIEz37zPuspgpGcOtNs7rhC88MHb3IQRycIl7tc152
1RuwHnZvHfKm8zS0qiYUJAt0XC8EGgYEJq4fANnVFjv1Gew19DE+G1zCk4vAe3vPyU+pEnvO4UjQ
KdxaHi3JlL1Z+a4E/V0tpm+A60G1rGwxY1jyPSysmydlTXzl+S5n4IPpKUGOgp1VZz/rXhrhywio
mXBqI4u0D4nNTzbwco+3oMUmLBuSMXgU6brH8TEiKpaWapjKVaNMlrvzXQjYL+8X4kNMMieYXkCu
HH5i4pRjzYxwOFWch4Vr3zwOQX25jcHqfeMXkwLSGRAN5mMpJx1kW4bcExQWOjCoMt1aACdPfpZW
UWRILKbe0e+IAxJ3Xm6zi8+geiejXlQoF4p0twn1G0r6k82u10WmT9IAH2W+RH5GbDKd1SVCCafO
K7grWcZeAji1bXSe0QEr1sZX9ufYRRx46vL/j5H5xsPYY8Z2DBNjhIYwSFoXr6MBEf7NA3T7Jo2O
uXqNZEcsDGKDluSuWd5OPdPnfb/DLpzmsObj0GhQnfHbKojMYtua23GGMOKSm/ZplOJT+NekgefP
8XdYBDjbH4LqKjI8bZ1Z3CPkelk8aKGu8TJ28yQEk1aOi8P7tapQ8q4RbXlB5B2UsABwfXoC990f
h8uzyd/WsneRQYirX+qDywno8A3Z3CcI3ztCwOw8Q2Gmfh8duldmqMYAqL43kC5cSckTeCtiIAyH
Y4wEbdT2SviPkH+SprpLX89mhuAv1Fegf0245TPobm1RfIwNKiDrfz1O2l/vHdtonmuK6I1J+wfm
toESXHoE5D9UEjx9PqqSqkNhiSRnoa249tqmZJTdGw9c/6x2WY1fLKbtoz4yaZpvt88Qwuyo3EnF
BI+iTERW2+OWNto17c/rrJFSvjOkbaY70GuVr6Dis+SLkWG/t9FaYIA/492ulBWKoyIXDDRwBay2
73tDL20qz1n5DCtULmD0/AOnsJCFj0Dp3Df8yiTDzXhA0LxLygN/mVZpvHumItmDTsIG0GO70n9A
gXs0qE13LHFpw1UrnI7rnvcrg8aduy5JPg3L//bTkYf54rI1jC3cmTTGFOQr4DJxly+DyEGKqmF+
Thndr9xoVaH7oUTUen1iwrdJnEdiVNzUrMrwZ3Ohk3rUq9l6ffGxytSVpqItmLDO/Yy8ZRVeMqnp
VuizKkNWA10RoqjnGornbIyArNN1eDIZRxJEtFAEGLfyi39QS3cEhtqKqw/DoUzRTgBFYeV3RASo
FlhZyTWvuC+sL/QSLTHCfErYp0hkboNQ+adjWPx04tYnEzqv/njftjnmSMPATSDP4Yy9mmrYKfKt
7yb4buobbE1sYZBFJt2RqHZU2k9opkveuu/1CBZvBONZ3y8/uRlAWBismWQV+kO3Xx3WSgp+vQQf
Vcbbimf2/PA2hCY3Veah18bCThT+6Il5mIBdLq6viLWWhfkewJs/1MAr6PYwI2sdTz64kIobNf9T
MyyJnLWFHSCp/QM3vaPuPOkFCQ6IiAaeF+fcq+DfSZDhDrsrqJY+mSMMhtzdwHBP9CWuCq7uiEgT
/JFuAD/x3E+hfb/SMSzaac1NjZ7doUSMFGKPZUI6TIqltE2c657NT6bAvvIs/fowxVZgbs2uv1k5
FdGn8S+ej97PxOtksjiOfYNtKYC5bYGJapmL3DthxxC9TkUv0qm9HnGdKAXMqi5p0YAgLVzSYDJP
RHM7hb5/nbFF394kl/VPAoygCQLeZYM+bVFWE9tqDdF5iVSAJaGnJeSPcbI/HqgZJAd3Dewzw5IB
W46cUWAksn6UlMR8/Pk/vYG2YiNKTpP/QqTFqZF/0Df51fQAu5BZG0LKFIb/ZLQv8NSY5HsVGq9R
B5bhNvtkZmSM4dBx+x7tCSZGZv+SaaYmRtBuHNTmNYs7xj35zYot8d3UTwpKuOI0yA8IPHHWwnon
zqilxV+KqCzSAY4/eoHYsojuelNrWDHKiHtthNZ3kXk/cvxpd2RcVZOWxGIrvfi3J0mzy4+ucVm3
bv4sWXP8TksTavAEZSArO+nJe0IxTw0Tajtn3bpyNyOZXIx1Nld2cer4Zi8yXRdOcBHk8HYk7hIn
5GN0Q7AwWXjKWQ1I61ePNq/BJprFAQ5aX29kFo1W30G2sFEX2kke3buPZrsSduw3whzek1HgLpey
w+AROZXjPdlXqvl09DJAnGrykOvKrBtRfAAzirf57tzzp9nVp8004z9DiG+Y187TNtjFwq23gbkw
lUbazTyDKms9NALELFhSfdubCJLDCRtxDaadljsbtSusIvbkTqytyjuR3d5tSMkPtK8FyllTqtZd
GlL6k0RbuGCqPSGJbY0cEqwDx0kczHynNGumOBL/glpA0UIsVggUhmXzJ8aPxdHEI4F9s4sB3++Q
wT50TKRGglQgPAX4PWy7JKElkJXgYoFL7AOQZrAqjrPLJZPDTeSDheIKn+QWQ/MBzLv3b6vDKi5k
TMtlPgQ8QLXPayOHbQxl1mhQ675Q0GX1688/Co4kBFzHCxkp/OLFTUwBf3UhbP9b8TdcFvPSlnIu
K20hFeRyIQFuUpVzW2YnPIFSZgivJnvaInegCpJ3P+9QfyLFfQfV1xHx0zhxD74WlaIeVZj4VlP+
qfQC0SaAGzrJLj263ETUYEctgzYVBZBaxh0J8oJG7bhTiipmqXLGEO4aX0S05lVmF48byLM/z+vv
m5BhyMsIYTkKGh00q7F5uN1EB8muDZNFK22nJpYNu7gfzYZcxo9yVlQwZ6oqaYjw/3eY3GdtJf4W
ER19KrO3sL2WVvxy8HVlItWTL0pX9FkllqfE/1UlyyZcMphy8ixnuXMlDKdkxIfkgEIGdGdUVfNs
R48Df9e5koFriVhTn1OWNQBib0Ndw8RYBv+3/x157PFJc5ib7aZPJnHUUCfKJ0zfJkIDm3dfDoJY
xq33/OV+PMf/FxDdQF0DKV72v8PTiTgl/DCwzCe5WgUn80bCo1m5tzBVdgOVeWY9JyhPChbbvuV5
TRSRtjfo9yGhna+gHFIm2n1jLKvuQr3EJCnq5fO7yeVYuw/P40pNpXVsE95UeKPBQZeEI7Dk7eSo
toIto+mxoAT414RlFQTplfxdzF8X7gOJlJAIXwcc3nE+m7Tko4uLZ3pQIN+sGlB2lkanad1k4V8o
yGDlB2NpmUSB9kFPPD/XhBaU4+j31GD7BMRKTC6Xi/rurzpLWwkezobXgV7wGPcQfJxfaMJUI7SB
kgFlh4YI64weeqlINEGIfF09ggHfwyEsmw/KhkcwGjWjBUXt+Ajzuo6zj5a8cqnUppPEzQvDkp0S
A9jfd8BJBgKE85gAxGTXIfq3d81bRZWAcC/LF45w3Cl8Av4FUf2U0W/JO+9YHqKDdtYAkuJo4+Hg
YJAY9iOqa3pD08EWl3CrHnlUrkDEjczQ909P+1Z6qVNs4CtBWBNaBb4kUtI1G0d+tJm+4uq7jASn
wCvyXNclt9NKjotDPySBrAQTVi0R1fU7xD/qO3uhS+CWkforuW6V9oYU4Ecbfdmzr6xA0ORuEOmu
4kMfZ70v3VM+yt/BB+7ANIreo+2zT+tNs5fN2SVsGutFuJy24QNj+AGcwTMvnUj9sFpb8MEVt067
6eX8yuOF24ScyUZFACFJ7Bjmkp1hq/MUYSsKTSZa3o3KuTBSjZafPLapJDpgFP+pz0/7DU8FuINb
xBN8aINbImQTU+p5lsNFsAvHD4OMItlvaAlhyoWohOH/jT14HFoKl8KOR5uFqt29ZBbOEf46PwoI
DBwXqq1qU09fDaq5sAXDcR8Lrev2XkFMz7XnFdojuVfMY1+IVvzKplLlHNZmitQN/UGHmDvU1JeP
3zitGojMX4KWfTwXYCSRHXYKhlq0F2g6LleAviWlU3CodGiAdJ79SmMTM/NRzbIDWtysPlvsasb5
AtsT2715WIdjf5ErHWgGREKqIsUWQwKSpBtRzURKyor9p4vbskRyri1OhrTRLrPS85DQXgLikVpq
YKOkC60QUT7GuX5FiXrY/tKCimFsolfO+ZU1hdaM5S097IAjmS53CGXK6zAjik2Soc6QIhagLk1D
C19Y/eNAVP8K0QJmaQX+haSOrpAfF/Co/yEAX2KHYelGiDC6PgJ/fy5mV7COz3I9YzVKpToTbNHi
JcMia4b1n+zx26o6xz3WW14vLOuUxuBJv7RqFjgry/80mvpZ5xrX+HKDe8OfcdxFdyKjBTQXgtkG
Pcqj/AjM5wLGtz7Bz3v43Xbfbg4sElEFnUJjIiBtp6a/S68Jr2/0jNkh1Svg1uotGvZSiCbzvAL1
AwazUEyBveWywqtqLkspjuQhcUgk8H6vNkwCIiLrfQG9cEufSNQu5YyK/InPcyO6Gfneprlfrc1Q
c8bcssUwG00AA60qR8pkWJU0CtCz8MJHU+YqnG0b2kNj6B5k7X6hTDSOt+bythouEqE2aHdZ8sAY
9aKihxsXz9L6wfj0YyDStmWt+mkWRk+O8trcTna5AazCeYkd/7wdfLWUjAy6cCzGDTFxb6Gjlnjj
AMRvUHHphycVGNRGlz5xGlZkWNzCbyALsNScgE5buWaq7yT2fZzO40mwNo7THNjeIGgwaAkS+fQw
WVCu7FYaZQEfutq83P9j3iW9BPUnIKT1vl3fqK4ueYvFKk7hcshum/sWk28a9kMwKAVnnHSOV+IS
YPeo98vfsXWTDU9gjAEzemGu0pcNm+xKGKFp4G4A/ewms6OcffRzL5KFeLgdsRERm/L8RHBX1ViN
2zvj9rxPsPXreR2NdPX3jruJYCz8rP36H0amJUsO2Gu8SWQA9S0Yeoj90wz9zJ79t5FXlKboqsEj
4VZfeIyM5dGNwbUiFqXIzOvF6b4B7OxBKX0EwIDFtonW/K0+0GOlQQGFbjTZBEfE6RkikKVLlKLJ
lXcH5lqUBazvM0Bk4G1QvHE5pKpNLK6XolssvkTkW6kPeETA0Zd1HLBaoJmyXQnSYxfMp13WVDEE
mDDSlA55CKXp3oeRvgpFOks5fYcKdy6jPrl9x/9Wvs0gh/2esenL9G1IW5Xj0/PQzks1+jwl43MX
Tgjdl3rJ6sBXjwkTv+750u9pR/14QmbRVelwXO1c1Qka9h/9SWDzO2XNdgOSR/XjzW3mso1/ztVD
1lUJihuL1eAmQ8a2zaB98sTXXLjogBPHYNsm5wjHHMLcD2icto93V0TP1sP997qdOXUyZ8KSx4Pr
2Atx1oSN+eQYkFgVA7wCj7HY2PshvuSGKaVihf84xiZwZuYtqc9B/9pVDedLm9G3Sr7+C5VX3O3H
FIEYcW8P0k/VKBf56Xtrf7V5QDCjiyMVlJfKa843pbZI3ejVzN03ieeoJ2Iu88Wxe9Ad/MTmTX/F
EJLLm/R+7XoQrpUeuNeVUUGsH1KCRAjZ5GuKb6UDjfhBhy+8WAbMepS0FBMo95yMxY/VgLJucZSK
fjRcgH471N173FgA+UA0AvIOTxiryLpVQF6Btiz3Q0X2T/f9s2KW2y7pgLqdmNmYEwZG/t5JVRVS
YrUVsYK1thC9RNvjv54zSPcz9GLBGdQyWHeKpgzEGCFt0mIa0w6ekY8nR8qdNrKFQk9F6t8BiaQo
l3zJCVjQA2j+l7tvTHiFin0RJtvny/y3Je2x2tbLHF9nl3Z64USoi8TwazHbw1zx57UaNzjUjoeF
GF5Ljkn4bTD06ltdynvJhCqXvLl2JTAHwKprqwKkAuGlK2Hek5y2xJENtF90rzsiTYdUNXjICC0k
Qjp7GCXiSRFc/xlY7aCUAxz7Sx2nuzJ8NJgnX8igM8BKj21uJjI4pcYNwv5IluEn61FJbUO0pbfa
hKx5beLLMFYXdBZ/E6I443jlxH2OPkm0OHXm77tl+HQtL6ZXswtlrMiLq+TVylaYiD3NkFnRIRaI
wDzHdVzwVsvI9nj7FJBq72yp/OHOkFww5nIJp0V1N8053bdPhn1RbCLdYu3GVeLH0wRtseqlpVhg
rWQE75H25a9w02GKH+qOpy2964gPFzg+kx1lA92lifFTiNyOpFdkemJAZvK8myPT2vsls7TPNiK3
/7NQU21enz7wgE0Fhu9cYSxKScU0v5EYhn06unTzwdk4U+GcDJA1AHFWyUfGeuPG4pk9a/Xsz/Ro
sgyPqv5/ZNiVAr/9ZqLbYrQkYInI/tXHb1ejtcO2rhi4KMRyaHnhEPIYrlfa0K8c0i7JYvZTuNn+
UUoNGh88JmnUsYBK07xb98GZN+Luua53dpCwadlpd0ELVJzTQneYZ3Ry+1VeTzIPcOnXOi7xJb4n
WfmA1LvMeI1VhsqjbRqihE8az35QUAoSlneXvkjAR5TN43QtWwWs9uBBO2oFzz1h13QrdMSzOEgi
oRTpNjiVS3//jYfxP/iGPoSzg83SwG46jxhSF4u9IkXCwjigZatqviWWODQasGeGJq+4ooMFjel7
6/ALwnV6tjW5MTEPXuvVzbqct3+e/TSq+uWykanJ51lvSy6dfum9S3k4BJm8VqTAwFckH6+HJSfu
HLUfsTMNmqhfyhMDnhQPPpkHngUAI18fr+2xVUKLYWrk4bWhxh/Dqn5oU58xUbxumUKOskU942Vi
8Vbkoca4K0OyDBoias4BeY+HOKD2nguOISoK+akm4+4eIlAdWqFk+pl4Zs7kPNG21MenTJhpDxI2
XrhS+HaIhK2AYjH4eKjCSE6xzr3fdDdNMHaRSZHeGk5br7AaZjXvacx8mNGhtJDt89WUeNn3TGs+
sT4jq4uxdY6LDYdt2Du5dJHCNgDYU2vEcOHlRR85DZcMhWxxZUX7LTWE8KpomK3Jb/NSdW1CddTc
Y8/JlnaQaZ4ypvPiRE3Otz5zJbK8KF5nFt0os1BegTEp4hpyRQhH4LUxefYiOmmWUNIgT+Odyl2a
/9THa32GMX6MVDMOL4uPHm0oVzLMejIfRalNjw2zYHR4tAhB8lzLdjPYxyhWJt/EoMrkFHes8vjK
m324zE9CugTxPKYTOkiJJQdrJwFYlATMkBy4pGCa0x/9WyIv4fUlrN6zLVW5KnBqUcF6CS5WfPh5
kCiaKpK/MoAq4cYLjy7AwJy7FTx+T7ZtCWN/EMXTXCwoqipedipTnbysNRyMEfLsTqVELPpA5eDR
/iJQ6u+/zEYrOFkgpPuUy/WmFMcbQ7nu8ekSa6bfd6IV/FKyNsiHMvNH3kAYf0O2q+AKYtkeHze2
QuNur0AluXaQnnHezw8cSrsoM5iwBLY0m9KYKM3C3HWHhrO/vDhTrt7GIn2wJZzJFDnBINcvVwAp
gIBGdUETcV2/RQSN29NyNWyiNAHPsTH3Tiwx96xCGnCL4Cz0+5JTDP00zsGkgYkqJ7DgG9hhKIZI
6ITcaAnU7NfBWusXFYWLks4mVePQmXOJQI4YfoRrCevYVIunvp6gnJWn+CkhI8/e7AarFNkuz70d
/N9jOu4WmmFSDVs617yIsI/OENGNOAbW6bn1jlW6rGt2p2sFjMWO3Cp9oDQZLaNM5gbuDPvpuPry
l+Ut/ypQQ5/OvoJYdcOEzQSh+oYK+i+UVI3/quhCCUhveaVQp+iOv8p5pkgocJO6WSkP6S4jm6D2
BJtkELXMmwScXl3Duxn0WlorbLhH5YgrTAOvlaveg6x1sMONnZ5cQ9pCc3Pg0C4zeaXGs73+xpcA
13O1XEJ/cvwl+MLuc6mSKbF6E7/5efbRNxRaq62JbH0mANtbvbT3JbqEHUQPGGs+7sRA2g70QzoV
B6M1u3nCzHdmm86GlEYxgJ23sO935Z4opZl6GwvEYMJ7wAVFph6wrt74m05x5ZRku+NbU6QP5cr0
BzFpfIf+EI/oKjzupKFOnsVc51WH+d9IH84m0NydByUyFZ2BweYkLoGfH/YnuoYjCaHWzyyPX6yP
4GKjv5tM5q7ybQB5PrjN9s0WoHSXi//r3kuQpVVIYQlJnBRTPZZKq2/SKzZrH452dKHf2NPabLtx
kvAKvOXlNlswkar2gBnZh4UGf52uWnG1n0LvvWqAYvDhuIL2EeA7jWgR+ligLEOuzYlIo3UExOnj
BAIdaQaTq/oZeXsigmhVvYL//Fld76X10F0it+Nlo0f566HivzfhElOCg6E8MIR46RFN6gr80j2q
1I1XrsCO1j9fSPN484G7JkxGSa3wvFTWjPKvobkIoFPavRL1EZd7ZRc3PLj0lNlh8m8oF6tob5o6
+8v4j/wtUL88wklfqU1sD4eVgnCuouFeKMe5ysHJgEESL/PvvK1OXyr7owkF1d8jEIETfbvaoBN1
xJuDhL+hfTGy837br3oYW5tsN0kts1j4wONb2U0DCVFiioZhJnWeswefJLu0f73cVbij0X2q1j2v
/doqzl+A9zm/5MWgay9PwAd3j+Tc//vdmsUXK5hi8or/YevDZ3kgNkZZWxq2bSOnGRRRz5kFV2B7
DTo57GKx34SuaSaQGiT2wO9bEtxcJhnjWjiEOUK0U94UyCWfh4n6nRQuUeQij293jBFYG6MB/9xS
0I4GBzTzDF8H0yFFQwzdRwzErJTooYG0MFlNNNEEyazcY4/C2qF3c2Zu+JhIWn0y16Hibns1EJ8x
gvNpjfCYqWIqSZfnaWApRPc0ut8csLJQcta7mYpKtQRYS9ExRMVX0NNkdWZceG7lNJIkodmTuajw
o2Qsa9nEqFieq9fUJIdhikgsn+fgig+99xvuXYBLJ04pHrS7ZCERXmXE/zLlsGL0PwtBkiPDSC73
xEboy8KDftxWO2kveDkaRIrES/E0JM5MGdhiXVZbzDB0ys6QK1hEyu7VU/vviMIau6/rn4q5xmTC
WDbSSjzapBp0ACTfL71wl/aphSdKHrhA7UwNQ0e5BnmeUITlodufhXR4192ewNhnJ3FUGUIC8vtW
kXQXwxhOwLDqEMY5rC51wMphHM9qBcsHQPKzGr7/zCuy9FFXgZjs66O4aVXu0DIq/gGko5wBPxUP
iQOVxr6HrnQIWONGC6rG7GQI9rXdDkIMHblN9GHgwtIKbQWeKcGRgpU08C6h28bFXFtBEyLdeN8Z
nFbCoaKd2gDX4IUw10nviKSCIxNUZZwnDIO5ZF4KTezwJODYWnqVNiUIOwAPFYPNHWAFtYpc2T4S
AjlBWZo9lXUWU+lE3/0KQTCeT5d4oYhaOZhxpY7rU5oCfSpQ8ph/GTfLoC8/59tnpFyOJ1d48qkN
4cEtlSjKbM1NZXp/NT1wLNamSDPgofXiLmTAC8ofYJdfy+yQ6vH4j0QvfL/1qa2t0b+J5cmWR0yU
1aBO2CxIn1fLcgZa0SN+2QibSdu1QiCP9DrAG7KB8g4MQGBQORkj7zDvZlydDWQoeI3zpLdMu/1h
c/dLxt2AKbcGg9DyLBdpkxlgCCN4uvI4E6lgD2pm0fsgzkLJYrtMDgFlDklRThD41kuGX5hm55iC
MIs+ONTIzNXZntom6QSueCQ06g8/UGR6xVWSEIcdzmaMfBMBRDTx9pctc8mJc0ss08avvdJ1wItk
69KnSIVNV/Wf31s3prI1UKCMGy8Fg+PM/gxeJ6Yhcut657lH3Fo5w0BRtojpsD99dgcMUnmfCfOU
Q6Z1Wp0yeJKlmLghKsNGUX3Yh/97xU69i+Nb/z7DJPOrZ1PLoDfXFl8q77OM2MVIm4xgjrXFDLhO
f6QGs5uhp8ebxc+rz4kKd6vkSklxzlo9iwIP2eIWn6Wc6ij4HWsq+Yr/Z7NtWHJu6Iwkw4nzwyHK
XAT9RLFsl7PA9mHvi1J8TrNTDivoolMoNrMFvjVNDPS3Rxl9UWNxHKkjI3GfhY5wbnNV4k29sA5n
46q+JFnj1GttZkWh881LEKAoFQMeRU5TtE+IouSSn8Ba4qe7oh6WoYp6bayhqGNTQYTae6bvFWF6
NceE2AR+XNBRfhNFbjRBwPtoEHxm5/SWjCd+IiarXYo1U5mm+HE6C7v5Z/Jnuzt4l0ljVFrJgawd
wJPHDy+XwIkAsvqKE6XFFucQEkMU9yvDXJxiNEzeA7D/InlUSIKI5uSxNViy8pHTYJiAxd9ZHMgI
7r91QAZEjyiYqI/ivsYUQMDf+pg196G+3M4SpT0EWcVAwOPNKtVx07QwX5+Co6CkZXkzZQad+tCl
7g733liyfUJgipNo2jrjD66ejbDGLwQ5Ex0KFOprB6DfuxNu2d5c7E6sGH2Idgj5aeAFnJSq/B1U
ZCqLeIw+dQluAqzswDHFnwfYA0EeRDnXlbS8EtqQTPiSjAI4Og4+bO+h0aAk2Knf094N1lrnvHKl
vICdP5sWoanvbUx61fE+wZUFyu1cfGE+jKLxd3f9IiQbIKgMDxZdY2H3ndI27xGHtdIMO4OPnBZA
D26r+aQPPbbZ7VczeNsE7CwfBqlOlEiI97PsVruq9JYHmg0Mf7j79+35CBo8Xfoc05+JSesn1FeK
tPf2pufoYjViJkyP9UiEeDT4aLjF8qUpr2ZopqHqqZYi4HLO2y0hD8y8EOWfeMCftN8kxmzohL+q
WL9fg72yGwaCRXubSDUYtY6AfTikmCh1TI8HUdYck6X+vIfyF1fso9CItPdu2TdgEWHspUxgLGGt
HyP3SIwCfdBomvggV4mmJKOQfjObPiZmAC0Z4hArWdrSK2blD9662+NFa9ekztzAayb0aHf4B+hs
Bxl4kQjORkEJHpEN3a7h31y0ZxZkZBuAvoHrvlD8Ul0j2GdH3osmtvSiPYMHeZ61R4sGtIb2B1gJ
dEzfLT9WAFWwFZc069VhG/nO9DOZavKMrihtI7m2m54tueDZtAgzwjKGWuYB2CW7KAkpmcNuzYhJ
gKX2Agnmd1ggPwEdbC5GEXPm9pVXcOUgGU8A93MnQPQeVhL2bzGE2SPsrT2So1t7GBj6ummlwnLr
0EhslYYS7RuGS6uI/8G6LZ/tW00ERScKWq9STCplPUUVzKSzerhH8Ro92erOpnFAu0QctggqhIdh
Zzv2mTOopTLUqOZCfc/dIxKZYjGRM7/lLNAWZvgeKhnrxENZhFeLMbMdyY9fwL0kHYfWRBKPmWpX
/Rn8TjvhNS3JXjpl/RwWsQOWYvrOe/f6DKxFTJDnVhVxGMCKDW6dGt5gSF/v8+7zkW6nLr59JJj+
/9zjgDyXjqtLbcNQMM0Xko+n/AzEEYZS+yJ7et0FPKe4Wo0jOgCHWLhJ+JERQtyUIzs0Q3H3yq/g
W7OvWVbyRSCRCpEsHZFm2W3rQ2Z0QexuVkoyPwnW9S42WL16HnnfQlkn7f3OseHNwuKF8aSFMbNE
83kSDO/hpCZci28E4sU4zaBO7ON2LMFJjbb8v/XVkvWPxpk8pApaLJ+JU3ULVCcNHu41J0ucPpVh
//L3i445WLgS3d5rVtajLKhY5ndgBW11nqoRzdh3Q0nIOJXOC3SBZJHP35LzH0l9BXLjE+lx/eOc
xf5ZDDst6amLDcdziScVXPBS5fDtnLApPs/2mB+lTf1oQMOFQo4s8YX4mJsj3txuEBIFvwK/W2PR
fmupg0qNwS9zSpq8vcH/rBHHgZ0N9oOERGklytnzl3zCKz3x4oSXqtlxwKd3WdTJvYKodms0ofmn
z/nbAwHwpBjJSW1tn7K9/5qQcdNTZkItfWoZI+dsOsLhTZMp0Hx0pLoCZ48U7wVQOXGDpWQnCWGs
W6cCyMjX0BuRoOAcGXHtnj6nmX+ndYLpVd5BqEjylxHeig4/p9076y88K710COVgcX9g6YfTkAHh
3ZGvVQAQscN1fMlOIDHGsTnBFZAKBA4FuK/hYatMhLFcM75THDi2UCA1pRA1Ol+ArvR8yA5omPAV
cUajMKMtU9OTKewhHpHibCIcdcOGx8oeFI54MjXxNpYu6xhUhE5qtbWFJfBAVkjqzCZlErWeFD/b
uspLX3IgB2v9ktvCZQrlukvfeRBs4F/yQ5ls7fioYaJjlKGc3R3RAxvaaSo7TzqNcxQ276Z1eOnP
szY4Ite1ovmm62vCR2g0wy02pAVgFJpZftahx7gAcpiX7g0FIxcQV596UHqsl592A28Q3ZTwSmvo
ItdkhHm2Dm6hUjso3qM44m8yDU1cg/8Z/mJOPqQgDOp7CJ7DHcfwj/1AEhQMYNrsU1g60b7KGe0a
UJspUd6naYkCckot9//F7zPW4UWiMirhYSDXByaF+PxUcnX0nXJno8YvCW2phJIcqsbwYKvEldUr
3krtEOneWY4hng12GchkKIpjNnV+y4542hBtTHJ9W/KPd/gYNGCSwJN6xQHXL8wZvkdmSDtbsIS2
S3xp/+k9paM8p5LkvDRqkdQCiSIzC3H+5xLzqJMbz6P3epy4Jal/FxcUQ7TP8BnpCLauU/LRDXUX
8hK+FKhM1gziVXS7K+2lCcEJrqhZc++pmibCRN7A5irMiOuvQu9Ee9T50hok4UORNcfCjnRuuQ0r
h7tfED/dg4GFK9CRuTisgcwK35zuuBFgs/wQh90yp1dQ/Mdw2tq0ATOZPWKGGxAsZZwGH7edt53/
XVXUBy+A5Frw1S/psJThqS6atRXuqaCI8lxHMGt4Bl4M+PQZA7R0LckHERs+IZ1kizmnrf6p6kxv
/YdPtyjFSBHnPtFTIcsDEosidICURVg5Trwh/PXIzhDsqS6FoSH9P51UH5QBPjuh/LBemjtaFu32
ulIHW9bK8N/SFcl4gAe5cnokXUjL7DoZsQMbdy13HGsNnVSh3TZqNFlKzmsZ+mGTzYaocbGgD4S4
A5VDzERWHqABi8bX0UARPFPUO76Vk8ZvLhirl2Kw7XuXRsCTdRgMQAJOFnyiMflQjqz2cQCAh5nC
SUA6tR8Q5tmqAllDqKI7hBrZOobCWvN4fIY1b16WS2rHuAfghJeKyNSwtHGniN+w/q4NGsDJaViK
jF+FIQcFxQzBb0Cv6eNeMH92v55k6vjXDM5mBbfG1h+UebtX7ZpYlo4JMuJ9QKp2uhpZgqH1X4IQ
uTAz7AQju/Vv2CKi+oU/vsXiu1M4qQFVPyYsxBvRrUBr9a5eCxilxcwcsnb8fITt6+MZa5RPDXRl
kDSwhrXO+db+l+Kzlz0MypKGWqMEw3poXrlbIFQtjyLZpgE24G5NLY+kErIpw2esLJl2seeHM8vg
IRIsUzBhlIyZ7OTftPaOFv86OfjDUT3vQGONF+5Ylj6IcJXaMJ1UGoZWo6WUupN3Ti+Cl/28g5od
P1WA6cf5YHxhYRR2MYuaH+V3Bfda+ESpdnk/CnXOqmzB7ZSoiy5+WyBOAl2VFUECcUqd2iHQzKg1
Nc5VfzNl/jprP1flusXERgvS+O6A4qbgCr6J0YlLddJN/9mKz+1kg5uOq2EBqR5kZ3ou/nNtoteF
gdZwFzIbHguBRbsgEMClfcsEn5Vxh5USsbMffkR9G1b/Co1UuZH+A5ZafS/zyKatE8JA6FjBqSOb
qaeb11eI30X718efu4nTsAcTMFz7Eo3KBUURwx/ga7BxwdWiNopWYfpG2EfqxwidZTd2hVxQZoX1
+mwDxM1HfUL+nP7y4Nm4MG+covzW/0Uk9Fw9cFs9yuHJEbvmDQryUEFml5Ws0IoR+iAWPFNP1/wi
UoAMl4pNpYNs6jybU7PEnBWNFBebI/XCvDByt06yOaRSkcbotWf1dNe18L5CJd1vuqxqWDaRHzAx
tygihqZ0aV74giDnOedr7a8ynK00IK/YbXkw0NcB8E5OCRku8ueHGno0l/45dhxewEl7th82wWtN
76dC3aOJgLOiK2akCGb4qIzAysNcPP9YoPWihKRja5LMGYzIlQ8LSykZJ3vR1f1CYjG2AInobu+l
b7pgMB+gcf3yRZMvHSILskqJSvVosyWz0fPddxoCsVlqQXRlMpQ+LNRVP2ZsxwEXNlRhlF+1adoI
NyOqtsbzZQBH6FiWIQ+fREtw7HrEZCTUluoZk87U2fgqEnZeBIVJAq4us0+Nd9GBsiTZ4tr9R0YZ
cvM5+FIMNga+VJQf8A2TOSfc6U+j9GmDVj3rtwc0IY+2EArtODicPD9atIwJqoG8J1ViXDr1vblL
lpNRkGnYwPV0ieiInNMenHuBLeBuv5mpSRkcz+zeiIUds0Squtw52GtRbxZywx1oCGbMoq85SbTA
3WC0OTt/ehescjecByoGjxBzuTPnGvZZu6JQmbb9LH8iI18zmP/lSx3lzQfp2if+L6pIvcrUq3Io
lNq7SfVf+ui/951m09ea2Wu+tQszJuuUn48h6BLbPxdkyqqC3flFsVeAyS4Kf3T7WwLA0p3ZmeA6
8OBQUZwPoAleuqeT+LhZVbEyqkEK+o5BTFeJZOUnEbhVWcAosM4gK2H+7o4cUwl5ZCiU8PJxrBSC
EC1kGy5gXu2LLApsj0hvCGRrKcu+t7ZKTEEPpwrzMHc8toWW689GQ75hYF0x/m/OZoLT08MVO2Bz
c+Ag0CVFb13rT2qfClG6sEkxxJvh5dpAMZ78CZlMN9fY6dwII0NAoArbK8dRuqTA0Qj4/nu1DRnp
7gHwxw63ri3M6p+UlO/t6aUDYi6pNRHIgtAkyYxsU+aZxEwPmgTOTO5VkQ0pXbEqQuCTiZtjOpfx
Sc5NU5uBqAlJlUyYBUv1SGs9cHlPDunW9iYjJ6aBUwzpodUj8WF+K7iOR3XZI23Gdo4m4Nq/S7VN
1OzRypRJqAjnyUevwulSePrqh3U4iekIVTOwIYyK74VEP6EMlsGtSfQHqdu0pGnQQk/5U6//o/RD
5gSNuZ6PBkt6MeHxcrU6x7oGySVDf00g6f3iU6XfdbpvgNenesfqaUqEHzWwhYGYB6xi2qpQ9G5j
YMtVTl75yDgAH1/0VNIoDAocUI5596F+yytNQtBlD/he/+ePswQRtFNHBxwDat+K+56m+rCKe+0/
pGRSznb13viDCpUmlJ47G6s2QGcoj+YmfPYxryZ2yLCdrMG9lC2S0SMzGWuKS3xSXbnvAxO5UJJr
IwYoTujwVgXeIvWrjA80F+3Pzb0IrHgnp1vvcR0uBzbb0BMHUv/VyAe5EEmQ3o5BrCloYDXfDDnK
HFSUdmQvaXMnltuy2WNhxWR3Itgp0rIOTcsOcBOjRS5Y8YF9w1fuEuiGPF4wkFw0kN6JaADuHTD7
Y4VWn3nOrJ7O39r/LeKIEjjbt7zRuW9HhvHSOkjoliRnxkQ4tDMoAAx03zHJI47KDrPFNZXiHvR0
07yNsXPk8SCcYtmMLmYdljGw84f4ciRRveTCShLuL1cDFKYFd/SHhvQhp+MHOI/GC6t0IzfTOmld
03yNOakah/B/7qo/A74IoVFBK1AYourOFxG1BGFGOXZAUZFPX/8XgjZyWjIXm3w32cDb1pf8a622
IB9XEYogfZqoQQaI2eYicuf315Lb7soQHdqLBFaXYifZ1WKMo4Y3giGE6P/ocDWV1kPHiGiOtj6V
9EdsM9jUrohvyqgVIv/+H8jt96T+Y/L8X02BTou5ktnZ9Emq1VpNUXEs6GO5o4fAffvUB81Dckx2
L312kpWeMhh6vrDzXEU5IzrRiSzUmHoKNiVp/6G7QEpcnlTxmNiJ9s/77hyNYtPFtWEqImZZdbr/
vOVwHHfG9cKwCiqgP9W/lJjesGBBgtI9taQod8wipn1DwGieT7vI/JJClWQGXB1RQblUgbStaXGB
wyjCH0EaUow4HMNNhNFzrOjnGW32gpAQW5is/Ds6ekwBYoq7rFa0i4kXoTy8E1ghOViRzgmgT2iy
dy5DhP4xt1OkhaWrgCJAv737lBonXyNkB1BVdIDay/ozm+3+eVLT2eUTbJot11UVvShNtO/2t5DS
3+tC0nU+ejc49NrBxN64umMleIQrRMyC5wBlkQWeQJUn7jHgFww4NwqSlXeHbv5Ok2GXppZBNWau
9/Bya5btIYWxzQ4PuUOqUmt4/t0W1pjgG60fXBoKA7CXZWQbK9t2Zv4pqqOE9yxGzJxSTjySXeZE
sKEeUuv5f8+PQyFsl6Hm6ParmU6TzpxoyVBtBB6wX8u5+aPpaXQPLRfPoyzJCRb4KjhJHk4HZ05Z
NC7aoFkw+RMCtTes3MSOh5NrIgx8N5mp/mlc3O7cHN+1ElN6dW/JdtABnXNZ+ofMtFzY/0j/FWjE
Z4+hB1ehneHLAIhqFWJGOU7UVuKF+QhpwXKjlrnD9BpprqHW+5RkS7nR92xRMgtpF2R0Yv1aSZa+
FTbAND+dRbtPy3+pmEE9+d8ykerrd5W6+fhJ3U0mACr/+YWqgnMgs4dlVidXRtD80oG4hi6JtMCF
/e4XpuSjGPpdm4FtpWPusaGru1nnNh8kElmADGCcmbPThsogneD8aJOn3NDiMMrUfTUPOTxNNT2u
Ytb4bjCjPNhZAm0/+7R80rLNvrn/A82Vp6jiw5JOrOJPZBY1b/JxRRm9vMsTehYdXTnK8ylgXxWC
8o4aHsNLbcZHsHhPL9q9BPZKnN2HV0qQ/4yLhgHnDlbf6suNS2FDnlEd2GNMtG9fAlsW5RjPnOP6
gXYUdZMJj+TSilfMqu+g03vOkWaLjCdY4lgRwUFNpSlAeTme5QAcVq0uT3YAcLYd1EN8py1A8Cym
i5iwK4cIqyvGbYamQSaiscFnMkKMeByf0o+uTAIHSNC04prVYYVD0MjWD3OTSuThqvP2guFC84aL
bF5atePHORBuUdx0cz07qpDRksV/EBQszo9moWKSxUmcUgCrSigRxNnbEZ3y2BHSoUrTpl/j61tC
Vk59mPVhw5UKlwhPN9iX91/QtszRH1djR/LCHe/UIJQozwYhDG6uMKpKHFux/Nh6+IGjZMnN8KVN
gaVJ1Tunc7YNLnG7ntIYSe3/NtXWNriWiTVnTJQ+mx1hxFgz1t2uPgrteVeigVNYi+tbD6Yl8J3T
jD2nnE/cDSsgtQygcUWZRNPxhYKySPIyocuR0Dwaf4hORqAYaJ50+rIk4rZjjaEHdGS7gklpw5vh
yg+uAx1ACVM3SZtW8FhDIbGTVnZsgFl5P58ojumhWaByVF0oCza9qK4HxElXys1//Jiy0ksZo0Qy
Rx1c27hOxrHjStvb/TUozNcOOwvl5cModYeOERqq8s6QkQAGNjIGItRL2ccL3hdlXun1pAHfzyJy
D6iRtoL1qky4GpKFIGICw1W0+UEuc91l10+T13iXsmLzEmcAyeRpsvNPUX7Xbm2eq8wlUWkv5xRb
TmKqnALuxo017mEe8aEQ0ZnG+vmneEGBxIxgV2IgeEcb7f/gv/gdcI4sIDtwvTM7yvc+pIc5wpgu
OJYs/UnaqL26goLhcJ8uno4OtEk/5Hr8bX6ORRCYEtjU/yeCDG7XDBNcuLkrN724BONtAa0Vfn47
PZMe/rgO5b0HAV14X6GCxzpuBS/IaL8WJoVv2hkOKIZKUhUH1scbz2BewLAuR5G4ZRwau5qsRSpc
MEEzaEa+HJco1ZyjgZTVWtGQNRmu4hc1eECw+C9yKHYBnfJNYivYu8m8eEkiGk2XTGB9ni3GpJKG
r5xIdTFZXxMT6W1CZPM5MJmCh5H/VtfKdm3UWUjcsIx6j9Pil0pIlhSo9Xel3RmaHBDtKt8FktBE
hosfxvtgWBTCMO6JDz0jcRpjp05P1ZZ1yDL0C4XVg/c7dAD+7V7VohZTr8wUuzE8/pAplA57WpM9
+BIfYjEpCqLrQCsS38DMy6LNKi4uV4euxgf4erfWcl4Fs/JTA9yMz8brZqrmrUCEIy57fdSNhnLW
aMqSbX7SuVMLyZhzgzB6+hjDTu9ELuL2A0Vwevt8vL16CYfbvP4s1g31KrDFhZiNsu9pMR4BOQGP
+tygPocDIKZ/qoo0aWGspQ9OuuQ6ue1mu/NO9Va/4uCWBnE6czHFDBdOtG8HLPzHJYDvuJDqgXWq
hIVDvFkyEjH1SKjyK97jjsFNsWhRx7APJ1D24BruP6cF7EY8JLQGK+Wi7l/xLfGbeJaEFY9vgOR0
ucZV5+ru8gxsS4SuSYP7UEC7YugBe4NvbpI9vOTM32R7J1AmLlzOTxWIoZXripfY2CAF1kYe+HXT
XHpoaVay/3dwbdbYtV/qZzZPReYMlnxv1VHIZwctOVbm5ypIdTwJROXrxtTjCK8zVdUm6fmbLluo
V/CSc7ZixSkcpRMN3UIpL+J3YmBQQ9N6tiqfLc2MN+AOQ6auq+VIwW38aJsoWvycO4WLtITt8ZRo
B6bJuHDUo//69tHmNRdL556bhH/MG5StK5CPyD8AucfjX2/UCYoqzyTjbV6L9+/ueRTLnXRFK7Za
z2pTMrOan4l1NZMQ8nEqNBhlSvPCoNKdaj0CgOxXiKgwcAscmLstbPjU5ei61Ld0akLHjRYDKSMl
++dMmcFfY/rx7+f1ye9L0gk3x6a5tyozvtbpgCifqgZXzeyW4tSy6dWW32BZqvXbcf+4o5qn/kra
i2gScLSx/dW3H+TLhavAh7GFie1d1SMG5zPvof9BVKZ66+6WaCbLq69veYNpAwtaxAPQ252B2YP+
tg0g+nT6GdyJnhmKYJMxMBZVzl5Lb4FfvCe9CQ1mt/YpQGrp7H+euf+PnnXdEW3H2DsNBGJhC5Gf
Ct93g80AMW7Ao43tjZLQJnkrajtPWHVlkO44PbFm7YTzdHGQZc8QGy5r4GTcuHgqfLuoXo2cryTl
rZ9Zrqy22vQvB21qIxkvziKzeCSCBj8iGgxyR6+KWNqJYOyp5wPd23HPC4Abq2400lSYEUPVRrjW
fr4MwpbV+XyOYhP/7hItcpP83tB1F60ku+f3semjQpR/+9rd0AOlHa5r3Sm3IpSpHz1vEextggOs
TumhaZii3gt8/EO/IRKsLmWLobNo0JPq0kEqzdc72RukT9H6yqwEzDMtUCn7meBvDyFS2mGB2boX
Vm1DCXZ5WW5tjRRcilmhaggGCMxnE+7DhELGr3/VhkBRgQnlGdPLX/CQEl7PzQekYBaVZfbD+9bF
CB6miX9DmGHUefSq0+zy0UnwStnS82MrhEuVtc9J6MOBpbPkTFqytpjHN2gcI61UqQtvm/T3+pNV
Mmpy2Mw8pAoblHYK5Fpxdci6eL3A8Bg6d9vF1YlkYPAD3nAWqMeXO4I7JKKayGpgM+WhOh2TRJwm
bJ2S8pWxmqmnM9KVp2NMnznPBoPli3zQAGm88IyDI7vNgNhiFXsBWmcoyFTk0iYB+sZATpdJEBPn
gX1FYflacJa1NzPODYfL8HLEQrGD1p40lAWq+DDc9GA+Q7/C5ccw51aRviwgWzfZqbSZjRG55Mu3
u5qbwsGD8zogjjKlG+UFmQ69N5v56EEDW3bGJvTsF94DgSotxWVdalyTVLIbiBnmiBonsF2e5yiS
fIO879Y0ojqQpjVVrDdLgHJTN4aaYtYEC0Emq63fqb93qmdcZzyet6zInFTyEQy+FpXUfBBfkC4K
yiR0vqaRSWmDEokZjCtg4/MLSuDcQYFj2ZCqjtsRCjxuUJGfU1vEzUH83s/pWfEBHypVSLtqaYM2
w9rVrEjbeoUc/ut4mr7KqM3OGIBI9uJujgNftrbuZ/9ti3iXAGLUNZiQLdet54xyJcaMWUHMc7di
5m2gVQv4o4Q0Ugdikh9uwHI4wIhsBRyTs13fCL2w+BPes/daE/36t7k2mReBK7xNkm7zoqb1cFvL
xBOjEXRakOjZphS62mYoVFg9BMdXRqq84XXQDY5NWrzRyqmBUae/YVrXj9pqg0wAhJo8/SUpCYdG
FmW/YJ0SxB2NVeI1qFuDUOAwD0dnOg80ZLDtqGa/M+Eu2Gl7ghDZtIxEWvz/kdONxg5ahJB4XODM
BweUj6odYt/GH/fb4FQaFDVBWP2dtwT+dDOAF6YDoUQVkq7IPAyPLqS5vfcwPMr+CUM5F/HxAxhI
NVRP0m330hrct5eDP0nrbGqfDQzTBdEkJ7ESOEGkF/EZePBA+kwYllrOQcIVUhE4KuCpcf9b2Seo
sFA/GK3WkG+/mxhAiMmmxpq9DG2Z4wXHFsflJz7SCDjTXPUlvkZL8l+n0nfVsJix/4l0McBQHDlc
GjpsUJnEuV2M4WLG3lZlsJVAeqrlTDBV4FSwckflNoBo1cD6nB237XFgV7ZOG9mrtilcmE8nc3wo
4s2p7528EcScOzf4+onj7QUcE/zWuo8O4BJBXgzVdR0gNOvdr9pwhsgw9AeI19A05vXFMs9RyOj2
lpdpA8pJCA3suePmJMDVg3hq9DxHKU/+fI6/5h6PQG3FnZUSy74EZV1wzrnNcFURBq8PPGC4AzfO
xL5xRNro+YS3Nde/a5R/PtHkkKKKAZyUsl22yWgi1c1pYvPyZQHHA82+krS+wFq6Fhbi+XuYPSHj
yy44XUK7Y78huKhTx6nR5IpJGuDVOX3R3hIeEyFMyvLPo0k3UO337Pg7SnWwd5uYvSN29fvIkAOS
SIuFZaZ02pe5NSEuOkcd8JNmN/5Ms9EbNq6PiWuse3dBARLoS3cBV+2quyU7V2YTW8v9Yj6wF/J1
YwKYuCY4/MtHlpN7CHjETCslv/yrqWuyxH2tzbR/4T+txvB3csslnbB62UW2MZBA8uySrdw/swAO
WTtqZ5x3NDtu6WK8TgN9foanlPtDWlcIpASvSixoBgxKaWPuQgSGSt190QA0nPqD8IXM5h50ltuq
YJTD5Q691Pj4QFaYixHBEZvKP+l6XCsi8Mth1d1JIX+MBI+7rRDL5s72ebQ1rY/xbtijfsO3DU/u
gKdRfMf9MV9ZP39vUm/skUkU9jcoEwqo/5eXDNHMJPvyOfOd1oDhFgjIEpEIO1H8yFX15ugOUnA9
aLlAAfXDJYmMzlLdJHuxjN4iWSDpIID2zCSsBtDwNKliwZ8jed/pmBq7qioo+SIcFTVkyhnNv4Bw
iBzfOD3d+kmXPLeuPdNC/a6IkGYAzYS23MUozZmIS18LEltAJKc2n6Il27vnluTwi2xykctoXaOk
N7mH1NUVtHMKDAw00uoakQ3RDBryeopCxAG9ogWGq4a+1AP1Fq9C8BX8fvmk5Ljtj3YfY7ktWswp
sK1jyPWjezURa9aU+Y9nnioseptsZSinfCXezhEOc++CC6KZSYaWb4zl2T1qtPYDJ3nhmKBtCm2V
KshKAZh5aC9VcgeylsiGaINcDRdCnGGakfoM7Me6EKOBH3jUDuaZZaD2c36waei76/d0i9gEQxWP
xPt3wdA3eXW2A61BKS9kLGUep/r1ogiwakpPaHmr+r0q8bBNumsD3eLIXHSu5917ZqdswI97e2BZ
Ug4dj7V63mgergKnAZinxrCHIuyH7VlyQvhA+3pz/sTnEzSGzaSq727YEta1CkKwxqbxWI02edgI
V71dLNofcaFWP1M3iOJvM4FEwc2PPW8Q1J6ZcHlPAdjfO+cPUx0PKsquzLHIjgrSJlU1cQcV0loj
TV/jfn87xwAf1/8pzzcSHa2wocfd5CPbORYnPiB9UnFSFCRd/6HqM63o7ZAZw4ztY77evHiyaOmW
CjPfRGZUezSDqxDxTHlJnRRKZDI493Ql+rTbSKdBWRXojX/TOUl/DHejU7ZyhMRmMzrBNw4sedTF
ANaG6Urgmc0OpdpORbSP0ZPF8rbfMEubwHfKQEqqPPR40d3BzljliJiH98YgCkEjRhTbKxAl05uc
6d+Xh9QwpzNTeuVgb85TD97Czdks0tSHVM9tAbtHvBBiBFVy5D/CY3FiFpb/3a1lDZRdHbfFZ6RO
p0PwAU6Pq/h3dV6Qgy3/ZtvoyhLz/UXXhDoOJ0htiLAnck9SOWqBZDp7HEb4Iff2kyqOCDPqD3Px
7ZpRmtjRjDl3aknJxmf/vkj7RbDxcvMHhtXj4iIAVW9YgIZnxEjD2y1lyzWFGeDTvpCZvEY9CtG4
g99fLC/yMKYRVnUyqGKv4//56WRWcVWi3dJMj9Rnb+UTysK/PTZWAu1TC5gqQ6QancPghA30b66w
CTLiqTE/V/mjtOMYHk61PgPw/da+sKAz7ziIYHlVxc6ffngcSpWRq5zUVvLCPwl/QK+BDRNB3/qO
MiWofx6UkztMcLWbJdHY4Fs6aQJ0uo4SHhiE9Xx6LUFHuXHIuiJKn6IptDBq1aQYsws9MobbhlyN
G4/AITAQLvNzJMqrESPUtcYc3++XzxB3TC6GCETVhALjueCd/ECkn46/yLrQfIKaNojJwsQvq+ZZ
KsvwG15U8XaW1TcdfG+fMvofOz5QtcNXHemw1bvpVqWqUxtRD/gNI7X09dlKzLYpfR5tPTIYTKiZ
qTc7ShzmbyOcdrmhX9SN+R8TWzuyWhhRsJFADWBVOV7N6kFsCrASj04AiFQBOuIXjH7cKDZSuYu5
73GIQOJm5iv6xnb0oZ/zaj/xp2aBnXdoAApy2lftj3VZ0mByoKDPSLjV3xSYW6Nh8ywW35WKmyyI
X29bMZsLSsn96jS/jbH3wJuWXCuV+o3vwS4A+GG7lBmFCubdQL9uELlfh5BHB01rTTOOoUVx1cLJ
Lc1XMroDigQ81+ZNHOf+5t1wUIvxOVpsHKpcNtkf2bbBKsdKLIKJ94tpqZ/+FDDKtdt8kEBw/jpN
2TmlaIRYJS/HSNcnW73sUWpkkCehZdPAgFDWBoxMiYCPq0ZIew1aMh4OfRMOjFGtlLxUJF1ybzwJ
BifbbJDTRAzmSmN8LY6zPE61JlXYuuQvYdwzUlkzQiJ8YVBqENUBkdH3yd82hpt3u3rkEWfi0C14
i91NevXTxldXDyXVJk8vTXeR92JEhNRLINzbHALrLKoH6XhwRhjrGrc5gApvDWhs/dsKhyqsGdi6
Yx1pEs3UM0TVYZFg2BpxUTOmef1GFKB5GjbWbyRoz4Bh2+a3hj1Lxis3NVakwZi5JVnnbpX4609J
hMZWXtyme3mJyrq8vu8duAIdauC6cVW1F1SHeSvFtxDwUtPBvPG7brfFxBPHDkmkYwcrclONvOOS
hB0OI8+dzkLPxhS4+k+NKXMCG8LteUU55a3mkwAEk53IpATM6obwzK/c5assM9DL76xO4xWqjnAj
gNThJHoO2Ws2xF0e4d4ttt7FRb1MKWjKsFO3wUw44lCToub2Omq4OuvCeve8264a/HXhgYOxCOgl
Vl8q3kHyBoxr152gY+goVGFpJF+GxdBGiIdH+syYhouDkoAwMAHW3O7D7qh3x4dvLI4bnIgaTbe1
ZDJSVHtDS4zQ1X1+9QjdJjGny2LRxMerw/j/TGQaEF4eqdobet+BTmFKSwl5kLsvkVAMoXLQ5sU8
lOhdr/e+27DhXbl65PX8H0A3z2wBXhGQvvNruw1fLd4h2FWtvVBZfrZsxVmdPPyjwGBhlr4HwFSU
BdYa8gev2YBOVXH3cspkBp+BNhJs4BQBJegz6CKeFdFliGRF6P/5hiuY2pLbPtLHq/2GPamgTp8e
g30MHWb+8FMPJSVduAfqYfjHpFy5DSPXSQZxUib/S+7Xnhcz1FhMWYKUy8WbXuCGTKi5aIy9KCFe
HoNaI/6hknIwsmjNIcdmv2u6srFCMHwvsYRVXQs3cZ/C6hAjWlmHb3nZe8NVQo9yPrfUprLUroiR
AmNPiWX1VKqiwWnM7s2dmBkI0PTfZuLeYgktQp9Qm2qzaYn1B5pXdBJQjpLUW8JW6gIYLl5vu2pE
2Pc2V4qkOEW/1ouMHh3k5dQzcTWNMB7SJwyzrIPCFs37wZRk2JME+xVMQtY2MFemL7clpFL9LyjQ
zV8JOTcjM9osdFoobyf/NQA6MQ+1o85xbhfM3pFHrjlB3UY5m5jC9m9FzRPF5cJiygEoyDPmF9hR
RCeFujsIgjOAJ9aWEYuZvISmKrj6OihLgvWvgBObxRQz8k4eBia+9KIR6osyCBN2CWThIjEq64en
BbX2vgL9DizW7O3FD45ZvG8pwa1tpJX4bi7Vzs1N9yk3DoSgT3srAJOX1TAqALVxeBPwZCIynDBs
zClAPj4Zwk57teCxZDa/GT72mJfu0X4Hrl6O8sYrWBx18zuWFPSjy/PvT3tC8so4xNTm5UUgIlaZ
eTi7u28EUGuHMj9XB2olo9Hzb0bB4AoVcjMIWNtVDRFj8BfeDo6eUVb/s0Z3hjfOi0Cg/vX554M+
YyZyTMaSlg7ljjebrsAN1YkL9SUuBl9BW/UwmNh5MHmHlq5iYWZnUFx9mQ94nSUdQbxrl3gc9V8y
djrVNkE/PqOLlAXopZWlH3rNx/Zpt8k8y4DWtJ8zcXR5nrdqGjwC5B+V565YZ7uaPEsA04Qb2L4u
S5diRap4H+XccAnWwJ5Tn55RjHHPICfzJjgamjQ3cO2VRrMno5+Mdyj3F0D982CBJsIpZVuqmlN3
S9W5PDAgXcN+QZY9HeHgddoFH56vBfn0THnNHrbVDhCLfWDESxaRMONeR1rindIQRVG3Al+iQ0bU
TX7sPSDjmW7zq7/Xb54m+D5rV2b6IiiWmG7SzBQhuiPVmo7pcuM8FUxukdMaByCWSHj4dhip/Jt6
QJKek7ND9BwHcuS1la8KEgvyHlaCvYatG97U98vpIasbaDRbhfVu/BS+YValjhn4wqe/QsiWL7S0
Hmy8XQEs28hzbI59PkSbqJE2+VeLGtid9XLKTY/beaAIT6BvMKccDtrdGACOhpDGGkNVhrvXGLRW
DrT9x3wor09XDKv4wnxUYbfWWIxpvfVxoUvhUFphvMr5VHcOsLvSyw88x2DNyDzSojjpkLBi4lsx
jWialZn0w7uWd5NxbAwiQoxmmZGaUc7dt3kJaxLwlT4FVn7ZneXEBeYJmLejFgf33h2iV7t/0XCx
0lBBUgyXaXymWHC3MmYYB/FkXwUGEseZiDJvG2xU83CR3GD3630+L6FlBjf21tnDNzF19P4qNdio
72Ozt54SGopMZ8cAFPemk/c4j+/hJsB0sOfYtwsMmHlBa/HaTyfif1j1srC5pmsCE+7VccXq7D1k
Vh0rZJiJq0FkzZ5QlnU+vDUnPErOJlWXEYAZjtDLZKS5/iTg/ZKNjRFyZykQ7PjHiSB5JNM1so5a
Xdw9YKt0dIk7J4n7+um13+18h95HPVv+W3JYw4e4rv465kZU+grVmvPti/vdk2VfCBPEaA2OR1Fp
sIHqTBqebQzfuaytAoQkVWWp9Ze+SVJKGzp2dtUhaVzMFiRQLB/N4YZwUvq+1eUDkXag4Olztz2p
S47SmX+lNZI/Z4aetZtuYhyinJZJNDWmvqPTN32GfoQuGxkzPrZg0rh9sf3bbtL1oyV1134hL+Fw
+577HDkdZz58RZOqcv23ax/e5UzPgS2bRgMaIQSWZsaMM0iDdOrAcBDhyaCNUHxV8LsnmK1LWLfZ
c3uOvlCDuFsQyAUawoxKJlAmZQPpcsqKr0QghD1OhUAV43qExRwwlwQopzPkoR3aPpAgmwdDomXI
YTfQ11mFz2xYVxT1qRFXT0Q/YPXlL+7F4R+PFNOALW1AyXxoDi098rk70/RcAIJ8zsr1z6VYt1uP
++V6Hz2+/Nehun8+DAmb5PIDHEdewptJfs13xXbZwYvIzuScUIxPGD5nGIcejkgo58bUrNKfaPnx
T0NYKN7RJcKAmTGVp2oE8x2VTk0/7m+zMAmhabELmTZhlNPEMhlOVOABWQ8RW7yyZwhzpS8xqLPu
KuJRJfPMNr6UicdLDYpt+daSct/4VRVYmNlhYE9XKsM1jeQlrnpR6MXPJH2lshWbQO0+FI0MZtUn
dXmsl4tIG5gU2SAqWD3QEEqAV0PI+Ba46QMQwvc1cpZLd8TZZtjIFdQfd7rZUOlQerE1H4ejjOih
L9hvv/aLk458VSORY+EqNTjkkXVH3kLBD1UMDLlBlJyzU+onCaPJ3+4Y2TEoUOdJ7JT2o0nUgbCX
6dp/24zO0M+xVpYcH05btvHMBHwvBpwlHVn4jRFfLI9bHwLWqJaP0KkTtoIHCFFs/8EFyoVHYdaA
ALpukhefoiM/KjjdySPDTNJOAV1akyBW88PzjfCj4g9qrgeL8jpTXN/xDHmiNhlaAG5oVYEDHDz1
aFmc0mQOpm7MGHzLt6e1XJIIQz+6KNjnzQYmmkIvj0xueSEHji/3vgylt3HRgOAtlKHpdgYMrYpk
FcLD+D4o9QlxQBg0/PMiqMjM44pJgWxRxwu+CrMbinpr0e8SmVnVCvptaeliowMbEmuPfZ+tXQ4I
cl4cvWlAhGhUMQdJA6bQUBvyNfPl1NeV2U7KUvq54u9uIA2s7gjKsj/j55AcpUn/qzBujV1yQcqB
BHdQsbUsSLLeOdhmiJ19sFC39r7u8sheHTlHAoTr7QMSH4r7GxKIsoNJhjxx56QJ+wQdAzH2N9Bx
F7m15OpnBoGN3TUpzwWmy77v1HgZaw9Uw05Xd+pmWW97uekodMjrdLDOHOx8h5w/2qENNMf3KtEE
nyIHji4R5jM9soV2x9ihG4Y/V+4z9fdQ9tnHsEtuxCL+hAP6dIi16j9EwRci77AmeoEhAhW9vswu
KvOw6S6XaAo2KOWCrcYq0wN/8YxBJrXs03ZvZN9eEFsgT+GKvXHX4KbssnJeZReJPAZTJB5IMhbU
8Tnx4kaeBtRHK++P40xNbIqtLxIoYTRcbCGjvJjo4rNNYuYogkXRBbk2xxHT9iNOijKZ40ruvoDb
qpovjags8recj068aiw0FIICR1hLAoOopDwUQwBePk4JtYT7L8U8PQswd8ok7suHqr27vml0Yn5C
k2vIFKkL/Cjwx2GAjTUpf6PHcS2VYKBe7kQzm5wdRreOAstzv/+dieatHRrosM7NOlvoio1/YiyX
QtL6UK5rKF76hFmMCQGkH2LYHe9VHPrcWYC9csU/dbpkGtDLoG+0QSW1TGqubxAFgBPtOYJ5evkn
48fAKWQ4Kr9aK5tlTlYulNtNqlfFTr9cNXhMupPMPz8SYtIO+zBEy/TEbfR2QVyBlHzQLTeUls8F
taFwHFJi7NTPlB3YVUh4UY5XnzSQPyA1gQlHexQlKURaDi14GE3R7OOzjZSA8CzQV+zquxShkMz7
bqMKFotU/E/2uy4esgUrTdFEXH3TUceAn/lZp61eL4bB1sTRj3NPYzuJSwyeA1ANkWW5KaDqLITl
lnAe0kAqat/fyMdjthz20DSmVkDntSqLFGB3qaqKaO9Tolw2LNnfOgWJ74KgLual89Z65UvV1+AB
tNzFU4raWmpV21W/LBAGpwq1GBQJ8KHQ1zqghVbtNMCntvmZOjbmdjl7PHAFhfxtbdxNEW6OI39W
5oQcgIAqYuxicB4NfeB4vfjGKvNHwUNQMAHGjHJUNYTEyxqV/9IwhXJ+M7C/ptcRPN3oB4E980Za
Cje91C47fDZ/mpuN0PNwQ0m5co3xZwYyf1a7Wibb0Wx+XBj+UWfXwIeTDOq42//nNj6ruYhGQI2F
bpVSmCI9MytS8G0u8D4iH0dHLvYmCmbmZhNRBolOpUFtY596HxpKXrL5B+7kBpqKJz9Fb/38T/i2
W6FnF6XW7HuDcg6KEGa01QhFhTfl+s5vVhbsXLggPWpq32wKUFZdK1Zbw3n7HLYON6JTdo1Eo6xT
PfTlA+LqlXlYinNcYACMo2vcCAuazWMz5kXKz4OAJioPa2a0duTJIX3z8PNQFBT68qseQfqwoPyJ
F3LFt1hd8BJPsNEsJoxwDfsQwl+2jTcFWakwwhzZCp3rIZw/Didvvj4dbosq0GF+JXvRKDh+53jg
JEX0oB3vpt69SWd2sqbzCaHFJ0ksYyGhzdx5beaOTpLY6EHJr7SHq+L+x/uU5cibXGwv+Rg0Tllj
HI5+0NHfXFnYLRday7QEHrSm+YbcxEFaHoIFqt6S9y8dkycPYba/aAIRbIF3GsJp3R6PhuLlzhJR
cud4tjxADfmpLTRZtUqrpPfrm33IteexrXk70Purt1FqkgvNNZQcSj9hw2FmdTf62iHexe2XjLbF
IbFg/atZ3NazY5kVykykyX+huBojxtGgq3vxYepMLsCOTfPofIK2E0yn505FUaba9QphY33vFUjW
WPKl6THkyuHIRBHD0QKvkiG+r54l4dP0FVjkLRhwaxEx9vVmc+gx3GxuP3zSAcjnsFmk9pSTY+aj
qxpF7goMzVe/RNU0Jlw1cqcXZM8BF0vwg5G2h4arCQxj80+CgTk8yY0pvuXdodSTPp5DW1pAUaae
8vDRJpQ4RLtMk6twdPyeDwZziCjbLUT96wu8IzmDOHuei1LFmLRecN1dW5HJ2cg6TasBfgJkXuYG
uwBnsqruPp9gl3UMoi4lgoOkoBJ51w6spKNWq2OEES7Elpb/ZERGNRKPRWz4iW/by3jqL0a5NXd6
vjH46Sddy0q98q6ec/1m1tTJSUahCaCS1uMTRlX9dshkJw/7jblYAQFOqyr6Vva41XNxWSTf/msP
AKW/7q7xM7QHgpIwEfAjuJmwrg4s4GqhUlaD7Fw+TCMjTIu2rRqJfVTQPh6NERnQ0D+2sNkCeVr+
y0oirVn3SsMB8hnr0f0uzT18qg8LI4EpYsrrLbH1vwh4Mvfx5pgULszkKvZl1488oOPfqiq0v6dL
r9bd1ixyYD2WElFZWAqGC5zLVhB4vdiHzLgRf4Vu6QO53rh8WaRdxHuUMI0CVlED8kzHtaailSbl
E6plUvRInuCf6/MCUd7UWUHHhKCTbGmBJUtrifbmSYkeflQAZtudXCCm6mWLsr5LoK3rnIeUKbzM
oFaOxAUKQhg2v1snNpG4AavOWaCj31rlcL1hkp84YFMqqSXfBHk8/3lXfAovKUAOQdAEt+pXSFvH
VIEarQc18Ein60p5kSLhnglVh/LunTIB6JTcMj/Y8tOZU7eIaZOPM194rVt1iyYm5/E5aLM41CDO
MP+ZKL/Z6URFRe/cVN7R3MlQL7VWo6LUwPKzWRooo4EISPCLN6OCx1aN7fCcxX9v6edNBOBPWvqx
So+PzQjM7Erfr7GBbMhXi3GJ6+i9ldwVTqgRgTBO8XzrJiaGS6Kio4lS/I4ytCkJ4aQjWPkNfeX1
OFDnvHrx3SmDFmCpwamWrlME/FSERGMKZuCn5tYE6wGiM05crcHJWVglN/rcqqi7p5Ablat3jTg+
rvXi/77E9cYrEJIoH+ZPh4hBAsyFq5rH6W1AYxkvsaFVARQAL8PbeJxb0YopaPBQtp3Yb4CpPA4f
bWIVs7tsf1WcXryyuvayWP8WX0T89wOyfhKIZjJL6XCqTGluBq/74M/z+bRYzjhQljSv8qMEN+N+
A6hciYMCFprYeISH62ycePHmn1aTQzBcFpORtt4sRW//iKmG7UvdLZ62DoDOaCxs3R0snoXtO9vc
XQ4LndDYnU6X5rEW311jFsep5WcCJgtih4fR5/dONW9kML/1LM2n+VWvjQgdAv+xtQ5cMFEYPaTH
8uT/3TFwRGFCpgChMCzuvMu2n1WCdEkhE+epCOxaARqBXdIvEbUky+WNVJzxVoMLe3v9gLiZHmIG
WlHraKHZrxcBlKKrhpI34wAEz9iqM3n5feg9kzK7Zufpl7+HjfsV5rvNerp7A38bBPJRmZnkmtSh
poCAfKi6Tze6kMbnV5+nucD2NNQa3i7Mn90jR2esmcolV3SSw+NnsOg5cNHqHbG3ZhGcGRXxXDa4
oAqlxbnDFh64NTaItsj9HzIJG96j45yzT90G8K6cReBKMzRWx9Tn0J8YbU9qxAKuC+3TBFthKKMp
o0oy26VAN9onuwOrLl99VMDEfPYUkCyNznGMXvJ0WqwsP/cqzfO197Pbhw2+wiXajHC7ertoEPFq
dslc1Wlkx4B+I5oerg28C7yFzvdGeKengCljjhLo5b6S0vxpbGRKXgTZykU2UlY2+P/hk9smH2yX
GlSWhV64nollAoEkXXyMOnkC2nzA3iiPcxkyifiXPO6e47PQJYA7oNOs7uhWnEourrnpSLHgj5kt
Sggcz4FRivjtqo/uCY/wAtAnXdAFvaRB2tyhOYXGTPPg+BV2QkHyFvL3tphLmQsSZyKwKOmWwYQI
NtflSHZWqogTcOWLl09Q2IhRBKT1mQxTqNBFdNRe30hQIB3bezq437BNbcspAnkKn+977SxwZdzh
tBqWkUbLLY0p/Rb9TngRWWH3mYXJrJsI06aXi2ytQF+oTMUBynv4suJ6AdhWUSEC0K5U3Me/leXe
Up9O8aMzFPOf6ocsj1eCOASk/YZ6nGrdf5UPQMYXsDVmjpKDSF9XYjfKdNn+Y3C/K1DnqgLNTVcG
j3Ph+cRmxbcftIiGcFo4zUjwzNfAqOtjkZlSkqxWLSMMV6aTZk2CUJ04zqitDeNssaiB6V96Zajo
FXpItFqNE77z/m8u24Tck4OKxr8Z+3vtTOk2caw1f5iTsnaS0QxN1c/9UcYOpmbTmWJx4arcd6bS
ozc5Uo8pIP8VKqnwVbaA/uakS/pSkLI4aKIwf/YHhr0Kx7cPax4X6+LYESGMjhN/pkbqmOECosQX
HDqtN7nQYS9axaKadeZBzgOc/N+Du7ZAoz+wTpTGRL7MvWKYJh136fECQrxyK9801ukAY+OPpCqe
XrL+iMzMaC6ByJQkAVmqKYd1zUC0ZF+7PNBhLGT2fzqyDy4LGLJpFgHOwCjmVvY9m+OKizivMMxW
AOxd1USI8Dc/MwQklO7/4GyqC3JWfmfRxkiUWtW679I+9BM9OM+H0eZTrqCan4NFa14hAHCQsYFo
4WMLCkX3mXkmbvS3bXi3NcK0ejn2w5goU5ODPPSAQNVV2mKceb2ziL7CkuSjB0Ekbf1JJtwjTYoK
WE3WurmOVcmGH17oK6HwXSlRCFShZWQ1jhPryH6K9ZkG3rirBKfj8uskluGE2UvSC5uEwh4PQLvW
rJa1JrrnvKAM46OpYrwXY3qAh9xAH/OHdF9K/c2oP5ddXSbi5iB0X7SGMjOzMwWwWqnYu1E8XFYQ
PDJREZhS34tlW9KIG2zT/p80aMdlBbF4JvVwEER67Ui+LwbN50euuzM60NIOq+iL1DlZ1YVHEpeG
6RPvBjnO4Cvo4Ys8fVnyVN+xSLW7C0wEFSE+ynjreSfEgUdw4Vm/RMKg0Jjtm9krQ6jdIHbBLXq7
/59FcHKiYKuZikSL5xEXgEi5srqUIez0r57zMN7GLscbiB7gGA2VV28Jj6vYoMW6jbwQYemJMwo5
eZBAZ+wNfbWBA2vpS7vE0W5Hypj3XfqQsnq+Mw1Fa7l2s4ZeogNAfUOaB471tMBUClF6lTmzbrlL
LYyI7YpAXKsObvtazTYbPHqxWla+L2VDuHECcF/QgFrX0GYPNtt0cW+awinBtOZ6FYceQdKFpSGz
fjzekzmhrMUkIoZ2dc3hWBJaiCejPjDzJVaxXNiToh3EbMUKBc4vlzCMIhodVZ3n2dSnKbKj2inK
NG2AZ7KYqMBijmW5f/CPACUN5ge7QRMgHHu/4gnty6trY9ZMvhU4nYURrHHF2ZxNQYToCaCrNFuv
+TGAyhF4A/nSvlcxzRtms43/mxfQ51TEDmDivKTnis6vytWrmyNK/OfJGbabUcM8eeUyaF81RnKS
mbPPpU590a95EV/2woAASmngZJf9biWaHCSXjRrKlY93EM1hHn+yZb947FedrcaYzBGz5E09XG3U
NDvv8AD74hEOSmXoSlgGwXZj8Jcw8eoK0jiktEqrGUQxCVHqC02F6y9nE1f2plXaIbMbEl7dh4aL
MH7R7Hzopd5RR6Ia/50PaQ4jJld3ElN6bXG7ZtYEkQmRkKcnDAludXyTLxt27xl7WAehvr6yq/Go
t2OP0ZGCV3zgZ+wilrBQBjrqODlRAbpRuZ2iQtAh+B95JZvQC+vGmnk37fQw5OWjfTcjUKapPVCs
8cyv5fwN4mliPTW09eAEyj5UEQz5YH+cBWNsYSMpILYyv4lfvL1/NIV1AweL/HLoszfBT5HOBX1v
Id4jXdF1Ki+saKB8krd8sbKEGpO5iB6nK8MvkFLhXPanMmkPgi1T1GrpCQnBsTh2H2Ur76CBRRFK
tX3qEF0jo96OKyujZxTQ+o2+YDe2s7gJrTCk3oL2mHIzs3OOKhdz4F/5HyjPii8448BDpoNF8fox
CjiAD4RLQfRDXiAM/Rq8PIc5f07eNbmoWvLpErHWXBvrkPGPy6yvNeO04xFvSbyxMfhaEZ4mpS8c
nnu77/Ph5/fun/XufHC7P22Zo/tlkkVTuonI+axeHwVj53CxGGCwwsY8Eq4mDT3OZBXraK+4/dyw
U4CSKbY6CYMSMkmW3og0mHYGKyLtXhKr+lk7qzvF5Ff8zulKRPfJfatVS3n0orSFXuy6p2bsu/9Q
ETG14uYuUBOu2pfD5df7+Wui1T6lj25sRs15aYE7AWs06pYrOX+WIeWEqy6kY9WHZS97+YCdOU6R
1z37x48FyFOtpQJPQcFoAyjc90xs1nj9I44GcZd7xIMdz5nPszWLgeCKAZozLoFT26toHaEFoRyJ
Ihqb6AxAf/8qTEQNIgd/k7W5uwiDPDM87eBmVZZCSZgWTJZa70GJNFItoz48PLdzSxuo+0o51wJV
v/LQdoxeoE/QniVc80A6+ybE5/UOPG1hj2eWSQ00e9fl+ex/5mdoynTjnKaqUtVff8AU3o4hMzeZ
lbmUN5ZzNgKl35ptlfXUvUfMH4/b+cDS+3SGfdt7qScLhNFc0/bZOEE6LTBvqNtObvJfBrJVI0RC
dutGJIY1ce8RPVu5h4DlgCfhi+vU856ERKa2t7dIm3eUW3GJUvOE8VVHxZUPbbvJMz+jLx8AuBJu
cs2IzXq2H8KEtDb69XVkpFJ6GBcv8wYdBZjLY6R4YuF+K8C1Aa4uwzyn97Qi+pHDzoc8oZbBu6pI
zNZWoUpXrPRPGO6eblIf7x4fQU/kD3nezETHSgRXsdJRG/ManHgTUkssWxOKyTC9nnRPQcTUyGQN
kG4oBehw6RqVTSzJUl/VioRYHMGR/FkbwgrJbE1sr8bNzrtcVSV8pG12MBDGh+q6j0qKSWZY3s+t
lju+RYGy65KvYV8c201ce8DpCkhy9MRQ4L07/vOZn0PUDiO3xLCWMWyJ0gEKIA8Ea5DjIKIqXVEc
63Iev0xVSlIiibwz0892Qm+5r9FnvUzxuhWi+3laUCLIQkgkMJ0RtVzDdny0T2FjmptZ+olH6xdv
bPSb9Td6YdyQ7jH7xqM6msfGeOAWA1MZ63WBZ9mr83zN5fwqHAsHStb+QhP1tVrxx/OY8KxDtmsP
BajVtKQ3/pCO/1VvI/alZx7B1qlQ9+yWAmpi1tK+rs+5Clf+OfS8XUPb2S1AzbJfgAlHTZimXNzh
+FeWaSQ9caCZtcvw3byWjV+mXaPHBe2ypFhwKxXNh7HXq3iS7G0PsQoiunXoz9/wAOGNKz3j6Q45
u0A+RModZlLuLgLEcAx7i2QGswG/yYeOxDaWa3E3Netjw+lk/VsGdxeGOOwTCe6/BZUQ8eoKQ/Mt
EfFTjjpOwYSjDt8uqAdkhFllk+l0mLAxa2fVJKrbkTXZ/zDkjw9QPGV0wtINqhmQZauMd6r8Aa4T
UPYg303pWxS4d9aC2qhiv4FR8xbEcjKhZTOOffrnuK3P+yAkuALcPOFvfeE2LDs0tBfS+5KCNiPq
jmrueH6UtyVFfv9Pu9lSEcBKrXKtjwaNYxtHdUItAB1IO8En1iIMPBuC7090IlAho8edLofK4zEg
w0M1p/TOPo4LS87gQvJEvF7RdFdH7MTaR+6mDwizQ46Sh30XBN76Wgo+Jr7iv02oGlP/U1qMdadu
nBUgsNO1Wm1Js1dV/j2YcAuh6k0JP0NWpHgr70VjVh1R5te2kB6ZX+dri0BIlJEeCS79IvaRH95g
uZLkLneHZXxQc5MxziyS7s0kD6uZwKgC66U2lnr0luVvQVsa9mJD4EVBDhkqAxKosXvvGDHDzVti
S+AwV+zJmax4dtrFEQ2o2CO6UOIvOCwz9jbtglVGAxWAejrKLD+K60ht+qnODjGe052+/0UV71QE
qW2DOdMA2kMO+pahWAyowKMezPLyoXdeyTagXQBF1fIkct6KPxuwoPMb1FyxZAm56qcvxNnT3oY2
nqwQ45Fvn+V3I1K2WuD1rbsYUcCLEOZVOU5zdD093quqm9Yb6ZCTLVsBkTrVrWHOuXgUsiClV0RX
K+YN9un34o1uZ05QIT9msjZFTodgZ57FjRe+DAq2E/PHw8hDALs/W3nyAHRFQtWExvnIhwMEJ/J8
QYKa8UqZrvcyPHpZ0oNZIiJhorA3A9qF6kl8NnoFYajXsA8x6jUWiUb1TCj8tgzS8hOyRaMay25c
ASiT+TVFns49ccLFhCpU0QLju2csG7wX25AFKR7+Aypih0/wIbZMYSo5WnvckklBml/Eqx1BXK2u
5JaICGtPHc0XfXa8dmlQXXlynMVIyLI/WjWnd7jbQzXIKug7tNSGUP2RbTqPf5pyXp4em9MkMyvG
qiaJ7ylFmTsWxSWqw6K1OTeTQtYOPBxwsSlKb6NpTFVUvdUDaMadlvSY2zzplY7LFKMtWtkgoqUm
40lJLoMcC7gXYYWiSYKw7RDr8yuMx6sFILOWGv52Ftgg0VGrsnPqf6qLYG+2jIFbaNzVEC9LjEiT
FPFwJz3o8tEaZ3KJB6k5TGfPMkh7aJQBGq52nfy03YnVF8Y0gFTAF2WfJyz4T09T2IfJlCb2ew8B
qgNJMBbKqHIGDrblBoU0Lq4NGEokY2Zcveqo1mt5+9oCXHn7F2eQirQ9Drdn4trJvNwHoDR67ROV
zK3m351Ncz++7cd8i7Vg2hcpF+hGvZFNpDvzuhjacoASrrFh2I0E6KEfOLNp2rnKahFc8zyjsjz3
LgYWAOE1/kJUKMMONF29qHMxSrValauR5EHbX5dFUA6aAm/k1b207Ik1jos6dl1G/Hs219AlhIoO
w5h607qt6WVRkO5jC8eCEENRPneCwZX9pZxifGspQGBZ+ZVoVBNGlqHiZvdDG3L/eVr90DnyFC7t
FczlBYaVy477+8LWni5e3uq4xMBeaXWaEve4cPgRql4e9sAJZKBfbgC4swi2Jf4afiNat5K0QsjV
VRXRwdzRtjUhRn2+ZpGDm5BIhKX5PaEgvGq8PW3hiCkWkb1iewVWn9ztN46KuCIlctclinAJafyn
dxzX3FwiYnGNi81Q68Bo14szuEkTZyh31FpPOzBiQsl9JChtJuwgog8N0+aSRlC6TjKCRJFPuhGV
HAJuj/jkuxQTAMr3KnX2BcJ3YhjE5ucU/rFCn5dN90E+Jrk7CFp1IXGCPd2dgKbOMW1E0JJUSEOS
SRnWj+d6Z3gCNItpLH4Bk6Jp/xzky39C++Bbsp934PToMt/CdyWkgia4zc7O92ESrwoB6quYKlyE
PueppHSttRMgKDbqDc1bnIgKx23Scb9fxCIH6I3ZyhMsXBxg/LJvRQffeHT6nGsVlMckOSgSyWJa
nWOz5jvmS0V50AQuW0dAAwwHPqqkIrj/Vcqh07/rK5Sg2P4LRnWFf9icV7WOhr7uJIAslsNoT441
PUZ8XVXWjdEjsn+L2/M/iq9KM9TMyMl1hb901OWFIAHil2awlIkGB3tC3Yt68GNaPOe/W0leOCwz
YCwH+uM9IQ01JqeGOwUjf+xW9NlyE1yF6Viyj7Mhunj3EHi7QHROhqoNoG87B7B3AN3Dbo454L8C
gPeMvsj3Pz9V9qodr6Ry5MJizTLyKyqXPZmAOdkca3QQ8HVvU4AaIEK51RLc/nyBwxlIL/suyD1N
t1fBL82kYDpK/LcbOel2BmMIaNFyKe5MA7f0gD5W7qYjVsIGGS1vx7gzMwDG2r1h5e/EKR51ouEi
XRYQON393ZmS33UrBEqyq2z5E+rwm2taEtdCKZ30rT6v5iQiVrTPeRvINtYBlw5EiMtrHxzb1Otp
2f+YqBZI+ASBvXlTJRBEygAJh4/ZYXNVSS60ae1rfr7yVYYKakao/LusARRDD2yLikGH3dY6+EqB
ip6qa6PglZyHywnKbPiDxPTsRGIHnM67t1wQSVmgqKgnb8kGBilUqlXvUfO3dSTNyO+yyPIkg72M
EYX+kHd5a7Id/BiIoYEbMpU41GwaiCcDbmDGDmj3awziqRS1TBqbA+Dz5lNrmJJpMLpRoMqoWqGD
ve2EF2vpJWe3LAtvQ/Hbz8JBFte5aP/whrpKjTfRtGTYy703WuozMQSTeuX40km4AcPjYaCL4tEI
TAd2IBgQ0Oyix0ZROPHpzR9IRgU00CEswNp7gqWKLVkrDFJZ2JQYACTyeYOQbkpr5mzdMWSexn2t
DZn5XlCZDb+CTMKgpqImr4EHD3NFsmseAfmSKxkLNnfEh3QllpF7NPKkKDzNxPTuGjlpnx+hElrC
CG/5JAFFkuBQvPqQjpI1kCk/poJ6q950/sbQPU7iTMaQDRGMA5+1LKyfuhhaP74x0VAMRwTA1+Io
l4FwNlkYr7yEsAcdfqmEbWAIn/jktLZXcNMaDUOZ9oGYORFtTi02+Wdl/ccYthCf/kfrIUTdOFZJ
moypVR3YTsWtxnRTiJ/pp28vkBLpBLUCTHynrnVtPkuN6TWWRsHVgbRO6u6RAI19WDBeOO6ugzeF
0nozAlgE0QVJTd0bNXhY/sqCE5qGy/yQC/rk9c9uGFgxK9nbOWjaBoitZW9C3mJTEKjo/pj9LFwc
CNtEYW1r2Es0wP1aCDux+fDK9ZCe/LxcFrqjMYEUWj+5E9kiXuKGq1Co3qKX+u/MDdI8GBoEJDdp
5mN+vd1GX9YnDcgKGbWDNqECX8dwlXD2XliOP+bwfrHJ1GaCEi0+q3zEseUCkWFn/LRUlY6GilNk
Mrv9nE4tPzoMhZlmzo0cv7OJlM/KqwmrYHHyXrvVbd2lbWLhvQisHN74kn43Jj4FPPHyX/izdGq+
AUd4+aktszqZrI8DWcl/2rkZnmQHjKcK5JPLYY01N2Xe5lVUwq135b+/YrpCfOW2qNsV2Iwy48Ou
V8BGRlRD+xwsLlIJKp2mTCuSWULWbJR+CgsAtj4x68R96ve4Zc+yRlI+QwLdc+F5pNnQ5177Rmdy
AyRdgzxCraUVRN0W7MO5HlTmUm5ff/LZoOn3ogfqbmXH/BUxvN6+nkYYzhoarJ4aMji/KMZwt9tp
DzUAVg0CdvLFgacY46LUY8bda5OR4ftR7YtCXZep6NV2uPRcfXQgcQ9ongl+HTgLD0OpcRy4mioJ
2xvx9jKlu86mntGOYvEPIce1XplE0QBlazzIpsBpfttgSyv1NH3jI98rC9QUjqdh55jj1XYxxLTq
/xwZTbl2f+ZUshN+xTIdHXuahniizIkA+/tzY4Q3zAuIhATC+6DqJQ6fJLohRbeMuEp5cJkXSkbs
VSaL15YQVZishbZQrt6GNwSReRJi1AFDXZYBxc9n0yQS2qqIuiiHCyYWuqSRFbAbhLewZaSZT+D0
sgQlQHQAEC9sg/5btEa2Eg6j0M/LKiakj3FseiGwR++dP3osnIvMmt1WiXUI2o9nSBzjIqmfI67j
ojN0XrEonIrZ9YZdfERQaiAKFoLWUwQEVIIzJmGT7+R2Vv2JoKD4gbqvvHJDohc+SH4zCVD0wXG/
ecel9AlICNzQpH8iQ3bodN+fchj2izMBiweSHS0Z4A8ODaT27ql16Lzues1ljAalJTb20lkXFVCp
lXxkbMIFt970p6U6V6n2MWAocFZJW0JUzurMlP+f5Vm6tMnCbPkCjlluB77UJ76bctQVwXw8jope
tms8ZPcz6N4CAde42bGqqA3w/FAk/ygoLp1HjBSkDUraFkhHNPzGFPdxqoqIwXUovVBmCkBrdZog
o/GZdHbQsSqG0yYvEdEIO7arZG1FZz01lDqmvKsWxbb5m6uUap8fWO2uwa5P2qNssZi+KLFQfXI0
Bn+c8nuMpvneHM4kBNKc4TfyDnttNtGTS+uerVAIP6IpfyL7am+7mU6tBTl/0jJpg1aV1jzpuN8M
gydbP0RR5VZyCUm8CY+Y4f16drRtji5OM9HCfEo+UnuvVFh8H0QzanassRxITQxm2rENTr7jUw6L
kD3BIF7GWK5D7Y/RTNAuN5XFkkVjJ0U16H5YwSv+9dEuVuaXV5AQiK0llzf+w/O2KBGHtaN5iax5
fIY27dJlfEKIYPJ/n9YeQMfgMqW/6hcal1ZQOa70gHYQmQTxcVl9qJi5HhyvZuUbedKGEAVKPSfI
gGt8ZoA+oI/bx0ss8Zwuj6NWs7K8dmCR3WnsewUXlT38Swjzb2TtZs89alSel5PRpMafEUk08oJH
ekgJPndXNjMY17Gz9yvSaJcjCZS4OzaxTGZElSrKpM9xDytio2rHtFou1pHuYSxCIgXKIUj6EHsu
U9YuOkcVsOkYucNgyL0OJuPV2my2x3l44PgxJSRndjaWFy1d6YLLSB6TIUZOkntRfzkHwGprMtu7
fUDgoME4m7Bsp3iCqvCOtjFs5aHsaeAFBcfGxAC6Ou2RzY0bdYgB6GPijtEsm6rWj6zjBm3nb7bo
avjSIGmjASbJA/dO3LyqQIzsNEe/ZawTJZpK+yU8Sg8n3coDVekhJHdcBmBA22rF0Fq8txXZk5ul
BPpgZmrkB2eG9po47dSKMdZKH3SEuRzvY5vRVDrkxOd3vZRMUAmwLMoFfSkVquFLnmKB1pYgN+T3
glm9om6OW6FQJhOeVEZE54w2a4CdA2IGyLdsbaI7/u5xvXIG2rGY4w7yzRvV/9PVoPx3SUYaGbbj
NMTmjvnQzjay7XPpFbHZ/zhsXweaC6AHaIPob0I1dmVn/RHfTjke4LnA878dpQikHvfld85ZbB2n
/PQWZrgrZVdXHxK4lf3TPeuuExhmTbi53v+nmkBqxuNQu6mmx9T2bzrPIBjDySQDXqe13GEWogPM
PR2lBk3bwxEVlO6MNPxclBmtN/I2NhgRl6GLe9jNVWiTSoKdDSlRgybwwQ7MpJyXkoUP6SWJaaAW
d/Rt7YiuFX4aCu9FhSGnHqHJ80xtiy/MQcLD24WOg0qx4SBayklASGHgo+YFyosCik3ExaW6ocsX
fQk6n3OQ0v/FKbKNgE13RY7xp1PWiqkaYRBVboU/mcEIK857uRc929PKdJsBzWWMgGbn0RqAgCh6
mCSNODxmDb/Ly+1K6Uk2wmKyv+X0+l9tf+j3WeDLg69OOYOY1UQGYlk2yKmWEqeg7pnFrBWmjrUy
kE+GhmQUd6rbkuGh1y3yCBhZr97Pxy3S8QTfBbpo89cuK5W42maHHqjFyivkTkBS+LnsIKUQIFw3
j0elTD7xO0moHN3KWUeUDiie5DLakraEn/+69juU18FvM+fp3HP1MZzhjq9R9fXuoBJn0ltflLQX
OGXdq+Pv4Rom36s4nq9BKHolo25lztKHCZAuhmmVcuW3GIDll6jsizW5xQoDY6xptzur3pXko6dO
owgOHG8jUoQqAsS2xlSe/6EtPztNVYRKV2JbXVIzLYr0SM3M6PMH0NTtUzTel4PmHJOdriCv+20y
GrP5/5rhUPguNdoiHcBy99OW9yrAywU+dzt9U0VDg5z2SiyamAqZ86dQ92dLpmVlZsAxDODWN/Ip
sJ3Oc7wd3S0mkm9kxgIOY9ZG5D1Zd8hAOEPlnhiHHECbphfyG4nxgdg1ML5uVr4UTPrXTC9E6pbc
qZvipA9aXK/doEwqEpfKvQeVEIPZIV5gIZc1Lgxho3j9xycVaD/Z5VlPyILGAaQjpSTOAeCmyTPH
JwTPulf0YK6yt65bnjj2qX5JjXJZk1rwwfbWu69Od06SPAqrQQZX3FLdMXXYRgw1ShJhu8RLyQwR
BZFsZXofPqgz15B3QxbY2OSTZvcdGWQ+v/jdymhBiRg+c/zjlS+osweh77cm8SyI55u9BjHQnbnh
N2pXEnORzxtsRi05sjf2rnvbPxO+jbhWFwnlKHwtqBcj0MLI66f0bzGi/1I9hujB7WZjcOkiJFIP
QXWdD6c3QSej2wyIfjoKto9Oc5PEWYW2PdbP+1E0KePIDIMytZ/QFzTdtW3fCJuLdDmD7I5m7h9x
ltaDXv9P5W3EA6VTOiFrgfI8fNPbOLFqV2uf7E7C/jT39nYWQ4r/xdGbHcdXVoBRrGvk1uQ0o2St
melG/Mf4wh1rfqN5vxIkOWjQdmCNzpGWOlD1SdUH33Ula1fCORRrscdgy3UA8BACE/FPhhp04aQa
zJOC1RbhaqPRDRGeG5uOd/TGMXv38QW+PC2jncIeHKvUS4hjfuGPtTWD+0qLAUBA4vSIqRUtYO/K
aJ5wt2ZtiHqzS7ylDqODklPjKF/ABq7jP9cM0lR2purYLlmvDxPh/YF4Vltbcf89O70FywjH3jKg
Z3gqGXwfghSoaSaSlTQk5J56gjyGPR0pV2CzcMEHdT7YgpRSnCNHaXZ7PSgtoPgVdB5Tub/3Ulih
RpneNGZZJ7TUmlhrrp+jSgNU2KtizJwckgiGual3OS58/5DLeIucWJVSMeE9aP4tiyeh5LbXaADf
hMfya9idLsuQkKiirpQp3iWbsxuDWO3RpD7PFLp3BlhFHxO/YsII5lV63rfJk94Q9FDXwtburB6k
mxXMIpYA1Jhni98F+Byyzq8Xd5ZIAyJgXxYpXAN5uXKPNfjWqgy7+PFRRoivUPKqPYrRF6W02NgM
9NwmbYqVrP3tsWU1nL7YjPY5iyJmm5NTu9P44MBcsu//zBj7Gk9LgW66Lv12hlimLVNLT/JCpS51
ltwMLIZSIOQY/XEFwDdmVo3FOos3fcXkUYs/8n+sfX3HZW3pozpODfDKXCc+XW1DA3IM3+ubpd2L
/F2eFD9FyHlBschJGYP0czd0eH9xd302iijGm1AgX1dfeehceEiNOFVX30HSzy37ta+g8IlB5i1H
pmO64+QUu1N9Jz1jYUjRNvop3tuEo/mXstbGh1x55/Esfkuwkcq1r9rtFipUsQU3fMGHtd6H4zfh
kZxx2ktA7iVq6vSAul2njgLpztGYcfEKUxSBlIxQoE0PrMVya0lA8/kVCWGK5uK1q731HexulxUM
0aJp6n4Mb6r1rYEke5Pul6Z10FGrU/h79yvTP212QjAE+AuDgIzHoSP667msDD62yZtYHOj8WTPR
sZsDdcRsfA5tjjUxXUjIvyihfX9VcAPqBUaK6wg4oskWArJmCh1EIaxpLTMl9CnZ9n6qk4AEZOBg
Bk1N+NYvarrqfeGNByKP07DmyeaNuMXQb5BhOa6IsmemcUHoFdI55ybYsy74EcWzPCsa+YfAtqpU
m+xgJVT6hTmCFEvA3mGre9d8iV6uYCEXC0FMBhzwYpQykpbw99WQVnWFSSWviAETNlFEp2K0pQI3
sowGkhmZd1NRhynW+54qFFeWmdFvog2fZsQFIVXU0HPckzeIutgAVJITRDYiP0nSzvJnryNH6MOx
ky2dC6dNO5T8kCUVWM8BEgiPd+3UUmzMbPwLIDzlyNu+Hhm/oboxhI5EWxVSRlXXG1mtsCLPOoZo
FxUj3BKFzqKcUm0PATITeru84hPfnD2nEE031B82HBbiJK52LZB3SktP2dH338IN/btgu0SA/VVS
9iGerJp1hey6jqt85DkkbwNKYBEUR2PPDW+jEGNJxeFpNupmaQZeoOSY6NLSYC/jhLCRdz/bKxdo
5vzO4AR9ahjH5EHR2C8Ts0aZQiW3dlDgQfxPtbXd5cE9DLec/Wj59PMgP84ohoKamGzPuWaMtK/X
4Wn6C/cdf+AOR6xPpN5Lq6i2U32ILvh3ZlwaOi++8m9A0qMKNdnPwZza3VhMBAqzrpuwwcmTcEuY
pBgBGY7rrNxZciBsw270SnV8Ofycwqe6mm+NmStNBqBFnPuxxwgZnCFLj33FXCO7VyvxnKYFGVrg
LUUb6cW1E2zS7aQzku054lwyliD3GYAmxOvcPMvpW8MA+fSu/yglH9NlzuA1OHCZkCpO9vnWB9uT
fOZxbVHHUsKcwBP4o4vWfkooq1e5fTTKsr4D3jvAP0b9hmT7VeHZ4AxMxNQLWcLrX3E/lR5FG5C8
DzWiCJJpXyVICxrZdZtvsUvYBaYQA4M706dwWk2Uaalf277Ga/YilS6guNSeqt/L39cKz24tl980
hs69lozX4pV+/GrDhnPvcOvJmQZly2CTsIDLQGy/ISmtslxyYE6ErSk+6UXkW7OGSUZZsDtCd1d+
U3PKDNysVbk5yGTUz9rkHlAHAqzj+gIJnrWkEnvtyF3rlxgR96Vt5kRXr6dNwAficJC0T9m3hyGl
RzfeDWYUfOxElN/qTtduWnz1GBykqupQhMkJJNsMiOo8BAuaL9lEvNrvmEF2y7QUqU/x2KbLBrJB
D4N4c5m/UFAK5e20Ace/kxfRH87OmFoOCKHqZTxAfztmx9nZ7J6rbvJY38ML7DPURcBZPsaID9Qu
LQ8S/Eq58z3EDLmMu+qd4vQQ21HVbSY2UXAs7WLmtLOQX3ze0jIvBnWxXNiSCaR8ImPTklh7WWDi
u8rqX/CuKCB+soKdKWQpy1YB0JPdcEtZ0lGHZRfIxFZ/OEGsQIXLv6qt+ManrmtSt4NxrAQFkmUs
koytHfl8ZiwjXmuwr0vctSTPYLqxHO1ZpJUEr82Cmi6AP3VyMIyVXj0VkhWpPv3BMHzKD8c/nSM4
mLebQl36m1eQS9vi0isOc36IwBmYGjRnSHAfMJM72Gf5Tv/ZO0qokeLgaSk74mv/ss/7WSPl6BwN
6escENMCU31vA+hys7H/zC65LrxjB+6d+B/eEI46FbkR1Ci9n0yONyawOeea5ZvdkEfcBuvuswom
ECyqEFHdiYEAIhPuGkizPsNJzhBaha3ppRnHAFCzmbeqNeqJ6zdBBb2JvWc5lS/PpzKMueMI2y9M
ZyPHl4e0lv2xK2Owo+qaTfWZ4hAPvRjBbG8t/H+vICxRfkfWf3zgUcj1sqEGFWAGp3kguKaot32s
Ri71S5EAWM0dBFmuTLjbu3Sj2X/03Gh1FSnSYXC2OEow11Qg/TKeW7SJ7e77/XNvw2FBfrYJLj1t
GVQwOFokFk0GTCOIeGnDGciiqgswdborK0Er8RXWfhYEid0UB1o6LPijOlCRXIe7dDylo1gD7Lme
eR5jj/IFy8b/sZuugPLLX6mjVHhGrX/d3tPaqmiNhRj8mg2hbpCp6mwdfkL9EieB5yyxVG1zAFOU
x+bX0XqZ831NqieJqIUs2MW+QRi8QFxLQsbN3UADTEOv13I6qDfomD+hd8euqjIe9otqkXUrjr3N
fpKK93G7slAEqDqTfaqN8BT8/OP71gF9PCc51QEJ9+YGhw98pSBJvQfHI8toQJIuEW0IxDBLDbFX
HrC/eOhOyvX9TMX3k5oBp8oLXXE/6tDeWwS9E5HaXBwcsvgHpoEnw2xJF4wZCxH6W2ahttRy140N
ay8iPCiag//atJ7Md65Zz/ssnobvTN7HLZ/qm2VeOayP81u4BeB2BPowq+ktn42PonqYPN8sV4b+
ZqkGLhc+ny9IrOblaw0QAhwDsOP9SxT52sRseDg9Vum6uGWfqD1C85kPSx99nOxoLMKHusfK2pBF
D8bLd+QGOVfjp5+ERfHx9nDwi5NZLt90ossTfEdRnVCjus25ziiLdGrSAhThpBgDr0FSvkrXUQ73
gUhGEZU14QNRNps7ebjAXaHV9nglxuKUi+dmM0WEcCRFY6337zT6JW8lASOsEEExJCUmDcHPOk0B
bXU16fKSioblTdRXYl/wG4FJNTEwU2wlic3aKsMvYLqkIpI9z65lEjW16eMHSI7Nn94uqGLAozMW
zk90ThMQE59s11aCcvIwTHb0XWGcGrAaycHM92MO5kktPaypIiYsU0hhMdVp6Kvy28Sx+ONrFEOu
4fHDBwXTI9ud+SUdvtGZkIRfEpnIR8oPEOSaHrEsYsAgduiS+r8mI99V9f/KqS/4thjP7NsrpK6F
YemimdkanCxSqdI5/RYQ9RibShAMf8p/hVW4VE2jBAPXJt+VTID69zS0uyW0MzC1eIfbx4KmpYQ7
frnuVAoP4Aq3Lv4PCw+p9ZO5At7Ugty+hOF3+CbQ3NeTz4cdIDVgG7di1CT8tMJVo4oMHJdHiqC0
L9TSp4ZHGoDQA+yHTibxFlAvAsWKu9auJiOSdvRY/+kTMgzqO3B9TqccAPRnV/UYSVp/J3NLDKRt
H5mlLAUpQkNyw1ZlDIvfwxz6esuxE1ZHuw5ReQvGaMe7xZQvApx52hE1TwSN/FZXa+4SqG7YOBe4
qSiYqZrlFrLCYcOKQSTwhc4LhITj6nTwritaGxuwuOjyR3IaFTZ7qrEKWHl/qrZP0y9pxNYmUihK
oF04ue2ooEV11k90ocwJWBaYc2PBk1MogqzPv0gQc4gqbTs9fPk1aCQxew51M+amKHn/xRDfVQLi
ECEGLiOxSliTANmtQ2Z1d6HNk0eRcvJSVUbRAaAfMGNNKGfArTqfb1afLBLmr1Z3hbfCb3uuUFho
L26JizhhI6QTtNBJKCvIddBzWafHojEXtloscy7eN3lxRBr0eLoTiE7vdou+qgDOzRKpYoaLZni6
JIpdCgSQJpNwJXA/WHBQRQaR7QsNoMuHh7d+hj9qdYb7Gogr0Plgt9JNkdLLqvRj979tvhailNwx
ppX6uKWTRsQZXz0S/MPHAh4g1tWmBMVixvy2YTuwC6OQMhgLdlJwTyNYuGnLbwgQii4oWXU4fz1f
Utmv8/Boj/IrkVrdMyZTrhkSkBxVjP/qpOu8pHTOsqtgf4gu0VVA16Ap94bZNrQDOWS3zZNM/yXZ
SaJkn3vmWj8QViLCU/eTjhCMUlu2emy6mJvt/9oyZSTFPCRMGCDV+aGGcXm9vIcWlhiunwm8cAeH
SpxwVh7cNtiIQvZ9V0Elvn+oZTpX3YWhDm1TqkNOfkIiHC0lFwLrXxR497M7TBa0dCBCFka0WpZq
J2/yfK4DTpZfljl/EFZInIlvYxRfYmjTbvZDLKdecTi4eC2LarayvEXnAuJ0yc6fGcK5/HeozeGz
mBPyDpfWkxCzHLlKLg+E1KNjwhxDN2PJL1VmMpfrnwlGLA90/82lguZmgmRXxxORw+WOsv1yfsdL
Lt78eCRwJy6X2oGPzElx7Ts5pYLw+KjXR/bocxCSE9SW8scFbcX55Ar9GNA6f73+EHZZ1Vo8UaS9
NO5SckK3OdgXHVB2az1bE4L9yUp+A5Ex4sURxuFLpMEvbHsMLfea3xwmDOcUnK4wo/D1NGFtRJwX
BoMMkwLQwadfp0OQkBN3lp9sTqi4OLA0FUG8dosto7Yppq5q3v/l5FduL1w0XIlTC854JXFCYTOU
RGsRiS8ntOs5WvZHnKwcyQGWbQU5wltChVJzDzeJ6utpTR2tPomkS9kYHWuN0wW1C1bvo6eY2NEi
wL2kEjee9y2c4fPP4csLulq9zHHBqQZa+U0dbkxlKlfDuJTPa4KG2eOxrqZvsQoXjSHaUf5fPCvY
r5Adi0NavCRKu14Rey1RolIZ01JPpCn7raD65TAEvFBjDBMi3IhOQSF1DRH3kI7guBg1utthmTAP
qIPwtZiTYs4rPyeII7Qge2i69fTGuyGL21Mq1CNRfaZXhoNTqfjdJ8ByKc9gfx44CvmOn6IwDxeN
3dKPBu9AR8W17VwCdv8+Z5Vn13pmkL381rqKskFS+VasdQh35d2rCWDsTS+5riRFWqxZompZ3Ppe
aoWK6TCWTY/iCDO8B0SGJPLt9rnixDaykm4Ftv6b3Ne9k2f85Zev/NcvZih4srl8myK70ItTMz8r
juLprOKbTGRzSUOYLqHEHnAl1RuaJRTVN67SJNSO9osmGz61pOvVyX66RH2goIx+avylLtvhCoNg
pC0zcweP1ZcO3h823FyLGfIcEsWkOi+lXFm8qX+oNc5HhTskgkIZqxemuLn2NzmW6NCCYYJpy6NJ
p4Q6iXRhro3GR2H/JK04icek13EbqNFjc0UG9FbrMDOogVTA96pYA4iSBLADOf+QQ70SG6uzHETV
rToVrPaHbDeTEb8I6RG9oF04ZLKyAIEoXTKD+uLBhDBifmVMgJIRzHx0ncySKUC0ET59/6W+l0Ty
F5ZM1VtB34WTxnBYHl6xfhZBO33ZhZDtWQp6L1DH8qkwC1BmSE3QciKEgnMVGcAsF2I+xJTUXQMZ
H64wgnDR1U42sAfu0uAe+FJOvUJbB7j7Cdp9f5D+DWKoZSEsWNQ86GiTBYPLU6yFmgd+a6FDoQ41
lvL0TjVVyU1cmTeeT9554EjRg7EpoKvBeZriTraYgqJpv31B5+R+ndb+Nbs001Y/XKqQoI5BhzfQ
jofbdIIkC8CulSH7p5pvYmUQ7Tzr/biL4Ru5anuC/EJUlbGiLrtWpGdLeylxfvO87kauC5IwYrei
Bx/GgkE3OqqRAAAd7HmWqwRxKl19dJcjMK0eKBkqcIjqjyAGRH5477QRwDjURuXAYxMrLvCoJIbL
21ftfBF+0k69Ivnf+JQa7gQ/FwEDMdGDkI5A7wy+hA6hJbH+Fl6nJy7T3Dw8wbLY/d+6uubGnlr5
zyLedhLUZW6yhie/GPQv2qKafOInS4/Uh/Co/N5iUPPTCjGvlShEQ/308uCf5L9mfmsDp1mv4a+W
u/ZMJPwweedTVwLHW9Jj7mF6InqSRRmlWpC/vA8/7ao9r2Z+vasNDOpzMaeDzvO9nkUMGnbna1Vu
BPTCaXyDucGMm7gy3/X5Dn6HWMCeR+Gylbb9FlUXDwov1ZXsmMM2z3DJPIfpIpFcbbcXHKiMcQtU
BP3CpVVOUKBntSbEIMfhhBfKtO2znrJS9s9h/aa9QpSeMLpgY850lZkr2jcGqCeuMmblnKKsOSye
q+2I9mnU/E08zvJA8NRbI6LsfIkeah7V3jf4a+T12opMCZgk1ngDQAxjHs34C0dLQwJZvkqxjyzg
8GIcv2gJ5shSrJZZvKgWmgsgVnCQJZrVSBvwh3T2wYs1aabeCmnbf11qoH3payskrqxxVrRB/YFO
8OIDWWz2GL/aWGJVmcPA/DwJI0PP8j+09AnbyJkgSJnhxQmMKSfhRTX348HZ9QoygKz7OyeaW4rd
S85GcRwE8v7KBaE+ak5QieL00uYkDvVF/unQMsCA9duXQNF1t9OMxb5cab3cDHOZEa05Y0ig6y2J
K7ITdKl7lxfxEn65JGHT4bSRv7bRboJQtmLf1ag/WB9m3nGu60JYQ4arvBt8TGsPZig+DWtfT7Qn
OmQXvWig8vjg9hcHYeChfPssSa1/+9bC+L4gMggvHQNU+XNeJ2eeCmEgxYnVkX414lidlG2SdFVv
cecFSgftw5bA8WP2kMUZH5ION/9FjZ476awPv8PGvMMy1zU/AnIyQKzztfnCMrgaOh59kC+jf2hu
jJ3SOqttziSoLTG5px1Xyi7pLb+Ku9kW8rJBvj0vsuMAzpsKs0V8xeBVpxJGamQ+msTJRR8W+l4/
MedJVxyzgENyjh2fgES1H4pdThvjB1Lf5iCneakkYDJZGslFpRlLQh02P7AOUodbM6U8OvJRmdrZ
D1+7Ix7AGL74SwPLGewdfReq19v7pyDide4petjcmWjFbBKWeKaI5kQoQFzRKz7s8pb1PZzAmjOe
BI6zmn6sqtWh8stx19LEvfRglRcqv2XsV+Hx1DmM0yjzFuTi30uqE9j4HbBupEl9ba7A8MCEMKye
ft14exj0TAwgRSnHg2ZOtb2ceLcK8Syoj/hkpxArT4WQBHLbhb/UFg+6dUA8DNLsAYxq7MjkrJvp
D5ujJwWeaBahOF7Qs9hrKky5bhasg3dgJTlO1b+1ERHzHT71kiPVUJXahB0w9J7yxdpTZH/38W15
F8gQknWOc9zXRzvqrHLU2EX33nxtDxQDHK6/byH+6KmfcbUosrNYMXVb6fdMaNwwfsgdTI0mA4r1
YBVcpbO/PqpAYZQin6DIxleW59gRaHwPYPZo2LMZwa4cy5kmKf/pySx5K0obVZ4lPYpkAKDXwQLR
oDuhvEU2ljXjpA08f75XvcQRXIacF5QJNN2H1ev8k64aavB0hm1mos2lXf/ih8Jgq6M7fGxslqLB
eKouIApMOruYUJQB6kZIAuu4jqOXD5y7dAbguBQwyh8tsUz0QoOPVpCjVmaK4wUGroD8lZ1lETNv
J/gFS9hYBfZydwPsoIJK4Ig/iuL/J7sw3fh3eilkdG1sU2XADQx6khQiz7eC7GiH06E8y26ceZRd
7+nq0MRrEC/Q4Yj7CoUZDR0MBLLOyBSysz19p+xDLqjp9c9EnA482ZTbTIYdUlRfKT2Xri5I9LD+
PcVivN9wXTBgWNPv3sTbgoW5feJjUUZrNZM8bHMA0EfZqBkDimDpMhtkgtavKR4l5Q2mjoj775u4
EfAeld5u7obV97LHgopWs3lcfhP16C2t8glR9zlJmGA5+x5VdhkYSp5GiY/Ox6rfW/uQI4pxBLYU
8dFUmZc0CgwXwmwXREjlrBCiEB4kUlvnmal1teMmRvN5OVxwxN1SI0HcwpeZnKGddUFzuT0qwHjR
4DeuilJP9kMjHcEbUfBW2g3mrn4EoicEHyaZcPt6qg0b7dL8eqUCnhHDFNSAeHD0Xx/eLGwM9IPv
di3rGzQOLjKsDe1r9KW+HrAjpi1RYd42NMUF0DD+xKs3luASgsgtuFHbksrkaJdUl3S/1KSw2xhs
urkEMuEm69Be6oGMMbFt6EkQ48IXFaYsgp+csAph1ky2T8wdfHkyHM8KBro6qROdhzeNEJFk2vBs
rFkClErsWz4qCX7eJmI6RGXhr27JrGblf/kFWcaASyMS+txXXV/vJPZE1/IJAs6CXBlfavFgQEL6
zXStzP1DjoO6pkEKNWb0TtNaWM2r/KR4Ud/KEe7ZukByCzAZtvD20iRTh+KsaMH8wMw9ZKCQWZHm
2zxopszOBuuFH6tHHgbEVyy/2UVY8dc6/WcmgiQM7bsWC03W89DwQCWR6Nxt3M45Kz8Frb3QozyC
pOrABqtTJ+PW1yI9y5wKmHrYb4HI2xCQuwyvYN9JTLvvL3okZUEgzmn3z2cmM3jWSl4X0jtlf3uM
LYuYhbi/aT3/TMEKShGvuCRf5eyFSvaMNHEtFXQXp1XiXqP1Gt0n27I7lCv4Zv4QezSG+DnxOpv/
tMJRpS95l9d4nQFOkOMl5HtW+c9sHesNJEJ2JqrFssk862wKMn1kV4DPMPm5h83F3TdlgDOdzD7/
R14NUjm8l45mWldqVwSfg8TTNKaTlHYUsFA4WfoNuRtEo3+58g9vBXOni2prkIiMGpQiXKJ6xBXm
hfdCoUDoxp8FTWrxuFahwgYtuM46HjHWJmpRKF60c6tB6z/aXDKA76d5IZX0aaGPDWyLdfhFWBDK
tUusAXpwQhmtgP/G0MxASJoLlWuMyXOYTxmmpH2frXmVOYDyuRqpCIbFHB6Bj6akEfSkcf7GQRb4
MAGHasDBhmye3SvKtzC6xUE73JZFMnxnYdGOPxZSLoahx8qF0puyv6PBT8ezKUsZ+2R9NYhetqil
GltXq8ejQpmZTs0eNT0b8/eVk+lLzuz+3zctcIVCFwb0libYGqOPRnuK6DPtoI4EF0HNf4Cbeoqd
9nDnZIrkX98VFwBqc38gf7Lu756iK5TGy8UlE9Rr32A8GQRrcuKeC/FJDcKlkD/dwFk3g1XeZaSC
jzR/d7A6wIyKo4G7IwAqi6Pf/IMfSEmaxDSqRCtH1BMBJLkKlSXAHQPPaxIg/nsmJ6aaM/7EpkDa
XNPF+NCluNZo0UBXlP1BiPP3k1VUsnumKRMW+fcFTBzAcMPcHh/yLCYy4KuA7rUSzJWUOgpWpcLR
jyOavrckx3iF/j/TzMFItZpa8PDbmK4sUdktW3dmveu7g4h2sSUX5/+YjH966tRnxbacCcOfTEES
tJgGDUuLUvR94PpLZ2uYKjfHeeHsMKaczY9zAaRdT1WKkrrfqwOarGWtHxnWZCzQnSfUyXJ0miFm
nB2SpS/BuZsNok9HilRLOG7+QtkkHRfF/X1p8fTU5XkMaVH5132rcLk0dqgPv1XeA7MXU+i8m8f2
0iwzEZeY2WzIjeF+HdwpjKlVSH3Kfcpd29Or7+c9bi0PPaMnVKagMV5pMgWDcRFs2EXvW7I4H4Ja
9IVXHeYVnhD/kCW+HYuH4e4l6eaDSv2jPmbd8m128mpKF+vBSdWroqOTzTc1zfFODJtJtfNKRjjF
nw0ukJ1OA46NPYpNNr+axkjgJwvTITzGKueNdwxuUAc9mVuCEhX945vCnw4V7d5WK1DSPnVetEk7
8uK6/kS6uNhl+EZMeH6WqLx/dPRNeXAX2xNYsqABiTHEFOORyEqgngagDQnlqZnQGcxSAsEHGWSV
bjQJgz+JGJLu4XFTE3DqkWskr+KAYWHYCa5kvdqVHvXQksi39IMDSVCmJRNHUBJW5/lODvnFmJsa
3mc+tYNXPWl4ruvqIwSebmQkFQ2SY8LD6d2Ek/eC13IuKw0FrERcRx+nsRoyVFxCzS0BQihl3oR4
MLAjmF+xeLQR8w6KMfKCjyElUwO1ABYFBE2eL6jHosytOjd8zEPvWDsBfT3NSgzvGeNkSoNvIpwe
ETr17Ahf7LEI1liiP9HAAxOGM1lxDWhfMWHFIhyoJ1P0NWCU020C1o/KaVHYTY1dZZ0J3fmXdJFn
37LOP9QwHdi7w1bnctAyKwLgZA6luEqTc60PKpmzaFbQO/DZIOFAr/JhdDo3xE5wnBfM6dvdQkpr
abO7oKrkrITyS6g7GvwZKpVrbvo0mQt2dUxmtlZMI9+rN4ix7rBcHBxlKKaV7Lq3BB7kP/nVNWp3
4CqiN/OwHpjmp4ITcsRMgb8kb9KZMZ3N1bG4jdYVH7rWZ4UtiLmVoIlCminGqu0BgeSpZeFFSWeF
OjMDcD82CumUBut8y2CuQzUm/W5JV7QAScYMxqbvMvC9ZZI4M2YR37MSXMx7xASoF1BGW7ytuQ/9
4NJ7QUu6bMLD0x6czdNQhI0Kr4q6iwNfVgWlTNQyr1KFy9J5beXbljZwd/ZpZ0EXxvNOiO0U+LR8
82DJNIXqqyF0mpj6ZNuWx+Iw97486VI1KHtYUNeDHBRfPm/IyxjCI8D2qGCRhq+8I/x+OzrfSEEL
leNjfxnQUuwlJuIE55X1lYRnfH/1t1uf9W8Iom7XUW1nindNUgNeo9WrqKRQ+tf7j6Cj9/TrXCiq
zXk/e16mVac52uJxT2+rhztdFjETKtg47wHk9WEZUtGFiZe6Q1vAUZQDvcdzBskBGSMAUxQmKaYp
ImAqyTsI1NvrpAzFMeD0nh+wl+LSL7ykE1I9P2SkPplEwU1D0yVTjM1Dqf7z2YLWq47Vckx8Oiyq
XbFavOfavR9WL+9PMc7PXlHo6e7ClbYQjR8cUPi44KMQOJKujd/CLybkwmf6MQMlj+PCwiNGrhn8
bmTcZtGYKT900KKXXkYu4WDeQ4l3CEVJo3WM+nAbomSuzVfvl7go5hx64Iri690IHBr5aX8BGNnI
D/OIMV+Z4QVQLvo2PrVlwF9PyDIYgfCTiewZ4X1miDpED/+bXSjnhg711+VJ58HU3civfT9BJbAc
yrXn+2OqtZ3X+hlk4TyElS3usje9KH2Ty9XX2y0aaZmiWef3rLx6qpzPi8c8HEmp3Mgfw7+4nH9P
jNtD5PyNAIPBLhcbpLJ06ERfxgjhFLvTzHIJ5dJUYD5kVc/y2El9wg6maGAM2BD0vQ+l2RzYa+s7
2gheCKzMJKMIw3jR0CpxwY6Jh86XNhheR7F7Du0f3O6gYZzLwk7TXon/KfdmgXNIGRz086dp8voM
bdYNrAQuw/1heQuTtvNapI+Jyzv13rRxZYTBU9CfaXyfNJt1NaVt9gpmXF6G7buNv60AZPC9x365
vtujERcNzOBDHkJw3SmW6j7HPkDDEMPVt7L8nUQgqf0cAzdwpYY2MO9EmWzvzZqsGVLvX3uUhPbz
Oqow+SH7dmzMdTtxLcupurZIL5UTYEAW4JroQOgKPS5pApfqDzMcVFOfWCxNictKxyRvuT6idXL7
9U/sHoOSebvd7CXDGEoDpVcMGm4Ocy72MTD6/WPhip65lSPYjQAFHDDxx3C91N3cKPAfAPWJyJtz
J3BoO4VkChxvQLaOmrSUEPWOyNueNzEEoS1izGJoXTxeqLNGqRHnU6DU9UNiaqSOz+yq7njOhDYh
2yR4kVki0YYPzOlMIhokbaY3MFO3smmjj6bz/OfyhRLw1YBE6mAfpoukyRcG/qJ4FOk2184ougQH
CW47hRKiVwNyqiPCNI4GvzFkke0oW78h7A57PCCMnmHH8nXNQiNZVqq22PBz10dGLQ4lIUlvdTMy
DJU7jEWheITck2mAMWRJFQAkKRyX8QCZqOaKl1/AWPzKBFoSkCWIAAIH1sHS3Z1M0wHwmpcKFa1v
/Bw/v0/7ItO1PsLz/YuieSKSQB8UExb+PUs5HsiE3UXxl0ZKkgJGX+YZM2V5LULlYHQmdxwPexkK
i0G8EvAUquDvkl6JDETdtlgC3mLkqxDM/Ac43YIRiMi5xnqMIah6m8Lymk+KUTnmo1UQrNgV944V
RL4x09t4VjYFjGyMJM4qlvf2xJwHOUgXGqU11/aN4SEAv7BIXF3BAvd/q1Ska2ZSL81XksFSDAuF
hJGrh4CYgPL5xvnhrfLtun1M/Z9O9sweSJ8Bq1euBdgF4iDvU7vaGepXb8TGiTSKWL1Osht1VzxJ
UA6BGBNQlClE0zo548OtCuSragxPUZ0+UTmk00uf0Ny5dRJIuSCOAPxzwe20biRcjSdG7sUhRT0H
3B8PPGc1Lh2XGl1yIDj63mY1kojJbWbDfBj3CdrihMEp14UuPSI0+caBLWD3ErLDAuuFCfAqNLbg
DZ9zSASgwT1F6pXuwLUMjz3ulp6K/pAEKEpa2ho6jZhq5it5G+XedlNGBujLee79yUE/NPRrX+Hw
HRWexF5F01Uh+fykDBqUYV1AsaEYw+hRoSM6g/WZAUIr+4z3wgEGDAK+G2ToyikoC4QEwhm1Hi/q
pzSKnCbSHwePcu1qwf2MhZCSvEBgjkPQB5i5JZfTXrrOfTxJVNmHXxE9sfh4dtd7lzjQMjHK/HEX
GUrqcoB7wa3oNylok902d3Bn6ND2fqUQJE5d7QKPzz3VrdhizZPsl6erhExSykIqm9BuH/u4GmEH
IpYsN/VuZ/sr+Sm3mavkbTwMa4f1QYoeTJuLGtsJsN/2Pi0212OjCI5MzAzkwS8nVb+phWA1RXTK
nL/Dr3+lvG00Cao8k8+jITFUL+Vad0VfSFkXkWu79O//u4KIEWpHJPaCjBiBU55hHkw9XzjahmdV
kp53DsJMKtDMcJchKW06NuhrpqOs3Ua2LbEFOcjGbrJcEdjSo9wRE3N5SrZxrYvDrsPzHbNdCBQQ
osOsukDXLqGwyQ4377Ho3yR0L1f/3Hf8t3sd1MvxpYZH7UBvwBuWFx5lkjgWUtbT7WnMtKfvbTqb
hpIO5TmAmp364TIgvBTD5nE3dCdgflXfyru1F4xifehHP/68ogQoiKOnJJEn1lYPfsaTa3j4kTzo
7jkZA2ZSCoEWURcWCCxK2SAVC4eV68F8F6SVvLUeHDNCZ+08rxLA7tVfk0M3Rn4ZwK3IJY/jnAML
NYyOwdcid29L+8kfTYi5XrQqWsGkdPHfkD0wHfL20KzX4xZzUwg3q1bqKRjRk2jaVpL33QZ8Vf0L
KUoIjOwieubjxVNSfLK0+fboBo3fqYRXtd2QXD4Pz4MsmrUtRcN9qJY5P2nqKim47Sb2Wz3BLn7d
XnXMj96H8F5FvhOmCIBAfO+UjE2Nq5Vk+veEq1mSoLIT/igdVLTLjvsPfs5gntu+e5Oz19n1Z8eA
IUZGUUSgca80Ilizlq13iz6K9NPlQxAgtuH6ZOUfRCD0RAivAp+NMhfU+/SYUPCxekJ76jeHL3PJ
GEs8q0LJNa8Oaff2sV8EsI0SB6uEIQHzq6bdWSQyTk5LzMCBqnIBdp9zlLlMl41rcDflgHwfgpdO
cFNdfemNYGOmHDV83aQY9ScWMHEQ1AJ+JiF+b/NXKRuibCEMGTTuR04NgWX0peHwy8F09o8aKZSS
nwSfcwUzEDaB2NTmFtl5IcQMqIMnQqTLEAYK0cb1Pfm5NPR6pOTIrHLatxGvxTWjDOrGNqZGS/6x
/YGs0DP0NjIGAkKDoztGeDirbRiUvqvavceQ5ZJFgPgXQscuDBn7jBonxd6pnpE0DX7KtB7t/6kF
GFvPrUejl/k3f2EWkhXJHJRYCGhTAFAjKvJxRzSppkaSThyjVO76Z66rVYJuPQLBVwwwC6uH/DQy
POGGtfdn/bwSMBqxmmiU7R9dci7gD4iANuo0WWklIMK3lvZKRg1H772NF/qTTdZaM0ppWCi9uCsG
lgh6n6/S7lGPlDssKxBP8J226o3pHEKar8CaXW3KyrGNVDmYsCp6a1eJBmDkeVr91hJi3OSgsuVj
uA4lsJLvfa14LaXYbxYgVrOy/uvlqF8DzY4bZ1hT5lYa4gUyGL5UvSz6oFZnk825OGXPO905l/Vn
1PmY7cw0hhUHDQGLSHHbiy1XJoqJHCPaxHFD2mINEDn73ukQnIXOfAHQC8IhcoCs9wAZach0G3Yt
YCWcwcYplO/lSnqo0JsQZlKW0tCKGESGJhr7O9iw5F2moPYgheBFCZpFLYvFOVKkhV6UWEDQwBod
Wz97aPrLJQhEYBLH9L2SsVEi+m/w5/6v1QGL0muKYncpjLn0ld+s7mXOFMAl7Mzz6l1rouPVEilT
aTITuoXgZWjJJv1qPwwTkJB/7MTN345PlqCjpqwD2hJm0ZVdH5GrFbmawwGUmBOuqOWKsiDcypTv
GuEB1Z4T1Ml6/2CkNkHaHPD0lKEEVP3W3hvejTRLQRyOLzfoX+Qy0kVVznNleVmvYloHgLCojeXu
L9hBhrN0hGOrFsNj3sxFuU98DnBqQdeI2xW0baFFUqBwzyFFg+snTNyUzsNpcohW5WNf89bJz39t
PiVsN8/UnrXIz6zN8fH7pyzgWZXPZI9R++0SmUCn8NBrzsEqjF0lmMnQl9EMpyFmq4FySHufyrOO
8EjQ6FSFDK/UsxLrDoNcmaliM2pUm+nObQpXKELx5S8iY9cO1/85TpcC/L3c6SrZbYkUVyrU9f3U
3stYAqi17ORaGL+7fr3j/ci6DVLUqy7RyO35YHVMKF/H3y+sBaAMEFuvo9AEqJTaVbplNsy+kQkj
lGbnmntRksPUokjW5QCIL/EveSvIXfyuJO4Om4hkGFOAi6ypS2JnemndXOMH717tZtYL1eYIcrKi
FnVVi9tX925eGajY8qEWGXGZCP2uKM/iJM2qOfD22APGpTRCF9YFYxBlvkfH6HtwVi1oGNJ7B0eO
WdwGzYLUrOx4kp6k9XQZhw/feghnjWwxlsmmtGwoJuTScIq1E7ydt017jgroxAId7tvqO2mZqiof
qjBRq0Ld3IQk7MjGgUtYjlCSO2qakRE5jhkWbuhD7e6iib2z/37nLL8hSehWoq7hXITSosdDMH3o
bDnrNizDbPcwbvq4p8DAa8aFKRSEsodWKBCpf1xxkOiVcZx+xkIevsjQJnxSfirB3kkIQ9R0Si2+
taSccauhLJL2bwwZl712PoR8c5Nzwg9vVDCcCvqrJConSQQOAieNC67GMURk4VEkVTajpOQZAt9Y
couAI/55R3hjVPrRaa4aW1MQvITBRHq6cVl7QQnmxiHYw/i6fi0iO8VSm9wgMiGeSaAWmLd+4rMK
H9o0gDXxYenZhSt3ZOA8zhEjF340jg2WaLRPlEdmJvOPL6xZ3Pzg9+StLyg6erenOEAK6P0bi2eb
FC3e3PWmId9tSBIjj6gl8OVJi9id5mNeCx04ZTw55VRxeuracMjdO55Z5fSG11h+WvzK+WCodFad
5d1DjC5ySYYBNYS8fORhatJbMLBsL7zBZQkaZbMp2RqrKv9bTQXXzq0VMK/LYpJxzhtFfdvWpv00
KyEU15+IdphYHakkVuE3bu6GtRlyOEwN5mVEs65VVIwq6+75fvmDspGMJJ6ZwV7EWMFUBnEZItcP
TdRtNrahlCpk4fdZ2/lcjgOHw6/jOZKhjGe1UqqZwZ0TwVB/VD9YPNqQuW1ucTzF/S1gog9t02HI
QcEq6gUKBjd+niiEZzRc1b8mNhH5xlcmGOkid/DuVuy13mzSbj8y5tAliVIQ2tgrlGrjiN3Hprz+
4mYrdaEpOihed83iLqChRklJbrSxuyAwsXyh5wQ+J2Zp5JjTK4DzaqNGSFv8BLOo2HpzmYYQuLNj
ZdbkZsKCQLdWResa7SOT2XW80b+rl66d+VrL5EXnDEeCqsi6fezrxva1NfxgGuLkvfUz0KOvbs7A
HdJOQJqU3P1qTqT3ywHWrjhckkEyDZWL1J3rvtIKAGyXQkeRMf43GGewIkelmJEjz1mZ+eITPYPA
4D/jC7ckdjnkJdDgkT8nr2ODVoFxqLHuHTWUMUIbfExduVQMNEOzst+uWdbqptJDy+xoMwwNzkVh
9wuIoRojfvuYRfzodiHQHl4VkKXjCEykmF91zwfHa4KqQ6ljfn0LByySXuCjMZOtTi591lDshWZr
uL5Pq6zocziY7tKGMn1q+M7fGZZFfNqvXQdxk6RJT6c27JyU5kOsBgkDrJ3Lf6BXhkRyKjYAVFuh
pMMrIy7v0Nc/X1l8sLfMNEPHv2FmPb7Nc9uTPHgBHLBsjzbZMXo9qGJN7GENWGKSU1sk6OJyMTII
SqfWRB6jCr2OhkHd5qz+okJFZy01j9+va0TEMAV8zOprZzK6gIOdUGqaBbLgFcEQ0m3M/lukoxP8
IEMUzJLdk/wWFa2mCprl1R7uVB+0FCppceSaGAYMCDh39BBqZOHOMUl6QRSbzTzaJXtkiMP4dnVG
5QWTAtOaZi4D2s8HO7fFISDW1Wh99D7Acfg8bKXVS0v+ng/lHsUI6cF4wBRxj/AQ0j76Rrva9PF2
jqa7eVHz3zh+46WcfaTZc4lz/p5Wu88/Z1QuozDSqVBRr7mqypUnF4QClzkIygxFjnQ1QPeGQFxq
aRmG5M/RcfLDiQo7aCuhkUs5q2yV7EX5Im2e5nGDjBaCy3glVtXeHnrjI/KwHG58SAEwAxH5ytTk
E61CwHpWLEwucMITWUJzphS6CdfCVwADaFrF9W1XNEL8ploNTwHzxT0Vn7TIShItCbvMHUcdd0c4
j2bFLIuNztTil6Nsmtxp4HE4nyy+CV/o/nTAC7mXpxOBikYvX7YRv1FDALbQirQ70QRYtQ+6nc1H
4NFp8gnGensY3zpSNz9c0QKHa1+brcpgczpnHxz/dOefZOdiGg+RHzuwyrLCpsqLd7qKkKbdB7xr
r59Hr5B+xJu6eEqqx+ubWG+LsMLZj83r+Iujele21CVNvIJ4LqhD0t47WzITwCkLy4bSb+d3Xq/Y
qotn444Z/MWOtw3mSBfg/JuIv2nNfGDndeZbbd3dqIzqvk3tfKSzopdmTflzkuoWGanPn+FVJCEz
35aKefvcwi+0p6Ii7ViPtlaPylTOmufmh2/HGcuVfNM5uvXe9n/5xfBca3HZglY9RHTeB1cl3fP/
dKwM3bHvInUB5s0W9TK8+JjCIEjHlqbY3FGS1/agVAQW85qnvm1k2/GeSxbjaq9VTj1Slh5Id7as
NkSIP6AexPiYCOqlxTeA9KRNTFc7IT4cW3tA9FmKcLSLnF3BLimGUrb1dZ2vHzvTbGWDa7zfsV7M
a5J3HaC6dyuF2i3kCT9YKMP5RNnFnsYLiKYQJgHiDxP6hfsiLU7rtb/rwyWKxqt4snguQ06XWUcx
oitQqxFRja53JHkXzhBE0U4OFbswVQZKosDwozFVB5d7aVPjLh70Nb2GTdB1j4RrrId8Sx2xtjNS
orDYp99TIBt/bhd8IhJnlYCTQFdMvylpMuhPR7v8DAnue7hxqvLsXXkbVtT/PTBkzYmN1uidN0JR
2ojrSkMNNfX+p0laAxTICW4cFNWiRaKgLZ9Dc2URQBsti410e9PMeJegwHyCtEN4/u2JBADA83FZ
CnfYdaJSIDqqKn49vxs1Sw/YxjsAnUjJZLxkkxKjTQgzK+2tr+H1BVBAn2/6R9Gyh9nlERmwQ0yV
yFU25I8qmNPfUomtPuuurujB/Tpz23JJa4KajMZSAxsAUy8hJncx6VTLH6POYg5hunbBm2EGfvmr
O0SI0xfU5fPrPEwS5mOrJ1x1iwUohGSVuIbYOq0v8wopmp9OOCrpQnURMw/SOMNE4QFdFymX8qsu
Je8BGd27qmMnMF0YYIjYYXpSu0qs5zilohd312u8NWn5we5XkEBt1eDKrpxt1YVXDpew4ZFL6Mss
LF8QQDn4EBEHOj7r9pb+aBvAvNfPDDydrmiCHRAmDYlcg5v+shgr1pH45Kke1X5TLrpWbLilQN6g
TB6q6yZof2+Bn3IweOdDhz7FlLHStWCoCpAfemf6QnX1JGAFJ5OkPfE40oYNCU+/GXWHOM8o4v37
kmAIPg18DjDifB8w9JnVhxJLQSNJCfZabzBHyG9WgPyamVKlkYSwimNu3tMZiV1e+UQHRoFdq9GY
G26TkTg8WLsM6k7yLdKYsouvRomBrJKJQM40Ef/PC8L4fsUvPszA2dJdjhixE+LURBzmpid70fA5
x7GRzfPPaQapRCRnkY0OPL6eR+32mwaLigQwfPtp9scuZzxTeRN/0T1ub2WX4Ju3k0Pu2htwGyIV
KaaadWCe+EFEmxzklCfCf32RNqxiOQP03YNJfX0l5mhInn7w17Ll0qzdn6v8+7bI0J4pNPBrjUX+
XtLl5pLHoGJ0S15LoZD6Hxbe5i7EqbFYgWxfLvuaAmWeC9PT8Qweu8GAwM6kPq4BkMOiGjvBLO4M
g5BpLjU/lrhY15jGFQ4JqOahtqXVkcg5NrW3ZS5QE2IdbiIntnC+cnVhorYc66bVL3qfoR3JNUHM
TOV7AzVRNqlw/gKrQHdZq0bd1U+41XNojG6Av7HUfy1MPFOZ+6uyu26yEf5C2iz7duQ4h6pY94um
6zKYvaqTMztYWmysLXJbeP+3WDqfoxJxysgDmOllz94y0r1yTttiAtd96XwrIFU1zVghdZbNZdII
GFLQTC0Qb/EQMU3ZtkEwtJ1yzdsRxT7orWUlGiYqq41ObMa2wEL7SUE430mPsvuXtFJ9qmGDFCn/
Catbv+U39nHG+1uf+07JMf+1vGDxAz3s15eb2NTqdRWMMF3PMr6oMZdDPIYqMKnO6HuNAZB4TNMV
ui0OpudKRzbVALBEQBzsDX96qO8q/YBgmdAxtliCT8OxKVXRk9/o5GADxakgo5YcaPrR1vnP/YGg
3k1SAUZYVVDw0eYWnB/aajSgPzYqKIXBORYdGmZRqY/wli9d5IswfuacNdG1wXJYpvGPuiXdEfIk
slCBuODBvZmrjv+hmqo9MqJqk48o1lezNJFDq7NdRvy3kxRhxA6eXVd8WcCfRTKvZ+K2I39ybmfL
nUj5hK21zyQWL1RKqSyuH9zH5K0shKV5cxYyZiI9CkuSnpcEtobBqVstSNLI3nVC/dPL22MBXZGU
QPvOIZMzyyS7oZ/mHd6rXdK6aSM0dnKtsD24N64e23NZEL+htZWQ0Fv9sB3lv2n7VeqbiASzOF9R
VZ3c824W+ECsYTgmpMhh5NBSDlHnKkPyG0bKzq3/GfzAjG1W5c2S6tTaNVGKNSEeXUW9JbgehGWL
2DY5g+wZwgig569XDQsz+Fl2yW2Q1ejH8SocPNo97MOmy3A2zCnNo8PSxrGz+FFavqAGQnG2Z8SK
t6pryu5W2vMqTrSHUjLM1rZxyBG7C+7vmngCY96HrBz8QNWYxy86fdlPIbOHYsRQQPOijrMTjs3d
2BBEP+nyhylqAm+u53B1dpnYGCZkcCpJ4DwqefqSm+Cx3nuA3B5CU40cmUjg+wlsOuzx281/TzEA
RD14Ro0nJUw6upSNUbmnfJ4TI4kStVOarUzUyjUOLzZRH8rOgGcxRIUHHMahx9hlwA8yZM4fVPAL
B04jym+7ajGS25EgQRkCfL3kpA3MwZ5e1IM4EM73rSG+4OS+Rapt7niV08Rike1Q0TwZCwajjutD
/RJhY7SLjSweh5wBWLOE5LeqODty+UQTiiY3B4K8SO7YNb1M12jwOHYPnNiq8vs+7uryJDpAAd1I
JlNfv0wC83JAqsbXePT5WuXCRNPBXsc+EGQxZP3yC3Jxy6EZl7NdI65r0o1c33zujuuGD7I3IXva
8O6Pj5XJQi4IpLAW2uiURtAoF54LrcnEERfqmIrGtEIsGLKW6rMQFt3MbFJ7oZsCuELS+Er2EXpo
RAs9ibvSSszEGGUEO+HLQAXPT1Y0X5ssP6ZHeeBInPYkhAvUNeA35AZTrA2Eelq9tuK8uSyMhaFx
HnGssRzHkWLFte7s69ITEIPCN1RkfDO31xSAFejeBpVoXYRH2J9yYor9ilEoRaLo/eI+UC0WdKkv
Eq00xN1ULdL/WTgm2UeqWSu0b+ChdZo1HCg/j7Gi15P4WtvSCFW9QBcEMm/jZEElpZABgXbjoRbR
SV+d8Z8ZSojZm4A96Qi/m4l2/wbIGDR2V41JcEppbmFVA8gECygN/icP+Dl7av+vKzNIslWTEHf9
NhdcJmoXt0/kpwTAc4BxGanz0KoqM+xCJNoQwsMCTapIL+L8x2vTBgw6RpPvO+L7YKZ8uaZKtvYs
P5RLLX9gCFkuapmtSENdPEZtAxoz9wmdpPTy7RtzcrNsRnLy7xLc2Wzwc9qLxcg5cdhGwsNtXv03
boC4XcouQEXPF6nbOu4uXgmVQX+b72WjOnY3UuY794FnN8ESRdzSq1ivwPy996J9hs17K7QUbpuQ
IfMGqbbuGv+79+nT/F7t2kmENHcEFwveInOv7JCamZAg2lKZBHkyBWKKKvss8AAqgwlz2CEkkK4u
xTGrzdNk0Qxu9iYsVXDFDJfCPvFTsdp1boloK68MqR5VzqXi6WCsMsjDvWiRCk1l9YZq3plVlCf+
kzaDscPtsfl1o8sSTxBcirz6m6NEM0Ip77UKxj7f85pkRBBE4tATThw0j4J5YW3/7FNIqsftk4Hz
BYcHOJf08NOfDbxxbE/k4w/fU6VuEfoU3bVbo/UD+ds4q4fXw6+bCm6H9Y5edFDuQMVxsvBkbyEC
EzPRyou7VmIX3dsSJr3s9RHTMRIvqaMYqAT8ibZiTj7JItogEPqcTsghNksI7nvMUTXOopTeSXvH
/Y1X1tXrEhkSh2mzoCcdvzHzODdUbtLE710XovyrefZWZgHQUI40Yg6uqqCTVt30+0TNsCKMQNNz
7qTEIWGGHz08XOvLs/aJYUPvKfErqWbzbo9KbZlgUKpiWX/eVRjvDh9FU1iKnjjdToJJbSQKxQbM
71OBnznVKNkCKVKkZNi/We5g4FLgoA8m3Mb8nuCSQHT/sz2h1Ri3cy5Td0Dsb7fxubPKV15/kyYk
EM/r6SLrAYcDNPL6Omkw6tS1aQw9MqnF0Ie4ICo+tUTiQCKZ0npstkoukSLxqr3EU4wSNvNOZzyb
GDw/Q4G+cWzxbqq3kMWFsM2vrwHYZs7VpZdgEw2vfIsUCerIo78VFnl0B+OBqaRbOJMbr3ulDX8k
GvC1VY6vvdupvC7+dgn8qiwxb5CWU/yZUlM1kgZlGcbab6NAp1YP32zjNdl/6vpjDqVIlB6GZgKz
b3IXwOA8RrVHvv2ubYB3Rrb0GqDnjyn1FINaXsOUSq1WniheMxlayOOD/jaQkbNHgSG7YfefjrWE
LPPPde++43flfdlpqphNKuXtWwksDppoeVeqK5nKwBmAl3R4x817vPIeljbo04nPQxQpbFM0nrow
biFwOLBfSaYzNGxl+h2ymQP5IXEx3mTpAFV6gz7d7b9KLpbRrw+1NHYiYeHJTV1pIQVFYeyTvHih
SA+r/QeMWRKBrgsalyBv6Oowt/zoiuFxpLbI3/PyvaGKkYCGGWdNZkCudys5BGF79/IIFrruXBdI
S2kYZa5rufFViDbiQxq6XxS45onCsgosJjTskZly7RTefRNiUV5ZMNqxr2I7F50g/wQhgfgAlryi
9lr1EwnknQDKn7mmpUO90vFfRdM6nnv1jJCryVWq5vs3NCueu0YkIxi6FT1Kdq8rQQOt05+YCd60
J3UcwI/CtLG1cgc4hj8sDrBB35UhCLATLGvG3IJvjOYf5VpYC+uigQnCO6rUDeO7lNSYgDQ3X4S3
745tsv3aGOALiZqSbAPa+dMeQ7comZquFTQ3REABcfyqCQaq2DjBmzPgb3M75j+5Z07k+Ma0kPbU
R6CzPqnE2ovo1k5YiHPxUSYLBt1g5MQC65wWjDHpk/pdSYk8GYmHaecvxU1/KbG50ldcJCTDE5gX
a9TWIemwfpnVK52tPtOq1i8Wtth43xjvXeKVSy5NTlQ9HUdsUTMd6r/qzzt9OIWk7dNQqBCzcF8G
4Kzvmbjnl71W004xV1yX+l9qeyA7i0EtPuxVaUkeMsZjIol/T70LQDtFdnOEgkvoLPxSGLR9nckO
lxzZHKtLfKocPYfMs0UkVkupKgWHApZJcJAjGQxk/B84k6KYvYdKbwjPypOOfUptPm3qI7ohFBUo
fhvMHzvwtAUIp9Zuxum3QMJ3UdSOnwP3jiyTfWG4APgeqO9nFZRLB7Y8K7+Al1S5nJjcAEuta1Hx
eqP9Hz33agmxesYOOqXAQj+mwW7SaVi71RmZsp1tTBsPtaX+1+N8bTZCSBDgJDmvdlBz+3GOX6kf
hFeQLcg/J2/qrJI2+Og8JL7Aff3bRfjqwMt4QoKnsGJxafTbWrHZZLei6+qO6Jq0rX5bMwCZSvjv
xhK9NN8ZeBbo27pegFyVUVwn5+Kehm/4pyxrdAP74dpDMUOTCKby7tKMRR9HPAFOhS1jBzvRF26Z
pACX1CT3GCX6L0tj2FXVXnrbmc0E5Bxn7lxIeucOLEhSEt/cko5ThTAt5n1zgZRQQhBdusB+QjQ6
ZqxwmodMstnqU0V8rPKH6bl6PrORuy1UgqpR3ouguNkapbj6V2P3tEjLAfLR8D1T+hmjt0MjluKH
hirxAzM+ht3YrK/XrNHg3Jdffl5vs1zirmcHM2f1HiHfkk1xaAYBXx8t5x4smQcDTFoVdKeA5hGN
39EOeVB/lRoPAvItCLEFLZzlnlCJOMfuM7KHWZZ9W3XQfgRiDp82PJU10P8VZ+WMrZjCw5eVYAVR
sH/aYKJD+La3gTFYGMtyttyf4k9E0e3OGLDDNdSFnX/3pqfIf4wVeIA0HB1hjlu1cAZdrDbOQLLq
w25bdkYusF9WJN28fvQDtNnxC5OsKum7wWVm9jiEilU5z9XzbyqeAQdgpiWGGP1K15X7YkL6S/Nx
QTtygoL3UPhlOyQFM+3L6weJFNtGK+vgsVTpD6cBrAjbkWX7RB5t5goqDjghCHM+t6ocoKdawX1d
D7Y9OvFNfUqj+QeR8aamUBJVsLjQmBmrXnI24BVP3OhNMSt2BUkDx/77NUf50Ryr5+YgMHlnPXyC
rb15yTagDej5NsCf7b0F61J3q8NVhLJH+kSQRrktotg15aYrKUDgzIOoa/d8Fx4GB1rMRkpl/GtY
+kWRd+3l8lPKQ1uoU5Vj7Po65P9e139LGrzYB8ojspABYAVqZXiNsovwdElZuZgWC5cD9BpRPJ8I
AszHb7hq7GJLjC/1mH2vubEf7bWA/tiqDuZeak5Gi1rERGLx+jEQDiHb2C2kJVPjOP1vuvEHQeHY
LVuCdZstFkGTZ3fzVu77IBvhIm5XeO4ZBT4k+9GG8+ej/s4/4JTziIjYgbMtLAeAhMJ5uhz94pYX
8lYpX6kvzYykbgm/Js1pQeBz4Fajx66CvUy++5HCTUVLTfsmPVgGzKRkRmFJE+xN3YkauHN4NYL/
HSSFmtMRAy5WkdJmm2uR/a3RjoaifIzekq8p4I6wyR6G6iqTwkyn8gkTstYHyd/eU47py0chiKy7
24gj3BvOffjM/xrCUVyINu3wbmWyI1ACQ6ACFWbwoDQODzO16njegVS+etioB6UNlJw803e5HzRY
NiRoghYLjiTWg/SSMrtWgeltErwMtWEMar+u+RluNUMR3w8sdTx03ZJHCK8GoUQ+D/y5RIVO0mXq
9Pl82/jwHyq4UHauNprMJEx46LESMRaCrdalSysCBrPyx0Gmhf4rMCUTAHfi8ND7uOTtw/Jb2id3
lbUExvZIH7M4SmfuOlFA4r34g1amJYM8gTsQ8g1K+icsKYmuDoKj08nKDH2EV8hpBMN2B4YfBEql
Z7Rwb7iRaYxrL5cEX9bhwEuDUTHA9pt+2470EuEZTFQai6DeYab7WmWF0vlZK5bvkhypddACWCEh
YyLYn9gjlUKumFoEjbYXZ4DFWCmmRjhTIXALxXaDeF2kfctQ9JhTnLpCYYEjAZQcsMIhYQHHrQp1
ydMVb6lUH7VI8hkBx/BxRTA5jpzdr6ibfFsvmdbOI7+UyY2RwJPrvowjejk+OE+U9jei30Q7Sj1n
DvGAv35MArO3jeArXrCHoJklrXI1IerDaO1rwLCnEDxpDwHcIbaHwsvXCXvx+Uh/APRUJlMw2beN
ot9Qmerd/cK1hpbJ8Pcodlgb5iT86RPP5zNS2jmWfNoPs5HbY+CuPEsB6wfA4b3mecZsWFikfgS9
6U8ypfriiGbyt+6X4f3O7Vo9cAUHKPPNa1V9QeXHsPPkufRn8r7RIZNwushs5P1sLhgbEP8bORlm
YwYXfJUPyp5PgF9VQEEogFA6VZ4NJnCGLHZ6jqQcHz/Qp60+PS8GBSm13mBoLtxkBUmxnIF1xs3r
WFvq1DgYxyYfEBEbq7CEVLHVm8D04T0VPpsiu9Vo+x8eZga0GApsQ/BM7TMzBjKAac12BFdjhDAf
Cn6QVy5T45c4wRLumLK5l33qdX/TT8NY0TE5lZ6dTh0CbgoJfKJ8m6Da+ZlBkgYzuycj8E9Y5M5N
Acro/VgNGV3HGeREJuGd51PQB8med+ZejlnlLXnkwgbgsabh4ww2kaZWF7Wcp03OrGWLZQALwxZF
I3l70TF5rZ88PB0hokvlKuz9/dXa0q+W6A35r+uD9J1RZl1sFyK2Ipi9APGRUM99yq8ZdcbwDAwg
XyZvNtam0zM7yXlmLc+piAdiz6TOcKk6p1skx4dzI/DrY1W3dMXW4LLixnoxPbN+Hdrim6b8JoL/
JE3mu7IXu0bMLlrtq7dXu19n4iHOF6VnQdv6izCCO6K7dMkraVdHTE2Oy4YBaB/yIge3ErnjsA+s
tdXDX2Ls3AQHrrQZLNwVWqraItThEHMRe78jm3a7SkvPt/jH69zZFZ/EtT+9ld/D2aB0aHROpz3M
yI8wZ2cUx3UL4rhbdAF7goe+BimgpS14LfO1cDAFwyHtdO5tRY3nXZH5DiTdgVx/k1n3VjoLHfie
cMEw3Aqwuw1OopMa8SgmrPTsS+p3s7oyn7BJKOO/ps1ej9aE0xsgUUYN9lsHjw5DGVCyXffXb5Up
DfgUVu8dr7neAGAE+YCRnxSUOkxGzcPhWh1tyQroh5rpGMFrnaEXlcH9A/aFWisua3hiLHGRre+R
9IquWsTeE0Njy/k4BeWlGsmxqTWXSIXFuFoisX5ovMsEGNuTTLzMZ623gvuL78pBQmCGESYF3COU
DaaBMQaOdJA0635d2evzJlrxwCSoFJkMbkNbEZGRkGJezccwAoFciDEmDwe8/PWZQoItx9ny+yad
fgC4r7jn/SarSF6PCb6FpbeE8exr5/S4TNXonL3Az+UEjTI42X2EwBMApJLl0F9ibl6RXyH2A6W5
ludHtkjLW3XAwlR/rKZTRJazQthVhANAe7/3UY90Qo2BnyYA4DK1EjBD8MPu7O0WcDd0rGnH1Frz
ZcdOURrNmUMOAXxyUNfv+Nt9bBx5rTuCvJouR4DiGFtU41cn6CKc3S6QeSDKua5NdpB73S0FpItp
kmPBFQ3vII5iS482UqKkPGfFeZz0U1uWSrKospduqK0CxruIhouZ76glrjvlprBbngyVz8i/rg1H
BTYWv6jLU/GyvOawHqjYbzJushmKIzgsirFXiY+xuCHQ21tS+/NrIUFsrYblZ0Kc+rxtEsdb+vO9
bL0gCVwUhG37letADvGD5ITohD6kA2MY1lcZIao7xYeVv7MEfcQfQNiuWr4u8Op9yryvrty4729N
tNTkoIzRNYiZe8EgLKl7gKgbqDzQywKRfTX+NxkkpP4RBUj2vgus+YPyWxga492Ru0QlFBs2SCJr
k18OPI5z3o/3v9TjzfZLTwZ9cH6AxcSJj6QXvBEekCAR8rC7VOumqKwSuSyFd3cKyTTgzOp+DEbm
lbqWmUcHKmn0Nc6dS4mRwgZK3JAGHpSSqB10/l/hWUjokhBKIBFBARJHhY6W+MmUbVsZ7p8Zz/mi
SeGQb7Zt46I8jFnnuvsUKJSxpfz+3mMo/8d/tBZD5EFpeB6MH38Xtz3DYboSOGR8XUJtK/h1sm3f
1QLKR2F59mg9n4Vj8rpFondK8YWkcbsqjQz+r9jolUnb0QDCnqWVPLE34Wv0e+jV7l7Uthiz87iP
hjjmQcwNs/byTvrcfXeXdIsQOmvpMPXAmixWdxQ5Fm1yzV0fsf9UCTcA82gc9lozXSNwv7FMuN2N
cfUGuOdeW2SFZyq44klGb7ooH4wImyjpIJej9c9GtTo9IQUTM8fuBO4ur+aD9obJrh+8nseWhDQQ
nd6pwiGDemR74YfD3RRdylCm6PxehrzYvr+lXAUtns8k4R92J/26unHTVXes4xUnjqWQtXhEzOsX
xKupeSbUYLl52Y2fscDbeAYL3MIDJqJYD742zoxrB2sjEK2MItgFpMUewz5EjAI9C48wMvvToGlH
RNYF7nYualeB2bg6yB9wY3oz7c1L1e8iEfpBjdAJx3ELJKpLvOwoNVEYUXwqPn0w6+FayyOelQ0T
mGPZp+8rERUoG1eMymmZxy/pj4EdV78g6ZUWsVA3VjFiRalOrStwzSZ4E5Ws2eW7G2wiN4OadaaL
jM2FG3uqLiEM5HoynPv8+K3uioqL8rM9yVL4R5aYy6vVDNZ9Ai6CRpLfdWW4GVuwYfK4eoWStcW2
JOoCRlhJ6i5itMYgt7Yfl+nOfG8tdKejtkU+8TbePR8M5UYP0iUnJ/7+ZvvLE7GhuErONXYVPGoB
UzHARe8Iro6y+KUUILtkjGD5fGdJyYso68UzZhqaf1akk2uKzK4XMAHVAiSxBGYOdEFMORGmcueH
itT2w3MWocIXjAlnLf++FtUJ0dx+CLG+0CQKH0FihRx6/zSWlnw1NcyKfLOmKdySZepmeoIvVFQR
xWixPkI/XFj+vyaoOCUbPsLM0Hf0HZ+iHsAXvvCyQOhfuwppdpesRbV8eAXeswt6pb76Ln/9rz9c
JM3XatOjtVUPvX46QwjuExXXGRaPUkbrv1U2ohS9ALfVloHs7AolRw3M2fTNngDZsFYTAfAwFDef
4KkuVAiQRMkPjxI5ZaKDMqr0mYXuaxGvq/bUxkUe9yV/3ADewpFbqsALL2Ifk+FZVWIZi/1UKQwF
bFkTtyqjt76ZqtMl6RLzG+Uxtzzk0qhgXuUVqw2Iug8p0pFMWraLU6TFSdZ92xx7picUQ9eJ1n89
TohrIh4XxEwUVYE+bgYQ1SBRKjOyh7675f+2LVo4rgwgIAhu1a8MKArE0GFiqhJqy97/eLk2AIjX
VDe/Fz/CynGZ+/ou7ediU7uhQ3RzEdHBkZsm/xfh85ZW4e2CnYQJV8G7wO92xk2Y0O+5pvb309Il
5hv4d7NIdEG1w18Y4odWnq6Gq6QohJp3ujzFcjSn8gPDNO4Rda5yIaDrE7lGOy/vffRXhDtWQeis
lPoFvTHCDgBZHryQoByyYgyO6vf71nfS6aNovxit2d836R6WYS8u6syOB1JH5UGv8AI3m1FOhoca
f3hjvQ/wzc24wuQgTgu3pH7LLPxQzysNsLqDAxZmHp4/zT5dur2OZbRjEsX63vtCjQvHxthuzBrB
5ylwueGR1CtwrD4MtXdTAGgfg0FR0Uy80VMHKn8EMkzJ+MnEz8e3bIrLcZswfGITzTL/L03qtUJl
66E2SlF1DlE9dcYhL1srmcEyrhwwMzWUyu1gg1E3U3NekeRTJR2nXibxYNPk/vPwI+2cejq7u5IQ
nEJI9yqyM+fPTm/9SM5FfoNpOvmEXem2GhL3mfjkDzjDyD2Ai0KeicI+blVDApTCnKnJMn/nX3xM
45lLrTdrrAmV/eYgstE1SDbdmJVtuxJ4OUzci5hJYgTjHCJ9EMi+kalLPztBLWFcX+WcObe2bHTI
ZQdpiz9WmHtfk446xT3pzk/QIiI6VuQ1bIuFHDNFuZsJrBp6Vb8W9bKfgepgGBVlcWptNx0wUKjY
4ktads/YFPmv8mFUI+4ELE7YCGG05HbuKF8lyfweIz8hTBf9RbGdyDRaa9byDTycrzuOpughnpS7
aoaecLXOJoww0xMFMtlpAep5yzvUxioFfAUI1sJwziE4KMFvGpI9nreMwFZDfHGM51hgZdsGF7St
bhioLZGdz+TP75qLvzO2XSAQuLEyN6Nw9i6EEf4OI3YzKwSpCNxpjcSxd12wdV56kdMKvSPaDsqc
XHe8aNeo7N1lv40WACTdp67IrIwmTNYfhxKsHkrMF26BOKu21KYjr1CTIunWw9+9SMttHSELC4xn
64OO31fXhyEsRbEReUGuw5rNGujytwliZUldOgMWVcoqu+kZhEPuV/wKjGbBXJwxEqjadwfHHv2G
Y7fti8xHAhYlHqq2OhgajPJNBWdLzSO2axOTWtEU9o+A20ejNav5RViFDZqx8UK9GflTLwd9Na3+
OLaZ0m58TemFuWmD5WiHTrPGzCe9kbUp9FmzutjeeBJ+7alSqbXCyaS8xrUSADyZUznRdhnmR7mZ
cbbUerFbSY7k8JDl6dQBcsbR4AoDOYTPxlBFvu9eBnEkUv/ItiyetTiWQ3WmtSeDz6W79Kl2siVe
+NE1R7IUkveXMQSQCnbqglV/7Uu1f69Uh47vEc2do2tjTlvYRFvdvODz9XrQ/RB6bxaxzvM9AduU
meV8tV4H2/6aCwiAlWGYKIs5/FIMnwWeHiJEUAOsW5+bPnknvdAWBjhrgZr6JmfW6wIrj+F/Gvlq
DBBP0B/J8T+BIvgCuqaFUbcwamlAfUfNyhNDbhytr2vSjpEHUQtf8RjEVXvErFubhXDAP47aRCGT
S460sh8SFcgwdb5rFiD0fZZTgV4uzcRvQ82A2vp0VPAAjNVmDvg/TkgQi2F2Hxa82wrTYCUCfoA2
ruyEZR/LdKROgQ0V1pYK1P4v2K54/D6ABEg0piTJuvD35So170Br0C4Z+xoaV/TsaV5CgkGFOoYB
y/eLwWdaGp/fuggBS3Kd//W2knTFGjq7t4OFwTtp08HXlKayPgeo+XRHIqghUyPoUckDRvy4mBtj
Rynr4JbFKeEQp2DU8YUixqI7g72EhU1u4ae9iqdW6hBx7f+nqBqtpo+JVxqoUCDRNlp1XvRxvwR7
m6PaKjFQKXY0TLGK4OOFiKem5qtHlVB3sbwR+Sh277KmYmGNyn8A+xOFc71apG4YNfyCAJNV088s
lXK0ZL75N8FV+SoMfmozRaSUrCQf0PNNa9ajAuI/3EH7acERlbyx7V7SesIco1rT3z5s9QhdqF5b
k7xhFAymzVGzeXB185q+5i1SJ6qCdcvb5GV6FjXsC/gwxzEGZedctVjWHPg/K9FX2CEZMajQ9+w/
wUUlA2jfAeFAdNEiH7/gnto0a75V25VdGp5FAPCsvJk+VQpWmTkiWX3JeFQaL4+gE7f2st0pa/g4
SGaf18NGyhnN9M9Zu8C5OyMuEv7lnQgo8DueOi7OvDQHHLYMdfa3Nz0ynKBr3ewMP7LUurLaJ7Rq
cFSvbofmPsiAkDgcfYTgK5Mfb3l5QeAfxNo80ZW6S2m9lGuGMVuuV6nHk31nDF28Ni69xCsPzpPz
YI62T+TvMUHO2qTZO26osGmBRl2QjSvTOLyYX30nDfvoAua7uc5SDFj3KTaXbTB6D4R6g1LbckmC
lX0h7wUS8pgeoJO8TYlBkjnIlND0+ncLdRb/CNzHTyMPzJHYbaYt+SDMoPgUiY8dsb+nIGujLPvw
GJoOUBtPrDz5XFnYRXAEt5+H3wnETSRIJ1a9hf4NTyFlLzAbvFdJyLl7ZfPDTZLFxYJabMpWpTsA
P7XC/KDioh+e5Xlu38hyjZak45+t7boLdnRUcfRYO831760BVIycGMgEtPotmFjYQ1ep8kLbhVjA
kJF5BRsJI6YjfPJ3mg+BigdEvYtdMSelpOF5YGiIeWN9H9Cwse7zA7iopFF+m1U9LXN20Px83Hbj
F0lT7N8y4IZEc1EmBn5zpwUGeXoS9Iyh8Y5mHg97RvB7VCwP2eqeC/tsTpVKF42AOAXCOZYElL+G
S5lxUMf12utPQoOgYvQVROnc8OB/KC8HnNcT7O48LNXEuEtnPSFMknqDJ47Psli+w+EIH11zNf3j
wn5Ds+TIC7rfkAT5amAZ1qlpS/FAQ6mAGdMDaTEjsnvC9jwUXyjPZGZ45fUKl9L13+d8FW0UrwUB
sLS58j5ow+qCly+XqhCndAcWYfAmh4JyvHkVZq18oZraziecz5TGiJnplyrdP+GISjKHBLAmYL+t
pBDhDDwvfgEaKMd34fKWRhZZ0oOm5S2zLbFkUNhn307aZ3UP9pN1ah2TzsA9Gjzp1XWO5hUxSn84
IRR2ft8CP2zQXF8SP9qrnH++xIqPUWMoXmLx+lGL8zPoPoxfo3OZOO5X7BxsAhQ7Klsj6lfwyg0z
WLHEpINnM/W+n2KjkAhqQUA644ew3hT01Vj75nXKIQZPCcT8CCdFE+/m41vN5Kp2KFQZlBRyKBOm
Dr2i4N8LYPpZmQWH/G9VSBCQDLB2fAFpaNz8I1ZnqmJyLnINM+VpYUUPvRpGUD27lAeoqqsF8xzw
a/13KC4Fa7vFBs4dB+QboEXL7DDVak/DPQPV28Y1dQRoUCxpy4TYqp0EFf7QQoM22/oU+wxhDZC5
23c9e9Cj0nttc8qfyurQDKyoZ5jlckDIJNknVRqvS8xBDRMRghjnYOkZtLGVls5yzvo7oPqXc6fZ
JByRheDggM+uaOUHVOcS1DsV6mxQ/2P9zjC2e4Wf4b2ha7/yP2XgJJO//0/THpvE7BYixz+50kLu
EjZWnCKxvqpTfu9v2YgkAOg0mAl6fszXMshbRn0HRAH8LVVOlFrNtJdQaV3bWV9rAJjYVVKvrHmO
48vXVXtrVvan85QBwfmeaK7ZzxX+/ovKw2IlxSBdCZROBs8ZubX3fK/9tbopbJ23mZbrBzBVssYB
s0z91RrR3jaPDW8LJzjFEQs5A2dOgB5k+8ahwqoM1O3Up6t9FjxHB8p+Q0OLXz1GUU06z1WCyMBe
RDEJ/M/YUklWtTv33bcp+VSoHzmIsP/9YwQdWvlsv+xZDUomJRkH6aCB1FDLIurfCSZWXQaJ0XnR
gUnAkiBFYtWeiUqRjotOHXEEva+FFk2u6A+DUmISvE83HWWGzBpu9Oris3aWG04KuB8WOFTIcSVE
TkZNPNMWLmgFGYoMNLedyTFsbC8wnO/DhZEkf102fFvmwDwAqQZwRA5YE+ARNvGXArlkWiwXShoZ
u9FrkcKRIBYgDub3l8m2qj1RHP7ih/kO+F9K18jREbEpGUMZRXXgWqoj0Wz18a0vX4Q3tqmJypkr
8VwLsaUEY/Q0j2dg0A7x2dyw329qihdTX8SjibzR5/AlcMWSBBfPYgs6Cf6QBydcTQ6NUrEm9x3G
CAGiGtpHILHxm9eFIl0hjN7bJGD+FyS8k782ow5pLRQGbEFKa7WtTy6aAX2rLNI4FWnGXyZ1FKka
T1sUujZbzTUhAbnspzWCK41k34pHVKM2FjCoL4xOetfEKKTwdeWTMZObeMv76m9skGXt25SbDO8A
dmpyQbjx0NVLDV1Xh4N25YLh4mPHyH7l9AcYw9kUsVWLsUCDOls9cfk74C78Ek/457t2/JGCplz+
F8qr2QONq0KP6H9FKf56vOWLMh/bEY4kE0oW4oWWDoIB0xtyIBefM4qsjPJ0F6bsy1ZBOporXwSI
GPV1Au6FAFkkNP5dqI3Pp11LveENNejiVIrefT/h+9QGTK4JF0e/acUM8BkMiD4ZtcSlU/8sktXE
Fi1SFNVTm0zCYWmNVz0hQSBJxnX00QuLSPfKFX2eSxKFt0bbImf5aNYWO8Fyb1JAvE/GE5QibRvB
CODZ6qir+74UFRj17dqCXMMWLCBJUf48LTKi1TBM0JSPqNcxikZh5TkM5f7eKqTYupNu+QzLQUij
8l+g/9O+hFBkU+jmDKjta5dqpgPLHW/5qAT3O6wOlDQpZ7F7+Mt8FrhfByWnf+5VOCC8sJqAOWLJ
+CehAFFYohxxt3620YSGTcciOpSx7Y4CrMPC9UF1bqDvA8qMVhG7B/kOVOla+6W94KAoUFIs9FG0
fSPwARNgnp4sEhMO0sw3kEJjUM9DKWeWCJ/Fgvr9H+SSwdFAqhhOqBWXT7YhWHlYcOOvB6Wbfywp
qZvKMyoSZdi4zNXsF6mjgyXrL0yVVJ0UkHYmL3BGhEe4ogVzUqRIQzZ6TMTBxGLnVDZDvoS5rA6P
lZWFJFJTzon1slJ/6drf3gGUFzbMngzhnmT0KHAlVoXPtkN1pcoS8LeH8ay/SsRVQojIUL6WVQ62
EjSCz69rsnJT+7kVgS+1Od4GuQEGQJ4WwctVmucGvX4ZJqdBRPEOmKRZUhzTwrhJnB4W0GABHv7Y
aZlh/YjdbOBqoWiGnlexSLWvLqNpyUDeDe7PrUv2VXTxyTBMONcak1cZRPnbpWoYm5CwCJdtbGt1
hzaMZl7OLAetcoDE11mCec/LO4lm6Ace8KFOH6BNNomRPa9ftdWgoDaRpzwfF2xY6hLaa8fVNmng
y2oYOmZyz+8kGqsJTsFSocV0V8/V3nqKN1iRDXWU/Gaec3oosYTdNt5ASTvOp76k+owzKg+f2QT0
WbORJHtn+92U6rL+Z1J05OYkZVdTFTv6ki3xzeJ/fgP0NQm+L82EtjrLGyXS+lyXa8MEb3eQnl1N
zbwa5H1u9+JSH9PtHMl7N45dbyYZrxUDrGMKFEwP/Lfj2zNoCbAiBDlQdfsC1CnSZFTOXhudpTfE
KIYaLiOTU0ja1YaMHx1Uy8WWZkYl+MCNnJBKocYD3tz9Kh+sCWNfWDnVea4SE74mE+NyerzXt0il
/PBHnEMnd3z2ar06g9WIzDjwGCMSzr9Y6ygiK0gKZq4z6izcgSATcPdgEWmEoIuVGD/Wn2j9SCTV
cFdwM9l53syO7PnwTlenD8tFU/tAkAdwW4j0qw19cH80h5N4/yABDnN4K51r1/AYrgNRguaJ9WNw
ezLiA7LINeNpEtI98C5+bdvvijIwuR3KVyX2kIAffMvvr/4bXDhyGlyqN98kcVTswhxtLMe9kEo1
p3vV9KipGORUWEm2tdivibIvx6+S9ehg4rUIaAEvNsQ6/q/UOTX7Ym657g+aULsN2JCGFEbsEf/+
DRC5bLvWLZQGTt9nlX/hjpmVkSxBHyD1KvdenrZPU5xpTW/ch4fEE/MUebRHr4PEQ5k23MuEKIaG
/8EFVstmHKrqo7arL0CeqlSKKeY8Mf6cVs1wO991CMTzwW3xClI3pQgM8+i5Bdla5LtKVg3hTwX1
cGcMFrnTzas1nmBi519XxoRJF4EuNVCIp8wekelOijhfqJRRIuzUu64CwDMoNU+ppjLdoNBNJC2Y
FGEYh08PsZ1iUU6CzYwqVYypCjBBRuud6IDPxLfLNh8XUTN+Gks4+b3TX5epIU03tljPh4K5SSK8
+w7K90oQC3dq3xGO6IKndyeBwS+iakn4C6Qj+T+ZIgVFa9Ur9Dc4tj7sw7jvONpCPS8mGV4R0C+I
nh1u9u/DDH9xxqHDRY8x8U22aCKSleBR88/8l0AFjpgNgNHbcfgeoUb6GjfE1aea2/1M9h5wQqjB
ZBCLDLXBcZQrQpPz8pk23ekwO/qNHPWu9Mfsj5oZSYK507dKOXqbsFWVHG7Xg0cG6eei1q5tzvP0
prSonimkBdl2WwQ/rQHblmEa1eW5Z36yZaPpwkGovvJrn393rdp3qCUrfjIeHwBTPgT4m36K/h2U
COYYrZHhgkpIoyVLgUL9//Pr0fG4NUA6d6/R2tyrSfLeoQgdfgTgu51Zt/VIdQa/FRkUVBknjlpo
se9JLDbeczKod9zxBvsvb4S5c3T6LekdRZK1i4VBqAORkgOdqsVAtyD5pBZ/Sx1fY8x8nJfjzDFV
9uwfA/J7i3ECU6LNqVTR9PxLBvRMiREVBgrki8kF/MQh5R1oeIJqdm7AaXTKDnp20P2knBXC6+4O
D1VMdmniGBUvnqC5eyspzEFlaE5LVyNwQQ2uypqSxdjgR1oJXzu9BQe4/b3BQqyEpRpeVvtNlTYZ
cSNxBJldbDKWD29ABn+/G4i9m6w30W1QvOLGmLapbdz3LN777GQazWIXvZfloMEjf3uZZm5Ybn15
OPBbTkF6BaL2DhVKKNVG8Flr1uWXbs2j12h8dFcUWjJTOHQeFyUQDrRgs1KDVs9OuBsTZUVzHWjI
pozL8cEqETGPfg+Ug5EORwyukXmXz0vtCplbgQtNx28gM4GsYGL9arRJDVB1KM0O4obZPnL86zfa
H6dVCHJNmkyLRSDBoXQfjFi86mbzlVbSfhZE5VMjXpWJl7QfcLAZMchJFdcTkw9tW1Xhbn/RpY0n
y8Oh1a8IqMnoIXddpEQ/BJSUOrRHPos7zcCeSD6ud1qgD5fB6fVZ8oxf9HLBJzex+mPdDXbwJ3AU
m9MGl4Us/inLHAVLF7LQr4QAAikcC7T1K7/j/tfFVc+aFviIZBFfMWCbrQAp+U9V5zGD+x9o5uhE
c4ukwrBhUR/2dPCdN5Vjo12vaWqHsFffP8wccK2ybJ5di61WLN/n4CXv/KpSDtBIM+PQYPw+2NE6
Ve1cXMkGkV6aXA0poZvnbg5fsOOvMXGt6l0Si3BhWD2YKo4O1sesQkxN3APjKFRx67OcyxwSYRXl
0+QMgOEnBLBnaG1RuuH5ENjmHI8uGOBhSJL7gq024MCRmQB9t9IUXBjs97glpTY35whwPwORfDw2
oT6XiP88SobZ89mkalETdVY1Ep8CmgrMsRmLbIlG8580DbsNmI7QOpRBPKXBtkDQvikqvYz564vd
M8o296KDLxDyt99PiTvefVRGjTcuadIcYeQpzVeEosX5c1z3AUXtv44gIsHy8C6K3oxz0ylf9r7V
aw/oki6eXT6QJewSW59vTrbP6a51XiDD5t0ENw7hnpA3biF4e0FUn2OXf/OuXdtwVzMlqtyimmYc
suNsfdz1T5pgbXvW/Zt8wgeLA8NiQTahGN9cLglIl7Zi8Vos/chQiFeIKfC7INuDGyTZL1Lzlp8J
P6Ducx/oyFTwRG1VN0jx8/ASioP/aVIylXk12etRopyJP9dEZOV3ybHKZvDVqiO+XCSWd+mN8N8M
y9zR8dWM9FaJqCPChablIaEGeUPz7ayqhW/PvEqRQSQB/V5akdYXXRlepMmtf48bzIfVg5wxARns
DfJlCIKkmEYFfCZp/Rrql/hDgIsa+OEt4mef0Wwl/ZijfWbM5p407qisEEFOyibeV0YVPNxAEP1M
FcMes0smd5nyyseYDLMZoUdPxtc4KmalGPJF+Eg3sKDXFotjCrIczxKSXTdOtPc7XRkJ7jA88au3
gkGw6yGhjiCpCqTJkVUKIh52HvsumUjo3OHD7Z92sIgD++i+xPsiXHUuFD2WPqSe4F55L8qIVgFZ
G17OqyZ45yBwf6AzhbokmiRkbQiRto64zMZExMrI4pNFHdnVeRRo1Q8v0PJnf8t3AWjPwgPbY2DC
SqA62Ktbmd44/y94cp6SYD90lw8Hfad9QatoCBJbWlaAgrmJropHVQHp0zUGcvRfO7LI2cqkPwfs
XhpeqZWPufN1RNWHSUVR0nOCFEk1uqm0W7cPYPLssYTf4XfGEMmYA92WKgfgjX+20sLpFllN0msd
idgrmqSEEq8pxQ52soIGw/VPRJYivt/emsxb2q3dDN5YqTIJYna+3BhJKHwICoeSfqpDwaKzmGBS
f/0UQwDBB/muFDSJs66Tr/tkhTbP8BerV7PAG17formLSu/t43pYsIbIbfyL9WEvrzaQrYo2c3C1
vY5O4GWsM+Bl975HN68Mw+AAmmbNq67iLm9jR++inZncruFuYrCkICEEodMfW4DigTLmdh+/9fOD
fSCPs6HvrbybZwXpZGt81F+Rul16u6N2h5MUy1nhHXvqF1DoTNtB6vT0O521OUd+LjmD4ozoY3Yf
dEvb6e5pJWnlDVjQv6PCj0WSqDYjKSo2rWsfoaHp1OMudp+/gPd2TNjHHDjPP0lGBlhXhoe+urIZ
hi74eYiO040USSakpGO+i5ZNCgMvKDXPC3eEXKZkJMYMVunJtV8ad9BHPo81a0qVUVnmccCD6EaK
xgUPH2l14NLefAFmY1zAwiGF595+YPw+VaPjIciYfEZvCsl5+aUUJmCwVpeXMjfcrzJ5DETFKo6/
AFrt6yzQqFCc/WFUOqPMYDVXlyl/lV0mKDp7B/CXg+4ExrQ4ndOGWNlMGZiQbc9LIpQW8cewwzhA
upXWX1kJCfsvsQpg9/0x/W2rJYpV47QA0Kj5IzD2FGkO1VG0wrMn5MiHQCvmdR9EZkPUqX4LEhrF
VdXi77LeYSqpYOeBXrrDwvtDso8AHctGN2kySVBRISnAugLOtHMYzfE8oSt8jKbkWci1GGjFfWhK
Nj87ovmNjcj3avToCf0zC60SKnvYGRqJMPurXOhJ2UfcuC/30lHKB8VBdblbQZ1nSerVQhhkoHpO
Iv1GB8VVYAsYRofc7YcbCorceQfjHDcdiRwFQSMNxQBQBYvYRXjqyO8D4AyU8zSciSN5rElnzxzb
5jTVVOKrs1pKquGeeUWt8AoMwSSki+ohlpbrFSVsoDsQQ9vm5jkByPnSUMLhBNwjh+r0J97R6GyW
XASHWYe+B//T4eFaA1+1L5qVtJck9O1qdxBcI9k/P1bfroOektVUAi4HljSUA5DB705qt+kpSOyr
NH0boOlBetNTc8PZWKlT6DlHcAO+Z1CKPJBzmsUtkOJ03/euNXv/RqGXSWMoVWuPvQ+ZPpw+uFgW
6nT624TILCcwqaJvm7Bj+s04bj0mqaUsNefYPo4ynEDkJS1SI1C4xMv3W/VW6kJQXG5TOdK3GZxs
xAI5A//HADlECmHn6AOD9QlTITX/pyVmK+/hW071C3JJnF9NsW5reqr33UfvAGR67ZrN9rAHzZbm
fYcnSWv/acO6cIypSRpm1ib2v1G7uB6nroWUDtboAGS/sewCu/z2ci3g49JpdfXQuPvdbB8kl19e
1PwGhO83M1/K+/IMgrbw0wD0NOCQe+PJExXHNAymrwzH0juhMjCirMbZByBkWVmGV5z6MspQ26/Q
JGwzhnI1rgWvoMyGbud6JAfn1SCAFWP3s2NBaONfZ9EbZ5CvHJsXqDdaXZVfSXqAB4jXfcfUyvGo
SyJlyf22gwfqqB/XUrHk5ZgDn/qUkokOVy/miuK0fsGGJXSDrxzRAMkFA5PaAC4xR3RcLQcRqyc2
cOhJSto7tRSw5JTIsWD/IOP78dzyY8LNm6WhjKQqo3RJhh47zfLWCcPQBjcEjI3JGPaPfrvRnakQ
cm5gNX6sfsZAGB/pkuIJ0XsabHKIwS+oGgfUCsrKQZktgz2VqnevGdYgt5huzWgViXtxASVhkPvv
PlUJyZeQf8TwCXfPpeNXkZB3IXuyEGItA7d7DsJgpcS6hFhk6Vn/NKgrWlqRgegz3lRN8sEKYwrI
XmBIFNrriuhVbUVCl31GaBjAaMPbibfn7kOmTp3WlEPDROR9/BnnXaVC5+d5UbqcL+FIPo/pffb6
bV2SBWGsN1bxc2fJUIg3cbP31OqErb+99nOJtuCosa6cT9tLlSD1CKDqFjLr0LhsURjmWqhHLkEY
K4koz8ImVV6rOCRL9wrkSlhALZ4WjhbZ1Jo2Ar8EKTnp7K9Rt4XfSwIwP88JmFVN3ZNnXt+NjODd
eM/Hcqimc0CwCZlp6MYDzyU6xV2Fgv2McsMbaAUjg81vYHc2KV5gbsHVXt1EgPad7dUU75l8ax6o
VzcLzYBVJlXZ06t0nut4CVypE63gSxKtGnrr0KApTZQqgSy883TK5F+o/O4QTC2+NPKLuD/+9CmQ
80ZCLwEZLTN57ErsR0wYDY/fGP7WlQ157v1q4TNn+WnRI652/TW/6JrvtnFvUybUuyaULPdK5Ey8
Xj2TjWpYnsTI1KT3tQTptKOexuKKPgBD7exc6h2Io4q8cC2jz/Lgk77Id0ion6d4ahtbAWRAYXFU
ZOKX9xY4BCjc19L8QZo4zcX+q4hhI4DjJ/WGPIwQKsmjlHqTH5aFZWmNB5jy3o+kVJirYYnhvYo6
6DcwJzt6YoJlB490ihHXDN9VYRI7e7fhtEvNepaRuHiqmwRN4rOjWBzsu45ikyzyxpYvWyQdpkU4
ZtE8GdGFEaZQZysfxv0iHwE7F+YCWOeFyxF6H4EdI9izfKQc1ft9oaUm6j9Vyk6gqW61ZfYBLqTr
9UqcafdpcblisyWCQTNgGFgj4HkGZGp5CD5hih9Jl3imLsTkvOXQq16oXB9a4SKfkEB6l107H1KK
4Gv76odTAphW7k7U93R0eA01uPpCb1yrYRCknQhOnTDhNC3OHwLfuMwhpMw2w7puZo559EMqBAU6
+hBZsMK8npkTmRXYw98Lz7Y9/3AVa+pvjMH6u4zlSG+1hqfWEFbnrni7OIvQ+vRe+RJ9Glh4Eojn
qaYpEr1s9KphYYZaigTBBcykYwvG5AxmLbHFnuwPfqglaKi76jD3kO0jhrDCCC3/bR8Sqm7nUkTw
Q+jKjvAetcJV0H9s5cMnI1iP5LP+hOOk8X+KVtArklW+GiUdSMuCOX8JqDE2LcOIijh4zID3zDjz
K6EyYg1km5qqquDzOJ/GO8R2tLI2CCYb3NALXRzBgCKEqMOHuDxhVjLUco/b+97wJf4GDTQw/v0G
ZpLVaslCXAlWyf2EvKMwdV6bzg8aG7g+ECOLHQLlByEdr0kTjma2vazUU75bkUwW+ar5I3defHMf
WUkR89vVuEha5whdjtVcC6TCHs9Gi/F8fbS4Is3slASVrdkoGnhVpe766Utt9Nl9M664cYSHW5Il
7u7XHFYqjjQ/QWY4BcAyOXAz4bEl4Et3HDOMI+0uBsXtRpnW9GKhDA0l8gX3WDhWsSPF5fJySyDy
qoNHKG+9Jy+hR/epoBxcAq1+I3dMTzZh2koX3p4mC44W9xWvXW1e2vFas+JNDi3Ivy6FROHWFDEP
N0OobKIdgoTisy0zh8fAhzNSxgpb2Qz2ZEh4aEY4Y3xaA12ftR9RTbroRYhbV/6MpGAkFX/Va5WQ
hHDIzOM1w51O2NjnkXlB1/FBHaSwRzpH4kaWu7GntrAMOYgAbRgWGqQ433xZZMcVekAv16QClNcR
dnVsfpGKHZ+nGI8+57o9tDVdZM0BIPFUbiLfZ6056nZ1MSG14WNw24Z9do9zkB33OwFK+/hWg4zN
N7uFBeiPwFsfnEvEWPm8K88knYOaZHR0KPzVIeWTP8DQOoNvFAFst+L8nnzNkHI+jNe06ewrd8/4
/rS+LZSdOPM4ZOOpKtCPzER+Gjpu/B3giToXO7mL8qD4+0LvNs46UHHU0cm7xv69co6x+tU3f2Ox
wXEnsbEQ6GIsbltgK/9/7JHXy1+y7URVOs23z8ogrRI7kje0o2Xps0epMxgjCb9ShVe3noemFM+a
EH1XSxRdl6RDp3llz2o0/XjZGGJkooIjcrNBXaEwN3FuTgdO8tzzbN8PNRcT+Y7nZWrEEOnF4gUD
ABHc+DS7hTf0wtHOfVGfQ/wyvv6+W6oANAMZh+JgKcqoQgKinY4XJxpFIm9rSmVaTdoLoXBumrVS
hkhD3Zinyu+VI6DLBmHlYms36zvGBus3eBZm6HtAcuXYpZFbEljK79YsmT1wyAhdTCL4VWc/5Ico
1vesccu+qWqgDhrTpqwiuMGtaheMlFWO4kcwEZYo8WNIEIrniGDdZG2FCJ/Oa3vIydWqbsHnWdrB
ntn3TJwnChEjoxuhnFOxPxH3wUxKQshPHv2X6FauN9fQCVNcwNIXhULo8d4rEwvfGeiaxz2P6peg
4Csk9Ncq/3JrgDI9b92yLuKkR6xZsykGkIrVURMQReyAZdko6ikycrGzHtEOarbmfcuLKCsKLCdo
PKS4mrTxZgQpUasEXbgXKDdGcImBTOw47O/DH4+tQ0faUDa6s92KZwNtYyXjftRoks73JNzPYsvs
+BNE+XWluHz0cHtpfJSTXJV2Qm47CVAbSzbF6fj5TioyBzM5VWMmXtoRvOGqmXoxYH9L7hjHLA6q
hMA3yWcsQ+8le51rIVF0X9r97s+U3P0RZk7+yLobwEAl+29ZgSrSYvaGaOWyKE2U+gdLquETYmmh
nw7xFb9BDr9HN6ZwdHO8bBpkQlh7TrzsQa9zpZs/hQWnZRg8E6dwp/FmP2AE/EbWERs8NglpVh/Z
blIpI5SeADp9F3G83vEkHp7K24svqdmnSD90eMiG2TcgeHhiuYgCD+r7sCayKSrDsgEM4hiJMibp
m1pNnRtze4MyA5E+vq39z0EhpGv7tYMYCgOxOFkKjrc0gzqCfLgWOUZ/gR1ZXO9GIB2z6YK5WKBE
RXqM8mPdLVGlhxRiDFFW9sEt2WWCaC7omxeK/OZdfLkZi3IXlRGH3+8Cdu7dmEr0xRVppBF8RSgU
7gYuWA5J13eYSNWK6QeHMttDu5jIVhfjBdtqUEwhCBl1qKeBo9etybBVu9bowCBSmbcxFIxzYsFl
nlLMIl9goYuQKhwPaeL8Pwn8YrqtwESgF5vZleMq73Z/WTcBTQlIV1R80SMejYfSSiYh6BGvEFul
ZxHOvg5A0s+Rzc8lIwF37zdpYl5NxzhW5Rq3qH1zs/uxfIvN7u50tEuFyWtK8BWUdqf80/X9BFqP
OgaFSNY9GHTMEkuvxRpp63CVo1GUHfmIQVDJgzGtugJoh43uYelG7bRhF3dhWH9bpFlzU4BCfZt5
/2L2+vLIWr8U9xK1u+bOkgeIzpZ8YVQGJhaTcFjQydvsdh1mN5biscmA/S0Ik2wssPmFRqx/fdVM
ss0d9rZUmDjT03Jtelcx85ioBqpomlWVwvhC/ajwLWDpg538ct2K3HTw91SFtoLJ7mQZZvq1TaHc
sgomZX6lGUZt1FJyt1XkhTleDfd31Y8AA2zuMiMm85KHWAxF2QksXiw0jsL119+UkOX11W86zYqg
tG7ESEMKw7tanM3pXEy0KFlMb3KRzgvBXAKaVw+qjO55we81tDXWUIpRtNDUSXwDtzICjBeK/g8H
+qaNQuZKDgMG51GuC53cHbyX8jkGmzruuiC6GpgrH5EyHuYYq0PipkB/aFUSUHHzWjwaXnzkf3oD
ZuLXpmZepYz8YT4yq1SoV8rgrWRWw243Z9+LpwflTp1I4HC5vf8RFeZlqyT2tvdNjqNZ7plNO5pB
ZGoMNa66EH4JiS47MRnNV+60MAIqcT1fcIQADtAVTd9QiqUDS1vLayUQgC2htuPXAudF0zbdhU25
zCqt69UhinHpV0h0DTK4QBim8nmFXZbFxBcnZf8VvLu+9OGVaeudt8Of0GF4uOeavwpsrXE5uFZ8
om1tuilmAYHSTwKTJLUZ1ZYUOoi8JbWfNVFZzKu9RGNx3w6ZBqPtXr0JkwYo/5UMmz9k3+LHu6Qv
FgbhOYHM+tJD77M69/BALtMvyvFzlxVFVXXete+sDpkPoAnZypXd41K/rP2znT7kRIbV5Zu6KuvZ
WchejjrnI8FpGCBEELVHtX9/1eyexFwlAPTgx/eW7kWfyWx20ErHfXZt63vmbRjFkslXFV/HGnf4
byz1baPNmLcsHX24IlUv/K5RI1C2AkIOqvX6R6i9MLVKsP7zItmlhw1CDciEuX9EtaNcjUW5R1Av
NJYyWO+gVBG+BKyDN4vYUDp7uhL2jpR3rWGqekngJ5Zykxg8lNenwUuQaJjytNPzJW7Gst9lkmkC
kFrU0OQLS2tXJzsXtwVOD/vJBww9pFlhHc6OvQTEgCvbchDVy6Zq15yU+V/6Ewo4/LyO6DkLbqie
I6gYh9gT7DsYn3AEjTHQAacMqHutZphh1VyBf55QN8cNGgfecWaeRfxgR3iUSiyTfvB2RPQL+D+8
zVNHcWnYBtyR82t/oN51kRnz3McjToQUsw+NqAkD2SlD/l+w8uk/5Bm9ZBYCNlVW4WyND8nAsnFZ
MkjB5+QMQ4iJMTr+Uwtc8GU+TfhnHocqYbB4fMUFngNYq8qQizK5Td5/HcPakG6nGyT9DIGImVb4
itKa+PBHTcUzaehKvju0PtiNJvSlbjXA86ifTPJ7yXxS2OTVyToMb6foBguB0qh+Rbi6jowA4F0v
L3Yj9sA2TKJE45zFJsseduWiTYsDc4AKt3Ig7x8X9Bm6zKuaT1cmOUTrk1zviYGUX90JwZeD/0pu
M6tASWoLTQRW2V1oNhfeUsGJIuAIUnLbWTLoBZns6cK8FHO0Rw5J/7rFf1hh7+C8RFFlrPMOU/MT
2kyJLZkM6/pHdlv+BUhnw9UiL4L+4O6zLd05zzVfPpd4ZJa6lWTmHNnF9W8snzMlWMGdwmLQosaF
0xB5LumT+u8I5BvMz4naqZ+u6ojxeGKITdB79DJh9v5zMkygIzFFJg/WWMsKYrPL3YJ1ErZmKNGJ
bsYj81ieO5xKkd5ym2vCNxDFphE7qudZp1gZMkBZUDmnZ6D9vtQMWMYg+9CYDLVIKLct+N9vIS5z
2ITO9n0Z+wVDNIKPcVezI4vSsqbloF/ViFXVwVEjq9XZijCjZKngB00GXBfSoeiR4CxRUA3ikO5/
gCIp/XX18W9g/Wy+NDk/SBejV08lG0jJLVS6WG/DHvFR28wz4gU+kY5PXxjdWhRFbdZi+3J5pMjs
iIBtmc0GHmaQQ5/ZRuHC0NKchcrrEBTQ5Qi8Ir7//QGptW8oUcdfHE/4ZW6W6elSf2HTMmWO5r/f
8ScloTCUYluR4ZAN5tdKni6KZI574uXokxgCm20OQBiht1I9L9Oa5bZloZTEsQBHTnVLKtZZoWL2
t7JxdTc6BSpGeorKecQb4a39yQb0hLauAtTvXUtxumrjWvNl2kq0usbUoWfTlZv4j1XO1ilNN8cS
/9tbfKsdopAnwFTy/EMVMrNGW4a19SW/7UjR6mH6xQSE24pk/BSU8g0NFb8IZJWEcorKYEutDJ3b
/10u6ePW0UgvUasZN86qJFuTiF2YcElq8IkbGAfKhauNNhoFPJBmJbHIVEy/31ZoW+5HurU+HYAH
U5Tn0IoYp1yuK3O+LwwQDgeumI/6yWFsjePNvt9ZL6WhEPPBAKQ/VdO0L1SX817m+waI/YhrQn0t
v+H0CI4Sgx70DHriT21hnsmb8ZV0jzuAZYnyd0aTJwfAR84IbXKsAd0HIV8Gc2lfuENxhcb/RhuB
9Pn6pJhY0Pb+Dw5DZ6hI4rjdqHPLPCkNc34a7bHAuZ/dySb1dpWO7fckQ6hkIOaCvw89PQzeMPic
pUUf97SV3q/qEGIhYGoqXeQ0idDruGdLtHvYQjj3Dour5F6oZD4N5JzUC+B061yZQopeyhvejNx0
yf0FSOyO3o8TtiVn48s4i7NQ2QWLNAcwCUI1SBXjZX401k7rtu8bH8rTXaoZOylonDdO0h3hCL58
/IzVRi6QoYO6nfxsSEQK8Qt9V9xhlHeZXmAcFxOXoXghp10h1GjkuNG/d/3TgdOQ1dT6bfmS+QNs
FE2SOw2o8A0SzIkcsBS/VK2ccsPqoLv/SWzeIRGaj+Gh29UlvwXqvrYsGxXnfPIIfeCPvZlUsE0Q
5Z6MSnTzKtsBSJkuiyrvXj0FGBq8I/qRJJh/eMrpsWErMtwDdDfgbSTD/9/R4Z/wDybfhFQmqiFI
TGq5iqDn9A9bkw1dkfLOTf41iNzXOnle4xxyjYEYyjTGjFJ3jsmZuNgwt33K+g5Rq+lksIUL7gI8
LX9+vKgx+UBOHEqF9Qo118WzhadRzrIR/tZzwjdFL7swaPgKR86Glcri05BlR0OCqxapvhY61OfL
8+EXvBqsM7ZinJ+4IM4EMHHVAtHyVPkg4Mb7VvFoc8x7vCUQXhkVx0JCMcIUu+DkvIfrrnfdnDvY
yvqZ1cPh+dHVFUK31cJi8npryzMOmVWSuCbp34Gr0IjlbsQk1PcYfdNcIdHx4obz4CVTbTYCnO5S
LEYmnBKu77gNJ5QDMUNgoVA9t0+WG1t2ERa0ZYUdlql9vTqB7ZiLylIfo4GcH6dSTjDmtXgm94h8
SurE+YZ6i2Ew/ldlsFnf0wNilv7FBDQNxBk4PqtwRBaRGU3Ra5Wxq/oLobmyij5GPANsleTpdAHF
4WX9twYvUac3mCKPfWuRbgTXO+Lyt3EO2Oiof6IQ8icvMjMG6FVwf0djL8occpuEo7d4H0doUVP3
cIEANxPv5b/lIm8CUCi9UHa2wYkAnmlEJU+RQ1cJ3VUaxXj7Oc6RDNnxgzXThCAhzu7fWJizrzNJ
2DP0zTC8uoF/BuOcFk20Dy0HU1TR6o7Rl0J5OrzikSRAEDntsG1uv12pXU17G8SppzuTfv6rz+/L
osc//69xDtxNgKzR6KoiINlSVtpuACWMqKspIDwunIGqaWbzsU1PkFnz/0zz1B5I9SCNXaj/qFQo
I0yp3twEglicr1Ta6Ipdf73QTJOOWSs3+l+UzqH39OkwXfh4V3ZLQ6j6ie4e3WVsaxLS2SUjE8gF
PLGIQcuS1AS87jg2ZSvTecMSZAaDDY2h/GelkpDMQf/UNp5XHGVvy4Um710eeHIfF0J2Qp/ejT5q
biVdNx68b8l8w5qtG3Pcxhx3zCyvo7WiXGoYN2Ugm+IFbSmLxFKD6CWAVqjTkLRr2hGUWMA3em12
i3GgrbQDVindvqekVudgwij8LMQLZvBbIn/wnM/w+9PuBjA9yaaXoHMGgEfvh9zL7HP/PZwHAz2W
SN4+pVZhmJy6HcsJiNMYSx9P1evCWxLWXimD4AZb4HnlHlZEbFKFVOV/XyuxejOPvL/qaCl4BQTD
n6XUtJ9Q/tE6RS95hV4f9ga4Z4GexnODNGMQtSPjIVuZZqHc74+oXUV4QrNlnTg/uEwHIXRNW0yt
0LafEDKFJLr0e0+sd1RGfF75pvqSRsQf0FNkEMj2Hlc+m4RblO2IVomnxEOoIp/9XkENPYDrdHf0
FAXQ35Dbl9Xghk1djgTfHYs2Bs/v4M7hH2FPQrt6uauJ3eYjZJpf0LmCuouEpaHgJ14pnJMiXIR9
7pDX9fEHo0M38Lkq1CUaMy0bzlkpy1aoeTlmJL4TongtDEkE7MUiEX8o/g/DeXZVXxAIS1JEruBW
zlIWmcsy05kUhSKT986j9Sy7PSKqojmZKPMRLODzlHdO2Rck4c1Fhd5iDHunerYEzOfdqMaAz9nC
ctcFB8YNICp9M7f/xggT/hjZjgf69ooBotYRsDMkY3HwP5EOCQRD9ns8W7mDGqbW2a1LQuAhnRue
qqS7uJBkcX+ho3utHixTlmVIbnnpKv1klJrKPFXwfiN5NIAXgGwbYX6i5gNKY+/RQFWI7P3v9x4I
b1FDB3elfpNUdAZrHRTjImhYUCqxXGMW90k7mjeThVQ9u3E9XEKqBQb4THdq0B4T8IVIbR8XgJzd
POkTCBHwfZKr8uTvxahyGhz/dvRIC1+gu4fLe5KHYQSzsU+SpSWUULCIEF72HZetnSXBt1V1Oqj1
MIRgVh5WtXXFOXXyPjT4e94V8EuJkIce2dfEKHXb5085k1V2WERlrbhDXE6ljUUfL5I+5KMNcy6v
aISM0vrfnt6qqcsXm7JoDzpeCUOe1unZh1+lP+qPutbAhQ9XpYxIC0Tuh02NWK0uTZOG/Vmk38Ti
sqp5wyq6Hjd/6upsqS1C7HI0nOSO6Ai0xTf4F5SHQpdnlRp8ooLFp2Fn0PL86jDKagAmKXfMNIqo
i+muFPsDv4vtaR8FEJf2SgAH1vMJYz6LH85dcubMMktYOvxWL8k2HDaVfk32E0RedHDUkj93llue
o53mFifMlC5hljZ91OIwt6G5IjB25eFEgmYUm7EpzKoF84kIOlF9xQQhXiDtUzhXbVJj9uc5LTfd
QOwgQbA1oZDhmmlfguiEhY9ctunE4VZI1AGcWxr78wlJKq8KaHeFXOfVzhavTIfJ3unFCIAOeTW8
VE8IBUksMHqTI8M2fN1xIOmR7SMpQtSUWH88wIZl6n8tNf0fTJCDa2DPimHcWcYLPcrt1Q0zJz7V
7dJuHhCePqb4j0UGUjTtmy53Y04HV8z7m9scPNkhg+S7p1TqhQKzilhJUd0piFFwsON+vByVVAZP
3gk95RtT09NQyIOwNwzHnTcpapU5u9FE3+wxmJf3SOacCLjfr6Nbh1rXye4QrlDaZIfYKUVSN42f
EPOQRn42LH2xd/p/LnkWgd6Hcvp6jBAfgouN81okMdmzXqIq3dxvYiVbnukO/3ZtjdstoMx3on1I
ROqfAJEnRQYXATlg5fTQQN1vQEnIy1hwHzL8JNjYeNHhRKrGLvrMsIdoNX/FHidF7UyF/V/P0kbe
rwspDPQXDHFLZ9Ft8f7ORGjQJIv1YmNcJDzHH0SOvtK5U4cXjRqfG2wETWpxsoIEbUKVcyeT+6u5
enM5bOlym17nZ7PhdYLsnNvj3Hcwfu/j7EQfXux9MM3lhX9cTwRQPLe6fsmWodBIAsLQ/qj+i2x2
ajFcMStkD3pEkftilpYL1n+z3uu9nH0sCMT4LcWG0xaF/18DCE/xOqIio9bIEUqJR9d3GJzQKeum
HbAHRu7aZ2DyAf4glrfD7J8QP9xLqlZR5ePPv6hu/ej1ShavRTo+aj0XMcgHSQpOF1+7kEVR8Cuq
+3BIlLAs191K7wpJZPs4DerZpFJflKEABbDweH+wKFAdx3WEhj4itQ+Lge6JCRt+vGiaZK5RZ4Sa
/XiSB9AKxOVOQ52Yke4wLtXdCjJO+kGshwN4ornSsdq26YPe1o7fipS9Dpbgud+Mds2DG5Zc69jZ
zaKxOORakrsdGiTlG7lYNEJnHcd4JBf3L7YzDRaA+TyTcnWpMiVs0k1nxcA1gs1a/QGhgPA4n2iZ
CSogiT8NFzM3gb8WQqlGeYu1/O3qR+udEF51lHI1XIf4H6CB0Tj1OYZEqAK78zmZXba8R/Mb5xZH
GVUVj2ygbik+m9bQ3jiaeYp1VPgvDCaQPj23WcyWSrMZFQRtERsl4rpwBjyXfmo9DRvVBCLNtP77
avIpdmzEAaNQ6rBnfadqCh7VvHoZ/83RCYwF8qHBy2wzarOBMtkVRxn0AIgpfVx76fByUUkU7eQ0
Q/hsMGbnmrWbmwyNZTvsC3fULKF0rTLmDvXWKYYMNrYN3eVz1QioAYsF9TMwyu3On0dK3KhdHrbi
jvLh7NQtmJ9DN3EDqniAMaPiqC6quf1Y3nM3YbKWI+BjuGnBg1d3NB3DFLSQDdBMjKPs4bWbjkGq
RwZlzCAFluQ76qNUi1yI47Edzrir5mbA1GGenduPvwg9+f7w4j2mfMdzQmx3htj0e36YlB2ogTVm
JSOCL82VYb3r3IzeI4uQQL2mvnbq75DOAGMP0zVnZWoXWmPbjlwRewyZ62mWMxpwyCQItbHHWIMo
f3cJ1t6zCbfAnPSnJSi+FaM/KUceyTKE3cSnp/idr4SvDjQpKX44OvYht6/Q3NSqfp/GCdzDm0p7
jAPEx4eafP4URFBY61GxfJ6S90fC67OqQOZ91IzbwCom/zEUEK8tktlhmzFt99aLCm7lPkGFD04G
GDlZK7/zNbwhNZ5izC5hlpnPqVPskZD4JhAjASXF80/EYJRqYKYhneGsIe1zaVk56NPRfPVcnnm6
AIRTPOY9exA5g9dF/gqdzx1oav/A44TfqR5PYFK5PdbI6bCdVq+qYepT8oDUic98xYB9tGkApc/2
5PA6Ru78CGj1FH1uGgJdcIJBoVz+GlK7E0BMFXGM8xK8iy2i41kXV1ZmvKyejAuhfI0teyJXo+s8
KZPmuqvDFiwGsTywViYSO+v9/Ep6Ftekg8SLm2+/rLP5RV0blmAlqspJKdpnv5bjCOseHq4bNqcq
k4RZWygUJ5kecngvYazUVZs4NN/QNElhHq9m9JubohmdDWYprD4K12OEkHlmEQly0kSeZSyPzZ8i
x6BAc9VWQoopMLcF/ZSE4nxgHPIP6wMYFC2s0lqtHTtpOYv09RUk015LgL47hW+HgZXdASPvgHV5
SGSr2IECS/5hvqpqhdHwpushjoBVtvkoz/0/t4n9ykqrM6Ksj4zxqtbEh4OByiK0+q4QRijVx28p
BMobTwdwZshycDXLgfQcZuflQW6FNG9t7VsbnQ7AHj0Z4NHN/bKDi0KPuSNbgEDjJIzBwNvZavdL
O5wR8XFgfSToqpnVB0QLZHNgmRZMYzTuneaGi86hQbPdzKk5Zo+xXH3xLKhTqTU6NDdCLo6hDxgq
IozDPpNfzP/dJu3Q/9zakmBDdzEKtEwVAQtrcptkzsewTR6b1xaPpx9IDMRGkoGpzlX6F1sPI6TE
k2LGv6bzNdjPGr8XrrVjcCNenpWdZw1BmQIaN4fLIWU3kheXiXWHgGMfI/iNOa4K8sxfpNB9lAUv
Z/8eDYlkYaOCU56NdB5MrbIFAcS8oC95JVtEGSZ+oNZ5xVDZxbTpIv+8/9phIEW6LGD8UmJWerpe
kWS2Lrzrrvt38ca1jrpc4gjRB7nV3meP6FlybTetdwO5cOcRUOUux+xCWaVgUclePu0Tfk9x7R8O
Ob8Jq+x2CLGatXynNB//dTeDW4wYeQj1NA8mGWLFeDSv/nJOlz7vdFVrwgSs9E9lN5bDf8xioAix
ZgW+bQeqvbysmKoAVx8zbFI/KKEMxxa4YpIkPx25rZCQtpEcE7/eSePIdpcESJ68JZh/g6HIqA2T
IjhXHURhWckFR3CsFXVyLStel5z9jb81NiNqF4Vqsvn/96vgeCNZysfEvdGrmqHD3EU5dA4CZiIh
E7mst3D/4utgd6hZH6iJjWuV+S2WUYO8LUY1umlrW9rQmSdb+WxOuyVxySdRLjLJR/4GqSJn21Yq
EzPL/w7LPx4IdWearKJIINpyuDEcOnfBHSe1Nf2D3VctLiO3kue3FEwNu/9qKEtR6LKUEz4bt8en
TXHue0+yhXSaycoabLgIzB8GzKp5nLTQruueav1I7c6XcTUV+VAEitBavtXuZjVSKy2ugbulQo+f
oaeNuPrxZTe2tcsieR71N5xrF83hZwjryFutCU61XiMF9kU2WKQF4sqam3292nJksUXwHvtwmuwd
Igb3xLY8kK9PqkfaSzcOlzNdCvC2miQu5XtIa7mNkkQTjqU8FvbI9TJAJrkLTA4glcTZdzt3gC/D
00DKfPFuKU7lEBe/a6MbYuMulYeaxd6utWGST3h3dDBAQH6b4qoXfOo4GEBd09UjyTDDtV6v1AGd
vC1b76TUvoISs/PJUonobeb2XEnifMfl5czvV4KzS1GlD3+rkbkcni5y8U4v/JZG/aHZ83h6fZ4l
ZhSJVt7ePHohV1O/JQadGScSxL2axBEh0qS80G70fiA3+jz/4Rd5Dl96MgL5KwTg0tYIval4c9Cx
J7BOAFXx11LaWDROaMa2w18bVPJa3rZzpAWI3Gk4aLVuWV67X4JebR0tQrMRQVTcmTRy4D0Uny+I
r9zx4QOAkDlfVtJtNbSvvzQZZ+lWAqjxSzZ6Z3+ZuC5/IBGQcpUfKJpAeZICOIjfQTXlVTL5HNtz
ZRfBv9l+atGArKabffcDD9S/J5g24uBDMzyeh//dMdO/OULQfBOIMyQqq2k3zQKbpEhrpx6nRBUY
czP2IxkjYYdBSMjqmS3YIDuHduNt7Bdjt3Xc/KIv7ql6T2fEMXF2GdFRcyoWgRMVndUULDhxKDBb
aCsK1QaRBDfbKSU2DVhEG0wtMap9eSSqQIJQLHOP/d0HsGvPpTGQYc+t3G4v7IUARF1+cXfQrFci
jmca0UQZt4l6lmJgCymPdTJt1Ly9ZVXfH9qSw3tm3RqA0qD8b2bpzgBqJnXSK9SNDTnKaqm/Sj36
v1k5M14PTV7ageLxnjilX0erDGN2J/eRjfdj7QY/5HX5O4V8c4BJ705rETr/JfSWGgyjrvkjosC2
26gCDg7f0iUj362t1r5M6/obQdD73WGItYJehcLTJZkWI72Efccbq4BjMI+tk4UTwwobpZcKt+cK
HO0Nm7CYwdnbb7d+NhzcCqME1w5SkKFytOWoJtQ5AhZPGtEcnP/WPWmzH+QskHkvOjCd+0WeQukt
uAPJGywLd/yWZ+CDAcyV+h6KZNsWu0DiEZ0i2EAfavlIBzHsT//jQIjvjsTWdF4NKXaSonc+Me0F
2HDQsX6nS2pmnlxcdgEYontU2u0P2+b4diRbSdQ8Q8hmAWxfzmIkMOoUMsFyGD/nq5OCcS32uZ/L
nZcVGv6/f6AsUyr+GWMn7USwZp3scjmIxCc2t9kjx9O9l5NqYpdr4ls5NUOEi8FnBr0k1bCXCbRr
RGw4hVzxwTBOaj7YZFWxW02xe06rUm+aRQQQT7dYEnmlsTFVIdprCat3NLNiGt39fV7gbkNPRfTZ
ocdeYvu+kgPYLpupsuJb52ofN/eSio8hbJ1jI9YK50gkCfou+QFurbwtEY4u6KOEZHQ8/aEv86De
oVDLV9klB+vpRuneQ4TKvoBZYzmT54AwWn8NlPZYj8frbrYa8wHYmJ4eqTaI2fZaAb4qYyK3lQF9
rcItuS7wTCCAuvlWOWFJm9j0Aks7lJeE+JiZF8leMInE8h8uNCDuYmkImZIExld1D0DvfpmSWPL9
DLAFLkNrMF9/cIKB1JzSVH0tQTx+zc5DEFyoYbi6M8RRJ+GiP4U2M57SHi/VBS/q5Yp6nIwTmvBb
EAgb0N7E4zsIe/YJLt6mq1s8FWyMh2FjRyXEmLcfa4qMZu8aDKYYD/ChBCgd1LLdP0w8uAuCYrXw
3/+0LDXe5qOVCTAk/l5BvuhIHJdIKeOXWt9WZbiPSakbgudFIWbQ9au7OYDES+DWIJUipLRpTGR6
in39KJ7fTCj4KNa3/8ktxgg+jrepE2PeIAL85hH71DKQzQcsCcKX9me6cLWhoucTKRmQyb2LHkhB
8uhm6l1GBmEJc1wwhL41V1jdWy0dquZxxAAuQPRypzy+D6BeUVRqPlza1m6/PdAy3u4oio2EAmZN
+nYmeWZtA2NUegKUikdYPHoMJpAC/hlCchDYpth3l2eqhU/MkEkizjT/JHXl++3QY388dRiRInmo
/mzKTUJlko/P5KgGsihe9ZPs9ed/ThPnu28b+RxRioh9KsDztZu6ltFLU8CecbVIeBcOzEzhD09n
yVS6I8cqMi0t1ijgaPXpsb8XDDtYcrWxkXbzk1PwjOczoVzbHOzTkQh3oZeSHkCiVxeIPCLH5MrV
flhYVE7CfmeXhV99XRGh/UJqohqNQR2WX7n743hUIsat6fWUhaNjdJ4AC4GpVm/SS5bV/G9X/6Uo
YTiX12gSAZ+3vsyG+9r0XXuyE41ReiL3Gn5fbjTKBFeSVRS5NwIGXZ9E+NJSc4zm1eb1gdbnEzJi
ALBbov8coAB4fZ/mYIy1vzTrFEt24UHpPk+LMTfTxjfUZJkPBL9KliL2UKGLcat60fgRuHoUV3Gs
SKdkr6tx/SMa1uvCj90MMcQIUu2Ac4fH6YXUuWoEXDiswm4UHfo3qmjVaOMGKoLI3IQQSPA45cTG
jQOzO1r8y80MYEt71ejplpqdRnLOTlZWRXEEgh18Het8r88Nsf10upDJjmc4czuqwsSrALBMzU0k
wCh5Q0d9/o72SyuNPYDhGKy8GaT71dBbQzwE/oW9azP/zlZHEALJ782h0d+RucOawiheE8P2Z4Kf
H3sXMSq+lMWI4quaV2cSCe3VTVQP7wwe84G2gf4O5n5oC6H3YMmQjfv7YaX0shpiEmhdToSYG1+1
tGpl77Gq5eDNzCWN8aK7FfmK+rQ8HJ9PH11/7wMI+R8kJt96H8rSWN5e3dSFVD9aEfEtt6BPcQfz
p3vN1bdJumUBFvFecXt8OsTbZcJmcmw/Re465qHvPFubFVVTZHk/dapS58kZq5H3b1+7ZsE/vTu6
wqa1A+89/RfCdzXvSzKXdAVAPJugRninVcleRF7+To9xaWwqq6rDJR5LisuxOhbikmQkzYcafRkX
9jCnObb2k2dXGpStHAxXmZXVrl4mb4cNWlv/c4I8+QCHql3oiy2kMEWrr2Vrxfnj2FZq4NYlQ0HP
LuNC/HA+rOlDZokp7r3R7RCQOokiNn32c3mOkdtJYtzcFjZ4kvtJHRbkikA4w28rqr1XBANxWAkT
XJRBpLVgLh7Op6T8zTDTg4w1mcbAV7BvwlsQP92VqfK+qQ2wP+By6SRX5+c0hWudUmxVRyA4/viY
WaM9EVfm5+0Igt0GsSARP/Yl91/qz+2YjPjsiig/kVv9Iciqlxn9MciQVxvFeo/HeVPZMcN6nzYM
6AM4IZLM06Sy3V7DwTWlXG8zJzpXDcjnGWtEWmL8Xj1v+mvY3QXwJX/6BwQfMPCstVQEKbpcbmQq
JJJtftBsdRAWww6IZ+ZP5pFldiCCjCL+p646zVH4sA7r+sh9ISUffWYYIoD4x8tfXXuIuhZby8A9
kT1I+Xr8fOAq5RVazvAg/OqzrXQqNi1K9Te4HaHzmm2iUotsissnPKWqSk5icTGSGzQAsxEKtAVc
IC5MDE3+Lj2AbSfYgiCSaNHsMs3CDrzRl2SvTtjkBDMmwko9cRKDF8HHpwzuMq0HmpSPaU18jX6Z
UubM7HUOmeJYs9ElutY230ZhuzdN8lgFQBKMgSeOqU5evsr+qxHJ3NK77kuMfuQomnuJE2D124vR
ZifUZI6rI3oG+ZurZQlXzTPcMc5VZdPBLbgYvvVIol0MSbZYfAhOtUESxe9KalV9kkeitGV/ZhRi
o6IK8hm2y9OgijitfRuYApZfILzOUv52TzjRX+AIKcad+WhxqzRNTCP/lFebxr3NaMOcoWb1fp0n
jngMMTCxZgKC57PaL87mVE15DGlcROLXSb1/53Ps5jh/vkzwzoOK8ckZv05fnuOQaWSbDn+FlXV/
68Q5QETg4hOnQmjsaARFcvkMUK5eDwF1/GAVw3jeFvY8G/3Pj2Hbl6gvYN/sfnVL9masA1nl6Y6y
1Yo3B/nKFB1+qo994OJ6Ubw3UjnePpIHbtk+5/BZuA/eLe1aR4bj7y17dx7w1gohNAcvYR2crRbx
JVBiNl5C7xMamU3z69oJ5XH/+RlxF4bfrVieT3j7G3Q/MIJiKWgHDVjx06Q/HxvfWozDKqpVdmgR
JlTcPZunhf9telyyD3/tXHNYJthWY69h841mrgTzJTN7SzpxbrSyfVIh0hwfKlH2t383MsAw5a3o
fX1qoiGLUsSlYB1bpoqCVED+V6yPgyEXK41hKouxF36Qwa0cg3ja/8ZCHdXMNSQ5o43bQ33ywgnn
65/AOc0Ohj2dKsEOifCVGY9Lgipftalk/o/KqpwjxDbPRgG+ehlJhtVkycLQK1fjEIf9ISIsxOpV
t9OS9GFLwjCui92tM8JpPV61y5+BhFmTUqRpyVas/QwSaCsRubaMM3YstFUzWvQZypXSsNxmSUWd
7Uw2ivHBeoya/ExtPVe3zrqSfjBCd/KDFAkvOI08ccM0l+n8yXo3qlttzbqNI8o9oIRsm4q2Dkh+
bWNZ3WNEtSq+Lxr9kYKMHjhzEH0wRW8RgMo1HnFBeLz1FHcDC5NIs4Y/EocMQREqmSG4hb1tVGO3
V45rOGaTYo+wsWZeY4+NGaPljoREKjh2L04dMWZOY5mvLzAlKqntV1NoDNsqlEN3tOmjdOYo2kx0
ONorYCpc6gb7ezC0WPI4yYwAP0IjdVBxIBMVlqxeiZkJ4+kvFvcUokoboR62mA/+j+wu0iQNGdDA
+JKxZGRi41AquSu0yy2tPYtgXtZAMxGbE5L4RyoTKv2R/YitXwjQ7uQKjAqnmY8UNUpLe7jq8e+Z
RE51K49occBVaZKe+EV1hR9Nl17ATDNq0qaJXZF4XZXkoU0rOjcrhNYKy15tEtTeMOzg1wLG8VkC
rnOuoNJRNs3PsNquDqRCpcoTv7npVkYl94dB6YWJhAo4dOmHjbGSA26CthyV0OY+HDlZr80FX1fB
3uJdd7eRlOcpSNxhFcQKO+biPxmyvQf9lMDvz8v9M2p2Sp0brZ13l29xt2XdZzwAcoilL88H7fMm
uq0kGPHA9EPAj2cMmgpeDzynzb8QKZgv53HfvHYvOOF53EYnxwiaMaQMPVjrXktzZ1y5Yc6ogbKS
J/Ofe01UpCA2cfuor7rdmwidBtlUlV1EoAVrMgnbgto7voexJE5tNtMD4P8O7KJn4OMNsDLUA7UW
CKgfnJNbCBcNJ4iVSD6XgXToMBmx0OGo7PD8CHHwfB9Acz9mE3vgS0S6oJTZroJelR1lRKJLdYCS
GBa6cPfzynRGIu3sZle86FAERfr5IgoAB7vEF/RD812dPVX84w3wt7WXwbPuzyLt/aojJALjZZDb
LnwoiXonza7yCTb6sA3sMAAwc924bs8hhhekDvPx2AMgVHNFIUzevf8YeuYaB6n4BUfwp5s6aBCQ
XjdaC1pqFUpnxCQoyBQZ347uWnZKR9CZFI8xh/dbMUIFOHZZ642nlPrDKip9A/h3PA3zXLYBufzE
hRz7iMBA0FgjLvrROX/rqO5SRwE9eRawykU3EsHWraPb/MZNMRVaAvaiFnc/HgpXOTtRC+ZWnPF4
wTGjyIRDY+HViKCc4R4TBzi5AlkEs4fEKyQzTEA/eZNUjqqvlg6xGkQgVlb/GOQ6xd33pa1NyB1p
ZVVqijJZ7BarmJzKVT7JsTiyuPhLhbnLLATq90ZK6E7asG3ghR5JC0AbsC6kSublizU/943+HDHJ
hqmBLnI1SGmqLc/FdmH/cIkFgzOkH1PYSF6kXWklary91r+WyZO+cYbVIXUp9T8qVLS/4gdKUnf9
69O9bLIPPVtdzZ93UpT1rV9Fz5VrDar4CFu6WoC/+flF5MxUpIiyB+HlASUDOx07Ahj7Kb+HWlfk
1UyIbw91NFcqx4vRHYyYc4GeSjreIo3mWJvnvKonoo/+Hi5P5Z3LqCBVSyfTB0fsDNvNQ88CJ0xx
T/nQEumBhRVtSTfZKe2xiQx/CIZPTH5klv6y7giMSypGPyRsrEZdxMp1XCQxGtxuDijX5CDb5eFL
0OJqaG146xb5ZXgMtlosn86nQmoY+zifjyg56tpCzujonsqbzpbUertlQDbMRw575wHZ/QrwXjz0
MiIKbSq80ht0NqUHeh7KZ7xrCnsJ+9Qhc/adEZiohuyIaTUo6CjH/lm63cBwM83COdRsauLzuG4f
1ZhW/metK8u5/WKpOltxhcuJUpwAxXfx+FaNfsAgm37UKIabCfxCswTF4bi4EFNoaH4lTFTMIb4w
8EAOv2IwisV3L1nBCWXwIxKWfA1mwdXxXyWAa4j1KkQd74kuBCdpkg7Yn0AJ6R8O+HP2z8qcvpNK
0EGV/7o3zG1cuycODYXDjaVdlMBSvBUcgh1viuyQyQbFkyZP+7Z2ab9U8jOs8gqUCmnkms5fQerp
KlrYO5PXYYPoUpvK7w/+kClika+os0rjE6B0BVRgIVNqvO4UbFz1rC4FbGq41M0EIErjrjhUchgG
0WqB2ciyGjGA0dOd8BqhUWuTUz6h/cM7EPrpBXeZ455ipDPKxKlao+c1dB64/M8skkHfVuemP1UK
4kw/9G4CvFMEZM2KYynLUFoMfiQXNAXKJTLYT/fpwU+bz3T5vDN9/OVhsu1BwxvQVxyk4PGCvtZV
syMFC+SCPazY6HXXxygLIHIC+CoUCCc80I1v9I8ueMkljWpbxyIhmLMTbqK3cGQCNSf39PxSEPMJ
mpthxVvOH4V9OAv/iA0ECSGg/p7wKwtFtwYlJXQAte0Yw89ByqM94+iNesXzkJRchvzug+PjT44/
iW+oKemaEp60c8CvtfDWOtpm1PJKkIryFdnqhDhcCaovhy2o6SslGO68uAee+LeYQ7fWr76/uKrx
yhArEV1x/mCN+UPN3s3dv/2Nd/qXgN53PelXlemTQuY6SS7NXTD9ktKWuh6N4DDINgCF0hYfAyNI
oIzwiyufb/z2VL+H9ar7IFJt+15QymZPoDd8zG7UTtzN5EqmmU1Gd1ezASNT+8ddOuMf9EH278Y4
ecx1ZTAy/r/lrtQBHOzFZae13N8gyc4U++Jtf0jgarMkjncneHIminLNdAG5RzVQzbptyWpjWCVL
Er+Zo3EgKjFM8Xy0i7TC7lQFxDknTxuUgaVZZ4z36e7ffpZMCoEeNzeV+xjqXF3RempO1XbyK3PQ
jNqwW0vri9Sa8ID8kWbph0vjZO4CrTMOfMDuITpzyGQPuRnzsRASl67Z7Sf616qlWO9vrqkU3nbD
fxkXPdVMu5kRalmRNdxMN/bhjBVq/DDvILqoZw9nVr1nbCVDhfJ+01m+lEhEyymlzKkCpNrVtko6
QsQXRunNH2GhLJIlEK1FSNK1p6YoObCeCsaNOOUoACKVWdng2cdVzzysq09tutCnSJMb41lZHVRt
UFCeUISVOZCL8LcMJV5/LB14sKJVj7JP3qW1PqwkVdPqy8ImqYR3b3c/t1fgfI7Fhjf9TXItz8LU
EmfzzQY7Q9gYVNQVJzzSLSL35vPLqZMXiqf03EGYxt8ABIakAwtJ4NyyrKoOHk4SDLsfykCmGRga
MSuJ0D7biQ73p9Sg0kL8u4X/QH4Wu8LiffRhs+soTJezSMuVGm3hN6PdEGKxkOifox1NxHzwldgo
imTa4cBLpNt/jUho4vGxGEDN7OWK7GB9aLseBl44ZYEAFFF5rUTxw3aZMFp8R9VyZ8ncA+g/ExsR
wCo4NuBxiRvlH66dsFQMuKaqAhH5IPWTxpI/JeltVjoZfxfBbzJG+4T3fYCoIPOOM8Ut+vQsTmoL
m+rgwrIXz0jKfDTEb/pD7MG+LuLzSSKa3IBWf+0VBhEXhtcdYtjHaaMYqL52yucuEvSO2qyawFMY
g6+H2pTtjhJbPGwvrl1TvmqoktFCxm4Y3rQKvQSOjeunRXEk9cy+4ICSxKYr6eNQ4inDFjUAbhpS
WFsgYCMv6Dm6UB+BRGhTT9XZZaDDg8SItCkGgwH75vmGFD4qY7HJTHqNLFe/HxvTcBIehBjX77kd
0dyMJvoofA9iV8nX97HeR5rRDxN9fxpwcBCEUBTH7NHiLP4VOPifUKAlRWuYSlUrxgfT2yhpGU4w
kfcz+133e8A2gRFVHUHtgqXK6CFmJ1XNYhrkeXkrHLkkPdu0qFhG7Jto0l/v/gshyge0TkM+S/ZL
sgzmgb+elzbVhoqDKOQrbg26SF3AxV1XdfHaJZMUxaWwuCgA0BevJivmafsoVQQcPiyp/hvtMDgI
H2VbKbFAL0krI6WDK9QuMm+6DExbSkU2geU9KtW23Dw/6lVGssRBPaU8hOwP0A/Zd6cLsZaGAiXX
QliH8TEoX1kXzcJAH1Z8hhJo0pQ/oxrIX9SuaWvv1I9iacRhLMmrQ1ZaMGauCMuUqy100paNbfB7
xdDW14Q57GYeafWHsmiJa/TJ3E+W36ewyXG9WtllWFK2Zdj5BoCXZMBfPam6IxoS6tlIdRw2lsAY
W+bVBo7zTy1zGxbAXfRYOBFW/C2TtknrNG30uASE29DYvPON+0CSX7L2EsB79+WUVAy7oSaGM3ZO
79jfaMWc6+jJgQKQjoADD6L74YjBlxDg3K1bLYkdQ+U99iXa9SeqPzPa+cenDMseOgsv/e0ss2HA
YQp1lfcxDB2wrhj4hs3JOCbiUNu8hslm1ETtnG52F68C8PmrEvTVQlVgSNNj9VHKToEsHAXj4UI0
lT42QSSeHzRpyH+OS4OdAbRNJXFWj2iU4ilp+id29ZMN5SgPagKkbbXMU6r9PrF5pM3QHuCEI1sA
dIw63fSoigWXEhiAOsh3sVmRAWDGRDQcxEjRNk7+JWvMtF/LK6r+WZZvpFeFMZsSVuJZrjuJswN1
E/S4MYQlDUEGONlIO27PpIHtpIYHdw/3uDd7cCCRZyLG/z16ONUvsK9P6n+zpM/aHAJYctZe2O5i
TvWMR7+ofmv598oQhGvsiOvw8n4DP/t13b9ZCESAxNsJinIs8Kdi6X7Tqzj8u5DAknbQOi6hwypl
rPzFrXKr5McQcOTt/3+O75gGqTCHbBo/QofOc6n1MTdBa0mBB3H7RBG7pb4BrJ2KyvfyQG6bUvVX
LGHt+iDrei3JMLMkwkIemyhp3BgNn4rmizCISD0+9SmXS/SDYL5d/Mv+liGJaFogtnPU3d2mkmWS
fb02xx3WIwl+A+NpRza587VxXHmEbYUyAyy07E/1sCQizfA7lmvSmkyFhjRZpnKLefXgvakbcBEg
boOz7l18s436DCnP+OoO6v3nijGtKU1si3Q6rq+PlM4URKDR132tTeAKCf3+IIGdkNT41yyVmJfA
hjPL0wnL0lT7SxNBhIvxsi61HgsU5Xo/KYb4Gp7I/s1maIdtbnJVy4DiCE+J4iQ80V/yuQtlorM9
8v6KxBsqfqh66lhMxlraJNtt69SmjRFkwwAAVZQ6/tpmoOkwXca8/nPF/cUC823MeBmiKR5dKHit
ZGnhVGGfLN9BX9K6hMWOLt6JK0j8SEIkQ5Tg+s3Na4dziSmcQJfS6Ng7K55UUcmZ+LYkSs2+Kf9n
Uv8JnGNM7sycWp0ROPnNOa4a6Yp6BL3n40Aczh4Vc8b8X4ltv/1JZWN8mkwDoBm2X+NG/9/BUUik
/3qY3yh9WJb7bNytkFkP23QarkYe/M2xBHnfYJRl7jq7M6gz44sA1+8jIlWbx5yqyalqMmQa4ufz
yo9oIqDU32kkGN3EsKkYflb+9GH131BjAY9wXWNfjCFyKCQq2l8/WjMoAybEseI//LSn18sWTd7e
tNyPTWF9ZnaHg4jGAd6JOx7ntX+RnvbSj72brc3gleIeD0v1Vf5voTm7xK+huNb77XHAP1Boio0/
1xMKlrBUzRzR4icHIURfaJgveEzmlhn8dy42ZYSQUvIgVA3rQZeYsCtQ3nIy1UWQlDP5FU6JF5gG
RuLb/6OZl5EJ9oc8vMpRb+T+90JZ9iStaNaBtXJSPJkgEt/mHi7AEeV6AW1jAiq1NUBsQiCkT8RW
mgN+UVcfoXrPKbgq8O2UaY+N43TTFBPVcBej0ClWbnZTtsFic70Fs9h3Lfj+kaHS5xlsFX/YwsHq
83rMO7SxytNdvqMJIQtPHLQoIoNqM8Bq6VBcEGaN49sD7o+SWX0I8xTt3IhkLsMGSW/OjuMUS3/b
x34oUSnZHq6ZiX89moCndsqr53fhwQ2AJ/OgHkPqDl0EYXbJxjwWlvw0ANBXPeFdnSbKKSa/d5pY
iivw7RMTS8weM+GRfMhiqdYw9ihzpISzDFQ0G4ZVT7RjDwUOgybBHcrNO5IFZw/WdF//1Fwa73Zz
o0WxMSgtOkihb+Lu8ye/zrXP68deN7aHDsw0RoCc4fNX04dVnt0NooqYvakdky3t3/o0xvloNg9m
ZkQfzdhMv+2pwW9G93VqjbaqknV5+aYJ5sa/gnLSQZiLPgbILwGT+/vLgMzYL1G4HCc1ZG7Q+MNr
H/sgtacAX66t0/FJHno38GKhYk8PHgnlKEj7J3MAMsXFK2L9wvMHrs+UIsYzV0aXnL/vS+/sTrU5
ulRausw+5mQWjx9MwfCun9N2O0qaHYUHEVScuMpbJtAQ3II+O40q6qhv3PXTC4hCO8TmgFUG3z6m
p3wFo1dmCI45eF0EwKUFzZm9O5ShbWy7ths/EcuwIz0lcNbUhRhbjVKV0aQDmvgpRjf2Igc4Kgi8
7VHjLoRhpR7bcDYwKSPg3ckAu7Ce7+535fMDf1PHdYGhtZ0avxnvxtzc5a+ZC9RuQ/nmMraIC8iz
wrot7//jsmd1zbWbws7ppGVR9ENPHFUK3tRLB7qxD3J7wL645CxIzsxyZKNl6o8BEq3CQe9dJpLq
szYUQoXvvmrjBZL5x7umvK91dwAYK+z6sF4CcBA5JeTN+w9ZuaCDJn/I46kHMTp+65rvx0/kfUJH
LVbJbYwNkCg2SQpCPXa3zV3brCMEj7omy2SELGMLwnjYv6IGpogFq3Ds+lOBOOUu7dkeVUu1lrC0
4eg/0w+hAyc9yNNaCh4o42tAYVAOnC4eiOimYiN02HWRPnwgkbhf5dTeL90jYgsSWhPg87RZxi0j
65/sskHY69w768Cd+vXyw3i+EEgjT4ub8/WrNT+2uGycdce47cUv4UZKE0N8asxoTkWA5U29udgN
yeAu0Jh4R8K+Ei/aCI3jmUWzDMDV9b1wiEHRnwZdeb5+RNG8U+ADQJpRPPfDCTtMSkBcdicaJh8G
DIqVJhltSaRa9GW27AUXxvx+tMkal7iky7RxwUUceEelqtwrSv3oGdTx197wEhiqPuf4UatVCcYA
ZSmpx5nl9t+g1FSDvah9HL0/kbYRe8/7SIjsETMxmdBLIIb8o/adxcFPD2rtB84KPWXAJiWI1K2I
dHCDKEjiplMU0sDXd5D6EWL1+VFuCT+WPFeCcldhF/HzlNP2ZJYUQVLF56MQBQk6Rh81AOzANTqh
R/9NffbX1+o9iZ8cEO545aRr8fr1ph4EaM48xjN0r0ANNSMsdbKr7MsPuz6kxb7Y3hfVbGnzfQpv
5pBSUMv2W7D8KTQldgLj2VaVsGf1RNBbq59PZvAhRSNcahjKPkqu8cgjKHpVg796Xk5wBn+ngTZE
+NgewadEjPst1iRX9WeH2oE7CnDFfBtC6ENHhGhQcbFspjQKkzaHeAjWKlV14MMlxN2yeJPtxELZ
LTunDpxFk7EJUfiyFwlqi0rFvO1jfcyl2TWljgSrhymbfTzSPzBqYBpoQpMjgs+mVbNy05E/NF3R
/z+JCpP22KSNq6AfYsM0JzwbrffqgmlMRqkTa2UdEOj26HS2pKDud4VT7FSa5SfrvOgFYO5T8yGU
xABpOSA4Kt7hbg04vZlY1jv44XK8hLAzbJkfYbyZb/k4WMA1R408WqcGwwSHtsSJ9vQWLBe9X1CW
RbD/Tprln9+Pp7qBQXbslpgXDPj5kL/uiFMG1gio0vAVyRiJ47eVowEN6TQO6AoXmD9AqUrp4/RE
vk5hBEE0A1G11Byii78egvUJnJViSucRC94d3LelXbNVGNQ79rmrGSuuDnEwJwG8+BIzYh9juNpG
ommSGf6+wd1Zxe2Kv6QMQZQKL0tE6RPrm+W9mtrVluheU9Dagg3D950cvpV8zs0t4M5IbgpAWcyU
6hKjAA+0LDypdPQCFc4EIZKH48L/ST3tXxjQcLPsRCiCaSVat9CAGW1neh4ja3EUi+LtUgsG1Rfc
5MkbEHchO/5j8WSRu79z119mP2c/oJw/IG2RfP8/6Q67mK6QZsT7FD/0760sBMYaxabY5aHmtnid
ZDQ+nQvBLG92FO+HWftSQ1G3eSCW+r0EUdbzV+ZGs7BuVQYePBksyOFHi4jD7Y+kUXUc9f1LVd6N
lUp1rIS+mu0Z/lwmaj3e2uQQMZMJL3Nv3P3Mo/HLRwkKlRiZ6IaWsZPPODM5NunK00Qg0MvH3YRZ
Ost6b6gzHrmkOjpbcDCyzBh5qB42XgkaBWvQJeV7yWTXTlojMY/LBRog9nCiK5BYZt19xDr2DL+O
KQe6D8SxlNbl2O6c8eeY85b5lyJpVhP4lEcOO17sclLTGlGhXCJTVTVv98gcWc7N9f6QXMNMO0TI
D1BctMeCX4xwyfLqTbN+8GidDP9Hu0+r0Hr3O5ln00ivlQPI5VqkhrPly/hgzim9bLDfXcaKIfq+
4fAM+s9XaSNcSgP6z3tJhon6rCzCcmf24/E7YOWKxIM6KN8AI5TpENArla2HJg3pEtzEPQW7kJzN
GrU53zMuwtpovIaktIWstQ9k1Ld0c3LGzuOKAF8xwe3sSk0Wx8jZt23xvQcDRX0rXC1YLyDYiqn5
ZuxQzQX0yPYN73HBrkbGTZFBg4++7eU0l6vQUFE04kUX2kLCWL1MkIPMWqcW6E9JWbuVGOwHkU9x
6ST2JGEBUP4FVwoZXpv1UKSCOJLnRLicqW/SZWPANpOn2z1woA9lrAh7cAOyWIkcPP3ZCa8jrMjT
Fk9givTJ2rsBtyT2tIW5NCkfRiMDL/bzETm9/jiNGA68JJsUfAqAD2C27cNqFnc4aZNjX65hVxiB
nqDzExnOGzJRNmUQSXEFO9Am9AQGuHdUkJg5f2KQFaIbWfTLgPbJHRalE9+pSUezhamAzouCQ4kM
UqUUR9ubWQTBNSASZwrh8Am9kXeyo/gjmh0aT1AOa/bRuc27gShHJ4DIpCp6VLKmEUiUP0/ElRxb
YKN4jl5v3+qx5KWrauPP7VFxczYnq4v2sXcuvrMIGrZPPVak0FsiGn+x+UiRevKYn46Duyqz6hOu
SRdPtmhKlr/VnTPo1VUJKNrYs7bBuxdGDRlk4OpKcKnh53O38R71+hivpVrJ1DxfRzQgtxXM+yDu
cl2KjUXNAj+G7hJiDw7xwsR4T++nyN+cY4n0uslq+//eVnBQD4rQfBSRu8+TvCebvQLxCsm4vs+P
QIYkxXp9UWHFIux2UAvmCny6KJDQT6ZbEwuwrrhjWmTLL7JXlPofS8oFN+13gUEsKexF49/3RcvU
Ijg6O1TKk825u9mdEAGN0wuM1sdw61dcQ0sNlaWdXMc2gEot4QLkwByADf5yr+TIPvNEb8POts59
Bpyu87M0N4rhu+cqwlkpOIpNuO3/5E012HZTzRCi+hmo5Ccq2R+8AxOzJyyV8pLY0Gnhw858IAmP
FsHvGCY5/CFzVmf7PQWObQoHLjmaUiNaAkrX9sdbigVFqudfWDJW75t+efDIo10lAyqm6LPRjqCC
dDEqYdut8Fw8b9RennjMWm5/9B9xBCWcfcFl2HF9NDtLBM9nm+UY2QKklvpuxW0+NWWdpytuPiQV
bgr1A+ekxa3LaDQRtPqNL1+V0+i+4gjtJRezrxSJAemjqRKtkP6DqbEujQUCMiRHCcQ68nQZfpgR
+XHFRtvCfeife17G9gBuyTiR2evWCd0ujWOm06z3W5WI9psVeu2JaeCvDf71ULMYmzN91yBKTTYk
A5wyhRPrfZyhYe94/2MYBR+TQ4AsJDBA1g1zVTZZwePLrmabh09E9RIYjiwziFI4lG/4AU/YLydg
zzWhVJm2Ifj+4QzWAYwf9IZnzfQdcIMMMhLS2iW4Q8FMAhiPLf/MgrfcaKaT3o88DR4tMDeJkWYf
XukW8ulcZDSK25m6AgmYxSq1zhlzbq9yaYR67WhRO7u17B5aTn27CE2hPl+mlRtFNY9t70uY7zyF
E0WJgCiqGi/9I6EM9Nev/gOMBqAXakgY3oYN2jGgX8/jifVmvl4uwMvXWGnbBLJ36fA5BCLKEFC8
JbFe5M+KJ/9GpccooquVIJd2rIsJOdTlJT+Yf0qPikoZNSEpvzsxJx2HYyjPhBnofBKqiyHOKcRM
f4eE27apIge7lwk9SYZKIi/A1gS8cFw05muj/Cj0pdDeuIhEINHaPpf5f99ULUMpwDTpCUeN7vSP
4i+yN/WxxVKyR3G52Q7giMXqqbAZIy9Ms9DZWNGydCJ0fMSR5Qv2EMEXr6hHJ9tmVuLCBayFrxgi
MPLfyLW58UQ1+ZcsLJFY2KSlJ6zZqZh4AofZTlQmuEZXfVOsL1QeU9xPCIXtqGxI9xnxpOUES2zz
TH0MJdHjnRfqQL4xAv6FviMhJv/tUhNFt/ynfDBomfIaEFIpSSs59DycUFKi7nZr5iCiq9VTP72Z
4GGt1FiAtXvi1uYH5BFvR58fcMDikQMG/Xho2JLOfW893wE4h1Q/PDj553/W0Qx2W2w4ZfvkgWW5
QUlSlgguDHrXZu3HoGLxdHYQw6EuWY4X9JQoW6DhTIXwvRkbbUrifuRoVeOEYBG36kzopQWMVDkz
N3ZnYF6I5O6otJlabGeY78heSzpQMH/6IXYSMvVz5J5+GQPeI+6tnLrUnlfmXuVWg1Zg8lWJkDgN
Z3pGlH5HFDvQ5fQdVOYZDUwgq5Z5gIPvZbIbKlDd3tCmK52gGwsqg9BC4FcXZbMSl7a/gfwJ4mOG
2a9lWHLvhBykREwClLtsJGXxt5gWZDiRsC7gCibKhTx8ixnfCbeq/HN2QQoAtWecjZq0DkLyL/AR
DD/pO/EY9KtENuTuOOAvjHFf1/UfehW5NiYnE+IN/oi7KQBsymV7/osD9DobZxe4Ma+/siILMtEM
hb3SxlryJV6s/lVGYdgs9XLF72ef4Ri+pxqL5Qq4xgmpvl+VoZVmZEvv6oSOcQS37SgKUoWPTMHG
xXER6riqDXBA5pT2nqbZ6MGJV98wX9EhGyjQa3h/YDXZgNSOCTNhSUkwQJdc0sZbtVectYeyv3RG
CGtE5AfjBzWC1stDHd6tmjtJb8UlvOUglOt98YEMN9cmrct3Xju3C3JESaHOSswbZg2xRZ1fOKFA
bSvFBUBoqTcnHbaj7PyOLHLGhp5YSAWfXCBBCmsYxwVh9NvvC+J25MWoPYeC6ZPB6gHBVNj7uaCu
/UoS7x5BsdeFnnxwy9cLx1HDYVu++7SYh2eL+ThYoZf00WzJu5PlUdt3LRgcofe6lAtLXTtTk+A9
3jpItFYadUksC5MrJi2/bJCVjoobqxKCkni/oxHwKkK9afdCnJtRchhZcpwCnc1ii15lNWu4rYPu
iD+uhIYexij2WXGmSznHNCUk9TFOBgKdwp9WCy8SjFJQFsSdm8+Jw/C0geerCNQY4jH85jyTgRQb
dN3PaIUurBmUzGBuJ3VjFB7dmq+4TtxHF49NyX4rizK5CODngd9L0AJROH8eyZv28WVICRuRU+ZJ
sjA3mHs7Ety1hB+m/Pi9MVgP2MTfuBi4pAoiujBR3AHhnefxjGKIVXsOdxQtrDuUtBrHrOeV85jR
CFS2vt9TqTUDnMtcbybvJ85f4N24obF9Nu8yrp8WWK8kpx1oChXjx/g5M+AhTNAlwoTFqNgy6PBB
Yey0w/anXxgQjw+raLds1P5whFtz1BiqEhgaCkDwiT/jJ1oTwG4SlnSu5hv/V5cahIgmyyId7nTK
j9hM9XvFZVcr/t+SH2J7BkKpQkuztwJO/lrI4SZANKrI47w+FAFz1QJNhplWlwKQQ17CYJtiJqJ1
vKIdvrQwERqSrFSqu919tQDJSopRHJbWJHmIG4clwipUfY0G2zEkjE/c4sybigySAfh+JAcRKFsh
CKTtegorIY0EFuiJGYaaPlxndd/wezl3/l9TAu90QVTcNMBvX0yeviudKFXTjC/Ca/wdd0S2TmJC
IO5mfEOmwaEyIu/zYRGoXaIw9svEdBYmX0CqZyntKDyzWaX8/W9S0E4xiIU2yRRsl7yXBD68+p6z
jnQ+rvCM9IgRaIYb14X5kzLP2+eGTFItS/zuwgkPGoc1QCzyTWAiSl1E0LPgsaOQ5L9q0VZk8C8L
zcMlDAxImTo5LHLqd+yybpUc3D/MP125cxLhk8sbzppX1zVyUf8PsXg3CroTqXLJPeUdtp7IuzW8
eZnItOeN1MNvjx3MUE0d90E7iGdVHXAgSXqwYpWaAqKH6GgMgwYurNVVr2roNqmn5+VKs3qfBjYN
aYnXB7lNbyMltEkASKNGCk52KeupQOTmCZD6B3b2JHLedJfyuN7fnQskRUSchVI+Q3pIGV50/598
SNHdzONC2tBSJ/3BGDd91/ilRFFEuyYiMlAivLCoQKU0sDGgtED1DPbUcnWwYCC/z4z4ja15fblY
cdc+hCU0/eoRpN8B3lkugVqp1Z/sN9j1XNWGUb7hHSUYfPbL7ytSX4x+2sbLPq2NZY2Gec2iXpsH
EtPaXVA1q8M0FVPoEm4Yr4JbFIUxeWWDC2g6hqs4Q06g2ys4vMwBq7H9sCTmPSMaBdsouM2WdxNv
5tT0/peN/jWQ2BCwTaMj7f4BxHRJir6BpuogcpfkSI7OU1BvuIflFQiCZ6ETVO1RWFwkCCBmYKn8
YMUnfaPtKaq46K5hFx2GzOb5IzjpjH+kXuuCm841gaaL5bRYaqA6ZsYD6uYfQ4U4GE0hFzG6q36u
sOF1FjzxluqO+eXJfQhu4l4FL7l7woghknoJgW6Bwp+44+84BYzLVRc/gy4tC+BOaiHggcxu7ZZi
e9MtlNOudm9iXwm86HuxB6TiL84oXLjkNNYCqLjEoJRFduzEmVm3+ZV7LZeVcXrUrkwiORI5VwGC
I5XGollJqA+oOgXWZip2lbrrW7RfJpDPhPz7DlO2Sejdn1FgiWsIWPsai50Yx/YM3+g+jxTRRmnx
lZxxczINhxy5JFMQhu2j8NtBJ9BS2P3iEE8stWjmBlneEuwX9rKrsJsi303KTO78aaHhZc7+MLeT
kvD+8d0+gARo2K/0dnzmntvoOVhRdSQ1tc5BkaK8rqZdlDCxBeDAjZdyNPoIb4cNHhCgZjnKysMw
p6p+jmRYHxzGWluV95DkOKKDOL1nUhJfqnc5bOj5KE3qHQ2ValmYEP8gZ2+9ddN/HuHjlEMcBUQ6
zKyRxAXBSBDwhgy33Ywk1CJcae42RBpmd1xQ5OTKzPl7UGbJGdEJwzVD61IBm3F20o/enVY1SBoR
6LkNeDcQpy6lUgMqVt8s0upr8N9iD7htaUcd1ddJmLyjydh9achgV6ZyOzWHwH0LTkvxQ476HRlh
uFBC+FNmseBmcw4cYhLxm522P4J8CuwPl9bqMOqSxplwZvG7R5nfy3FJX9p+BIElqK56v91sYOM3
lvp3fncwKViBugaePdD/VOAcXzs+sW5HyPulPUoKPFJtnlxxFlJUHMq0m2vlsrFE44JA/XbIVuFS
Tr6BR1ffOo5TLZH5Mta42iBdaOLEWgeSZ2pXSbGMSFz6Qhc8/E/O1uNlWpBjidIYiUZZ95kK7ynS
+8IyMof6eR4RxjzF3InQAz+6dk9DVj79r2ZWYK4JH2tPLNy+qbkg1fk3lVIvHCYIiGLXuOcpc8RG
eMSGYuMhYnZKJG1M8OnVk5l40iIAeazHBQSsgaUvxJThk+CUMnWVi9NBjetc2vYI909pQFnw4Zlx
9MiOOSSBLPyvfQXm3pfRjE02IyLnpjpfwdcg8EAYT5Ib3EjHZSWsFFEyJKCEiv1nus/0i9T7zTAk
UQJPA8Gw5dV5kKrFpK9SVZbGvypexb2G8WsRZxr7bLr8r8cN+ZMhItW5TsJCH8nY9alD//U5GEWf
sxkNjjrp9D4lWiw6DaUMwdBChXOI410RznYYoMxEy80zuHUDzm/Vk13xhncT8iO3PGR1n5L9NjC4
8hpVOpg2Cxl1IrYF+uRRD8QUjVuw2KUXKvUHpR1im6ocl0W5ho6rtmi7S6pUZmyegJdcF+zoypbm
R5UZ/Ke6Y57iEgr5cJn16eS7x42HSxt7mHpjBMOQmegVtPwBCx3j2a6nGd5MhbvvyQUM+S0Xhtg6
jPKuPKiWQmF7Sq6FHAcrNIqFE4ZYmYAawIb4GR2Iz3FQWlLRHldsln1pIiWuWuCQ9x1tCF3vZ7qN
o+apUuuXVLy+oCDbAJRUASgXK1miOAdtQdU4f9jncyYkYaEYkep78AfUYe7pVyAD/E707BBzP86u
f6rooAtFJsQx5gyLnXpHcbCzTci46oDp2DXIEG/YW+IP61p8tvLz8FN5fuXuLTQFXgw3RhYzmTei
neI5hnbHf5KQuJfRVGQ37GRkE3kVwfmkidy3b90zn298umHGhujoOwK9hQF6eI5MCcPRmYDovumA
awThjfL1C2DOGI7c/yPaKVm174Oyn1MAZwIb3tCsJ+WVnsct00pBxMx4EJ7jTAF3h35TiekLYhHQ
K/m2xhnsnIqRsMlsLtSygjHVIES+SzZiiEHijp7pjDkRiYYPM5MJx0eI4u43ZkkubmToGA/nCIdw
bCEl9ds64Y1UFdMouaL/nm4zBi56KFqo7ONNf/JYzDuMjXMpSidoQXJ2LBHMrG+TQcjrCBTrJm+A
xdGy9BcZVESCwRqSzPOVuTa/jYwK7Rj59PwJXTq39N7yah7FBFTX2Q2oOZlG4Alf6NZQNdPqJB51
i6jPtTpSJCY0NsnC/b3RQl0Og8H/mc4q0ePQrY68iMk9HEWxIK8BR7dP/6SfoJJlpNKBa5Tln6TM
WpPsLjVFtlWJsOEBI1iP8cKkNYT4l2RAciWlWMRdwnhw6EIk+RHYNLGqnXydwgr4f3nvkKVHQjPV
R0nwETg94clvDgLHHCTpSNFOm9xM996JlPW8js31Lf8okF+KA/Zz4HXZqzZvk3MrZrtpm5O/KSaD
cRxCOM2PhZCdmaMZUBfxYqnd68lsnW/Ceti4YYemfht0Ey8eq6s4/Ntiwy2CSmsRHMTC5u886tgy
4noq+qXMF6A9g2iw2v3rAY4RQHaa6kckwUEaZMDrH3PP8UH3geUqBt1NLO91px+Ren6iYpCA+zW+
ccDowMKaMeoz3B1E8Khlr3fpGsYxhMwqJLjZw+qBsCa6ZNrn4h1bv+Bf9SyVSBZe1hdjLSfjfK0a
UEZwMvfnchwMEdoO5UiiYs+Lgunnxi1rPjpFQSpVQF7ztBx0Ae+TN8yA9LxKOuro/KW3ijVI+evT
XDu5qGXeanl4ydNhVQLXRmrjOs54fe/rIBw6M9ZBfpWx/8OvSDMo4+NdrXGuaYco62x7l/RryMxn
/rpSMUAucmgCjRRheqzEU5kjCe2cefyWjtmn6do/CC1WRN9U80BxR57FhFwZ1Y+nAg5AAyJDdiKV
W4uxFTPVWtAQlHauieqH4Q/XCQt/lWzpwT03wKqe5v+r01tcsPrG/XYjhI0O567LPQAsN6tm5LZ+
n15G6rg548i/Omzfv5ZJ8Vz1xhxuKHz4M68rGuvZuas/BmaZDezWV822dOxhnvqq3TFhLBCySGFq
pOswTEb5eD6Ij0ibJp+KATdluMdXF4xgxgwpHcpDOiXbiFj8q7i8zKZZt9h6AOWOjsBIE44uhmjg
VZ9hOYW9JUvhzPp0yL7r++lR6oNM6PGmLeqIbwFw37SbQjcnAUh6KxXOCPtZTMPwqXdoaHeyrgj1
QgfMrGB5vfpZiEVbp06ZcfXJqOa0UpaGr7vpqnEJd9g8efgGph9haXWsnmxk9+ZhPevm2hNB/FnQ
H/mJCE9N8BrNBzPEhvVlRvahNJbVUGG0s95K+z8FUbSFRpdH5e7SGplTZRRdsakX5TZ6VqqyblOy
Z3VwMXKngQluEEjz6EwZsKEdh8X5PKTfBgNkOFMgwTtA8I1BzOH4WHXx5l/ThW1pPX1eAfgPwpS+
ltGcDfLQsv1V4+6IrcEvNMMfUaAWO0NQexajvrtprG2fIYeIkWYb7Hv7vfkNDQxSkMOv7woqbcBB
gzSonBC6LwDSmAs6XdZCtu4dDtRKz+r2L+wBkLPaKOgKAI7xg8h6y7+I6llGMKyjQsX+w5pOWVkd
w8D95uYcgSAw3Gdw5dFGCZoMnfFctU8FFk2GMxGKuQnvEOIZ2kyxZ1UyBVwjXVYCFncv9cDO945O
3s1NMlLHZTx+tFN/hv39moY7CHn3JwmKthPnClynUyHPWJXoVxZNVSy8CuGX/558HQfZ6RQpUbAH
tT9AKBTMh0c+KTmiQ91D3JrQm5S74HgjKZWEH0lLKOk6nZw/RYKnFRIF0lQzdqBISjcfl1Sl5/Fm
N9uVBQPIv9QwerUE2zxpwmAm3w3vmaZ3SwtrqA6LfWV6uj1cwgl/aJbFo9hAJ4XAf+ASK7XEjExR
drRhCkKBmszK8hmcGW5SUAHB0s+vmDS4or4ghWsz4K6uvqROx2QXGQe8zIS/eWTdd7d0OkqFwtEX
EKFW1ucf9IYTq11hgJS2+CgHymd8EUngic/f2910S+Y+ciMgsUmtIT9pjFfUo38yLnXa2yHN3Dif
FZGTSvum6lcmx8MKrCvECVW1spUUN3x9xAt+1XXaaS0Jhv1GfSD+5mRDRrandukmS2i2JupmfgFQ
sbH7V6C0Mc9FVTjJHL8YItBwskxCqniXSlC7DZdTPpoFL2W2pO4FZkpnyNndhMo9f+sMWvlo0SGB
o2iWSwmbN92MmGnkiz29/376pVqecbA/ut/XkllMnA9A4ZaFsYTvqi/y8reyMxNbBQaROMvDSw1V
YNV3rEMQWf4LGl46D/tJPC2tPyTqWW+NqsHdkPUbL1NuJsyMYDlIoYBlQ0PXmTm8NxYrCKBnJ4of
R1n11C0cTRwDlhqdM7R/ahkANQy4/eZp6hONtBINJ7VYgK26YHeP9jaeszj2lZqRbfe7rtIx4FgZ
WYdviW987vkhn/7w6nPO5AkaZ5rRsJxu/r+70rAw+Rg9mVvlx33U0SfueZA+FqG4Q6zc4tIdyGC2
Zv6cjiWvELf/cQpzcbT+mmlCe/OMxoyQrkRahY4QX3zXu9tmjoHifvOTTl7PzcdVM5dggNgGZ9TZ
gEDl87ZA4ku+HS3N0jo1Kj7XA9jtsOJc774vt5cORo1iAEtuA0Jz9gdAFquxNXzP5HEkpggHNniK
5o1z7y7ojvR57TBwPS+D6MfinNXq/l/F9DEtGQbkAuhKoGZhb877ZUhc4k/FdAFY1tQsMjX78TXB
zysiEALOF3gLx9qPnu1QmamvEo7umDfrS90Q+elExLs/uB/9r1BE6A04Hs8HovjG8uh0ZXfgrELr
T9mgQQH/2EQxGXTFDw7M9Zxa6ic3LNYx/z+Od+5BQhtGs/nFAJ4otdReVEYJMXWY0CYgdbYBUwcz
mFYc59XKl38N/9+ntX2UmvQne6JRInJBkvWluF6cF/n0Q2RYpmtAso0Co+VJTkYgkEofmihnl6Li
pEVa8lWAYTkx4N/CWar7yC9pq+N1ffKMdIQmavk5F3AhZ5ELf68CXOxPcB68BnO8idBapGcfSX/q
tntb8CFKmFnJM6sxr6qmCna9zPypvoQrnKb8Np4RuR5xL2MNGjwoiJufpxpGzdcU4hGw+UIhWEIP
4dAtOBgzp41hIVwxYtXo7oUYHE3fHig8civgiIXdwMCMSiGqLDvUzIBUtwlYEabuwQLTKhaTJgZ2
o7hpP37m08a/f702l2yz6YR2fSIno/PgA1nt2Y9UTBxdkAzjUcGjXRagkXbdOrloq0Xdd542LYcz
qVFkBLayrpKACsGkfJpxynqYmHDaxXxJcwXoNO4sWpxk385wuN2Sn213/r4quWh9Xet3ZU+2OixB
BDvXj5WWH8zirpfxILWFfdzWeOvPB+8CZ05KsU1L8cA/gZrv0mRAV/Yxq7US8Pp7PMlqAxIVvcNG
U3EEhTodDYBi6TyUoh19vTkQp3j2UCVm1P/wK34rgm+TfL2KuX35GDAmbrBuYubgS9JmRP8tjUF2
n+NlG7RWlk0Yuo6hpxMBcHnrsfrUYuQSC4t6VRJPpXEyK/6BhCi4CfjmZNX7mWltXEnDALKTNkFt
ST/Ok0gJU+ob+10+B0yzNLtNWHrcTQwpMG4hzyQHmto4v8SHXX9poKCxyHcaN/b5cEKYSE7VKTP2
N3xDfCG/almVT7Zj/DXk2PCI6hdF75pQRI/tjr/NdU2Ipdbiu/NCcc2Z43YNqIvqwOJiaq1KjGeA
0RjnPdD5ykVjXfqrTuXYYdXk99XENlBapiupULWswP0UzS+XZu2n9S1V5SJU9GRMWBy4kassRtDy
X76ZbvGG5CfoozZtUeBZyXKABamnbuKxfzaqj4dJGVBAhBqNicpb6juPMmzRVZXSqboaUu1wRs8H
NCd3XCJ+8LSWhSMcxAlvXTXyrHKP+vAVS7h1Xtm/NXfWv5zF7Yuy483mIxe0kWkWm7RPPXeAH/wt
jwBY2hSLt52C0NVIEsZ9LnuAENFsMZ/HhrtBH6Wrt/7y8jhflHIjIoYOL+yGvKSiQ86aoh8Lp7Ju
7UxTG/yYmRff9Go4k2M5xIfT0iEuEkQpzFNHjADm+q9bZUTfTXLZoRhGznDNXAbzGKVeSiYKvJZe
NWSaZ1ebScwL3ZdytLlJDIdJ4UqArRt+zwKl8BgK//CATGxPre71wYh4MsigAyzVnuQsTVXXNG+1
kclEGbo0WbkcG5yewF2DCER3tcqABykpzhMbZimKbfQXjB9HoJq/9saR/vLr/Wj219GNdz8GgdG0
fK74u1a/qxMT2LEK9DJoxGWCjt+D/F2MPdtPDnWz2jMOiPAX8GDYA2s2GApMlE35oW1awbXG+0ED
3Q1tH6za7ndyZFdrDvHlhHYL3O2WwUjbFF9DQA4c/MdMRRn8WqWfAa28dsdm749YUTylGMSHec00
t7t4Dcq6GmgHO+pYKHIdQcdkE+a0MdUAcWtPVcnpGHOJkDjLV+svpJ8PGIQ6XrPoo7rfPZI7OEhy
uuU6G+E8uw71cq8h2IIc1gtLFsEnDIgT4Eg4B68KwETFz0VmYwxq6zvTjAR9c2gPJCfQlJu93JmR
Q+uzn32J88hcex26BBfRwfS/PWPphyQYZqJdFh28GmeE0LqioYQtVlgC5tI1Dl54RU/9LvjzapOk
UjgDUD5KgDKA52RvYs0P774E2gJwx6QivwoY5bsh78mChFxujrtvPfC7brTW78eVAdSlv8SmwxGA
ivE7L0d3vP6/ExO46ZZWl8SxScREa/xTqktpOoD/Yf1lEXEl8s+bWi/ukyg7Sha3I1pYgmPe4SW3
HkPU19nuSs8+eGqjt27/7eKMjvoemUxahqCLIbHhMv2J7tBSdWvbc88PD4ArhXQCLavnbf1CA6Q9
F1r13SSpRxskJMBJYFp/X2l63NL+gKXmd98gKPErc3f8eMSr9yTZi3Gv8+C8XhIFh2xZkcQ5Drfp
3TuPMeIiHQ19zxtfeUMmrCBYigRQfkVQjLQcTPCAJ6/pGFShQoKuaMHx1K1PXIahn3kdvQOH8LWn
qeYFmd/jTT8jl6vqFnJMmA0sByZMi0cg4XMssnQ/cQJcPr0+8VTiqz46aaUPLSnnv+mOxZ9KR+G+
Gc8gAttwvWbCzuDC2yuuKfJWl2yJFtAlMfuKvpdUWjtu8mQty4lrTnbtclNwdPN0iaOSFtDY3N8Z
5F/nKu+z+uxVh7S6ySyff91fdnbhd4g3EDNI//sVGtConsfdhu5LYkuVqSt7Nj/3e33dWKyzBWIz
p7l1AwbNV78R4WZumRbYWxNDGrow3mfo1QnWcc6w9LsLr4aT0HnNfQc5Xc1oMcSsUswMdn7590vO
7IzCJ3OcmgXrIbnJ9MQDxxj1ebFgTlxB1Lyh51gSLKM9RdgEnkynw3FNzdSwtnovQ1yMW+E+wbLq
Hc7/eZiAsUAn8xyiIvdq1sBvN0STKqOPvyFJg1RtXjh7t7frYrRGqyLspbzLfnppeJsCKuAwZJJ9
pN6zL7l/GEdHXwrZhFrbuq0+BaYQS0Onayugf3X9qkKE75oh4PpRdHs6BdaFer68QEP3beK/e6VW
YXAZPajaUrsmsi3TM/ZIs8TGjBwlGiTFJ7UUX+1LF2agCGuLfJG9oHgHf2rWHYZH69f3MY8PUeFy
kdrlJ/p3yyDaxzGNhghuiu9KgzjC1bUu6imq9bAMLTLRZLv2gXSpfbKvE/BJARrmoPpAPJmmwnfl
KtLNORM7G0OC3lVssYjEZpPgkJ/BbI8ZypCQXsEY7Z0dkw3/QkJTXd+crA7RBp6ZYQVt5491u5O3
MLXydW/TYgbY62TRmlsvcstNNnHNAomHdhuSYZHSPmrPEH3mW91PWctvQPjP1FEzkx2Mw4pC36vF
2c8VwjsRU6MXh0N5tRMFVZ9zJgnUHOwAMT7MitvcpOlZhRCjVyLiwFAYWzTz7FdgB5UKeBlnqiQh
OjNli6bTOXZsT9Kt0ZGQB1VJS19YXm+HQMvlGpJafNFztXLa75Q+tSIN9S+kY/Nx9k++U2nGHIEm
l0b5J1Tcw+pUQcqenWnK8RiAZOsIbgVPEmU4vqVcr7Pn87fRx1zAuD8p1LxBhq0336TzFiLc20LR
59sBUEvsiiIJmtYjIKwd+Q5Oy/qVB06r4Qxoa0yCgW2XHtkSYztQ0hIH/fAEhLot5aIRaFOG9UUO
tAhNvkQ3xV4LDxG2GpNq12LrNo9D6BsoTvuib8Ml9B2gp5IvUHtWstpFALvEiaHb0hEiDE07NtRd
4qwGB/UDHkjR97Ye+AVqY+AcMzYfv9S8x7siLRB+AAQYqaieCsI6KkjwwxbDIt2CVwmBoy2o1txe
BcJDx9eTmI+VnpZsfbQmf32HikhbgZIkBXTq02h/8fUA30E2+GUCoAEubXTz3IS5sYZIqpwB0+L5
/76c8fCnLWcVZepdER2TtCK53IuHjpu6lPTdsfGFPH3s4R/aXWfuzKnAN/UoQD2blNZ8IWlo/ARr
qxl+73STbSWCW5BJXOkHMxt3aGftzDUuOxYrY9Yuioaz5wqftdg1+NLuWThi3bdja5hQzVdDTUSo
Yli7dp2cNqKJBu2mogAZ95LPE24lz13aroMEHmmxSdQQpr7Cyt9CSNMd0j0qaWLU86jlTSL/BT1h
UOVr0qiYGiWcz1CJkTvLTe5X9irZ86miauSQBINH9lFlptXtsjKYumkq86KyeU3GnJ0UN9nm53+S
17kr+G9uRz7SK4JtM/xxJ4aC42BfrB1Vi0AREboczyFJZLeJZ5Oo3d2bKq3AB4q+ohSrPDFYMl3t
vJz2OixcT8qVZkMzvehzTfdnnvWeJXwYBsx6RNYecKtX2EZQcJOXj448y0Vx2DMujK0Ij6j1ttKa
1ig8ynUW8PIku+7fM1WJ7lLO8tv1exq0ZqytQfWR6OUYzii05l2dvmlEifLU3/YX/FqMQTMUdI1u
N2EJMAtqwHf32bBqwNNiJeCPI1xOIM47eaqLMTaa2jtBvSQS1t24aA2RvXcGREm7Rcy/pc12AfT0
miB1EFVJ2ZUgjV8wakxr3tZueV/H5Ba24YaHF4R378ck7QNgFIFDfA3GCtbwaTLnQzYrKGnU9TZf
5x+ihyGDan3hQQ5NURazCAgbk/nk+bkaY9nhS3dxdx2PpHHxcnZ8+8hDaIQiQ35IgwswrSl21bk+
M4vX9v9qGB8uoocjfcmo94BqMWqeCHFuH/SsSqsoIzt8kxQ05nsf4cSd/YvCxacd+H4Jl/wQ5WpO
xMplXhR9o3k898wITlw5roKvlxMfHiUyEJq2+R4I1cv2cvAHPH8AvBNUwOkzBqt2aO5obIJmoUnZ
nqaM1k8N4jKXNpcCS0WkcXt2i+yRgTwbVAhPdRO+nDKpPDWbCQO3aMS0maJAZH13I97SvaybV9Zr
iZpPpOIu31UJzMU3bzVoV74NQ68etCJ7uzo8LuUUyiXZovC2CJJFGp6deKgmySgD25RLUkLrm//P
DdV6vN7WyTB8JNPZ2hqdoSzUgPuUB/RAsbTu4HRNfBy1CshmQVY0AbZ9aOIL+7eRGZK/DzTmUnOE
aw2o5R2q33Cx5SJ2q6iM65xwri54ITWJOW04GFPCD+bO/kMuwCOdE79cqoMoZmCXTHpdZQcRusQb
6eMY8twIhRLSGa9d0fmESDMDwVdMSu/7MVy116uANFlbaRgfxI8H+txliiZn/v3Qhxonn/Fbbq4Y
a+wXhKhi9OBHDHThzBjPWDh/UaupobP+9OIamBBQMLUiZ0Hvw73miITEBfH6918mSTHj1UBpn1h1
5nkOvN5nifKzb9C48qW71aQW8Zfdraw8/uBr+QrWB9YHn3Naizja/x+GjIb7JC5aLZkxm1e96Nl/
EdSHCe96lg68+srrfY0u9v0Ey4joB2XIMSlrM6M3NEPL3w+Wpamv7fGympxmOkEtZFlB8vg9NkJY
MG8aRKTmUILMC2JVWxauxENzV7Au/tCYfhYP9NS/0aWKWf9Fw4YRcEIkJ/WHlwxXwfAsCSrD24O6
B4IzTzLfNkix7kjTC5C8eQEl/9tqPaefeIzSs53cuP9vWrZmbOiERCxVcHqsCJZIK0NXqYvijz6D
Y/LgHhNOTANTMJmim5fxCC5+vA8cng8EhLlKQV466pxaitQySVDIffgfFc8vkomyTcxhK3B8/v4g
9vkIie376ShfH8VQ4YZLcZB7LKKHLpqaHUwODUc9u2Hgsu3uaHM0NCZ+07SKBpsJZohuRg6j+8x4
eEZXspNCIqciBz8t5UYpOGrcd9E9oqnWenyccknJyZE9UCbjCvhpALX9BJ/zDpkGtxCy7h9w48sr
WIPGdNU9oc47Ix8M+CZwSvCUNjASmWIiKYOASUzn5taBQBrCLvv1/1wwkdOpfv4UQiEujQG6tuPX
HjxLy0Bgg05Nh/JR6j7R+47hkK8FY17DtCSxKqcivkBs/ubO6LEHNgD5MUngnPUrZ4i2+jtedAFp
tL63wIOO2q+Nga/facHrTpgbnpLArXux5LaJzvcp7QchmCDfHG3cC7pYWNSne+xDOAM3AznNrHK6
gxojZOiSYkYfQ8XjyAvXQvBy09xqVepH0gO9Lj9CCpWo2THfJB/qw/5BGumHnh8JVG7fYg0TIHFU
sEdqWL6LiAAuZ/d9zVujGPQG4jt/zPzfPoWfx8qBmuO/F2sOkZzHnPViS4D+LDCInwBXmi7KMaxu
0ANNXRoO4G0h6D2GLEoJ6VwtC29rBwEy8TmZoFV7+rLVNgaRzMwsRkLviiedXBkiLkWCZF1AGqX8
QmK5iP+wrufZjUngSbz/AB1m38bRW12Ui2hwNvudHL4ukIPI/bW1Evv6Wp/ZkMketZTkLSYAs1R2
pNh0905gomeq+SXQJ+IvPLio9gC9o9hbUcKnIYp6peqwyGsY4U3bQNR5cUO/Wax+vhUBLs0Dq63L
vhaAG0fPriUknxiisCF9hq9AgCgxJ2jbXdHIVhJS5+/78C65Kd2d6raeWijvZxRVaAQvyJ5fK89X
CVhCM2QaLir9zoe13xT3uk7AAZHvdjXH3B7BCiwZI8Gysqeko/MIs77SKUsImg6Yl0zEMfDMcHVr
PGSCIGPlOZLBlqKRp76wNlzQo6o5iwS87Ab2fvDmdX9fGDX5lqxJtU+oRdXUoGJ1rX7w+GhSIlzM
lm6U3cqzrRnMN0DSV6FmgRCB1xfTkG1vx43jz0aBFaHXx6UmNiVCqwwYKcB6pDZGsoTGk54ZLDpm
X8/AqvtHJkvONh8fXII3IXcP3BsS/Udo/Liwp29HsnAPzskU1VcRi3riVZpxVALNDjzlsMKloH8T
BGDoD+NjABlDDVyULOSSvSPlAq1twZSY2Jo2S7FsVEvbRdOPO5wwXkVqFGQ5Hn5fFI4Dbtq1DerF
4IaHVeEfTy0hsBE3dlBfPvnFRnQRXQhZNSO9itBUx+iXuOU7zg+cOx3PyczmHFv/b1WcgPKjlgII
H3naK0VINIcc/0GdMwHqz8BEvPxFJk3jr7wruswPI1e4Oj31jmSQhOsswd8zsvTdt+kr49KYoldR
fPeW4kQ2a78E+HORA7TLza5b9iOSg1ncGI4X0sFoKBR1k5PSE7/Qe9nGzP26zzRyefjGYxZ9NKfW
AMtFVeQwMGABrr8cIePHcIDicLfAPn63PbMkvbOcaP6w/6fvFyZWs/vezB2w5tkJIKfOTrto5Esu
X4sBfalILEvvGDVLs90MR9kKUzndb5y9MEbI0MC847Mt9MzmmiaO/mNX3AZWCnGxSIxXT1vWRP3z
QNNb7Zrx5b6uXxPjJI2ZlASBg7i157Suk5V+V3kPdwLxOW5OiGbB2tHV1zwIvX9kIxyrDf8Yvdpi
KwnHmvVDxdPLEN5ebyROngu5K7sy81H58JOaUEQ3hcvAUn8wzR4a7XkjpgITrzJfpZf8AdQuXR4D
msIDeYo/KB6Af08rc8CT0nXubYvEbQJBpFZSTJshZ4nFsCe9G8U8/sajqI7EibHEDMQ5oEsXzBoi
t5XaE13eXAf7/5SHXJqUwHrAe1lmkSsKsq6rcWmUnezg9rvgBFL7mtF1LT2Og17i/t+0XJly8Ulm
BP/lfvoUlj3Wh2wxpbz0bAcPrnY0u5JyEVY1GGafrbq3mhHJaNCEujxhtvuNmd6zT+NnZSX/SRCs
p0pQFPMs2ten4Tl/Z1aXa5x8nKYnhheWNN8QA8Yxqkw5mxPKqiSdq3b+Vw8tl+dya++NyOan3yJp
7ssWaYKLHaAWWcOBNGGNq4pMzoLkumJ9PtabvxKWVJPB35xyoDCwyD8GM+V1MU61qSv8zyISwO+z
YRypLHddZls030sddBsQvXQXem8iIw/VYK7amWNFu8S11PNbDONMJGfnMuMb0JYmz33YI5OPazic
1zEOcf8DxKMopKK1tLDefk27HZ/YXSotW/XGeCEcv/H40/A5PJye80iugPnNtNKDmAxGcWhQDLwv
d41phjJlv6Qk5MrRhqXXBqv/KsTuEa1flUUemUZIXu3ov06EdLEYf9QpXCEDapvKiaaE22Td+v62
rTMifpdPnxSjok4jX0E0lw9IbwI5aefrhffbwVwOmIIXdlvbNk6SJBzLT2LDsljBndojP3Kiopfi
UaWPY8JqcgaJ8wazPcgPhEEj+2Vo4PX5Gw/V+yF+yjM0BYMkdCb4ABZHPs7EWSYjRMBTAg+i7pWt
MJmdXRmcsog6gBf+hk9kIkIfXH3VVnJQcBMpy6wUmI2Vhp7fk5FpN4hkjZKZ2Q/ZGVtFjUDds4nZ
1teG0Xx80vNq6aYeNfSyRVm9WAwy139DMaa7NTchzKs24FfsgLisbdM2OGAjKS2+QJ8cK7qH0QsA
CukgEq5qVmytqVN0QMWwm3viTDcHMUEnWgcWBuxd/P2N+Kkd2pSGAtmuRC0faDJF3FNqjZZm2fmw
P/ke/EGhdgOT0+gZ3zJtg/QEXCCQeBH7kRRc98jTRCBt3rOT+BzWtBFT4XQDnicP2Pef9c/2ks+P
ydiz8fMXCmfpO+MFs7VqmXHoACTbb9cUfKiiqoJ+h9KbJtRr9Vfm1GnC/vQNsG3o6JQbk94Efb+B
iXcp7AcDStHjdMtx0ZyZgo5YGz77sQHBdm3oigMwpMgRADoa3/3aq8NaThbpxL4mC5BE/s7L/Rq5
QEeZs3qJ/JEWt3eQ5E5PX47zhw8PSSHVMDcG4dLYKKdDKKarcQlW4HusN1KefAqkct9ztkggIfXW
fYLFrhwFmeaVnjj5VGrsUCR5+j7Vw/Zq4XhB2vq8gdQ3D1L6QZ4ahA3lHW+Ik0AiK2CibA0Qx6/g
ejam7eCweUmF7ENIT6I/Qi4v16j0v+ofx2DKUlbuQJQF11IUbgIon97Dh2PNkTe/DzYkaWR162CQ
RdLZtoburd+9/WnaYfiUohE8xhANnCz3Y1Ku6O3jTAQnY4CtXCoxqQFxWYIB1pbg2IyZHUAqPcrV
rBrUn313kuKk1BaTmVtu6d9aIgbsu5CmInR1MtlZPeQ+92SKkoM6VmVGr5+jNrT3fL4esw/CpSLl
3BhPJ79oLrwtWeSZ9tOS5eDQ1D3vzuuby81f+D51Znxjl6A8+hV4uDMj5IPIpp0Gh5Z/Y1a+RfCT
5rzrrYKgtflEy01AVusdg4h15EBMB/2Mcl3nLr22RyLGZaAM0bjtE5gl2CI375CwFnxAdT5XxUCv
g8BR3zPv5IGPEuXMDGPWswNmtOUdMZ54WuC3kxSTfZw/AYm6RBXdSEpJu6dEe9uUAOyYyOvMoS8h
qDu7VxYrdnHufNHOEKO9QRUIcdpu/26vjPEiLdQramHVZv1bmjHg4wxzAV75VxIHq4zqDdJakO2I
K51yt/bcRH3/F2BkYFZpbDtW7MEfgglAL734MdiB1A0J9Byf7ikj8eLJA8WhOE3kz/Sj7525JpYN
1j7fbOvRgiSy13RtRu0ugRqtV/b0jEd+DwknI2dSmxmi6gAS62Kr7YjL/tdHebBusGhwdvTo08Yg
bG99Lo5CYXJYCW+DX1m/YzIlwAjWcB8B9rlsKKIPTXuJqEM5cOql8iRDkcSM0hhtHLK9BH0qerzW
uMDzINdnbNLonIS7GEuOrpiGtWvYQ3NKwviWIVPG8o9YWtcuShEkMCpqxb+WuKLW/vkMHVKw8+Ik
dgdqRe7NS3ZTO+PD84uMb7p9ImwJZBmiiC3GkhIk/a8RIIJFK5woetDqKjzdGOVOiKl4RyGXSRIj
7qM2Nk/CFA6pjEZFOisZpJim/HbSc43mX+XoQCmM1eFpzNqU89dbGp3a8PxNjKGCUUNB1R0ltWww
mo9e75IqjqBcc1LZnuYE4hSr0WF4tzXk+MVVb6h2kH4wuvZLC72kJ3h4KMt+an9d/z95MfaWfUDY
6O9vXfEc/WN8J7t8KmuSNWkuufbho5zc81YR0oolLWN2ONQHgmAGGMN1WIX61Lvgkehl10zG990f
orRyesb8KgNm8f+QJf32Dn2A1PuZ6vf3SE7GiZqlcreiGbmAmT+KQAW1cP9CKawX7St8900zU/DK
6KzBWLqXLbQSxHF8EYFzdWxGncnwo7mxBUloJWh9Td875DxH4OaqKbeauPsE8aUxTcvJpBv7VCme
yfu6ATH2fo2OwR//LRQ3E18KA6gnFl7CxVjJulpUmNrmqB7QQNo8HSX+bqn/fP1uF1KN4Zag/VEp
OMFjg1cdCNv4MTM7QPIElrkK37fheBB+n+7cBtpoUJvwKPFpOoN5EKRmyvGqv2JZXteZudKV2oLq
LHFaWkhwUd1stMLC4O2bu7tEiiFSE7Dl+Df4aF8y+NyXQY9ZtQYq2QAlupouW2jNSzZ656bZQKka
uPieRRWC8R1bJ+V6zMbUg1VUKxLvfavvNC+kyuoUsjSppNccGYqjNBJEX7VHSSaSc0WzSeCUcFGx
Uq+W6KBCKsw6e1dMGa+TSarWgxVwLEkSRHguPI29ig64cJpccVcUiFdKrkf32D1AShhQQePtfp1c
H4LKpiYSpnXAjpvjJX/W5DGsarpxVLwA13yVcPI1jK2Z+Y5k3f8rBb8jL3h8o+pAbt2IuqfYeKa6
4OBgRsqJiQHZfpOk5WjIhKg+Rel+SiZFgz+7+hxTm4NOTzLRoOZ9eA3zpZog99p3H95QZIjjOt+I
AO0M+X2ESZzONV2STEKdqzhGaBefRqGBvIlWiugYS7tXSSqbCTMAtrVICoGbZILnvTRzyqyI33mC
B1egRHwN9R6dkzDGDsZq650hbRRZ40RBD5HK+4aO1Rdi0NhIK5oNqC1Ax7MSFrVQZ7DEBaBkzllv
XBUC5Ez2FQGIn1FNJbhiuc9ZtfjuX5WG2hSnZ52AeRkxT4OxPm0JvTE78xGyOEQ5XU5Y3VTzTsRN
7nrnan0wQUMgYK/hQcK1QitdFvjvhaUGEdYTg57O30d+VBVyBz2TVaOXoXSHMNuuyHmtY5C8KWFm
LVM/aXUAGaIhhnDnHR2aY5VmP9ZXJhmiU8cs3qZslr7lsymT/EMpqoefM7zODEUPsYEM4pqwol6L
QsnREMvVrD9S9x2AYqu1P5LlgYtkE3RBkn5YZh9qj/ElHTc+14ngmpS8ii4qNL04BmbhL/PNJabL
kz1DBLoJ9pjBcaat7aGxG16TL+8VUtyMt80lziyNXSQhPfp0jiwkgJMihwu113vE36F04njOf7Hx
n6LLYkwJCbNAbrxW54qOW2ooqGWyJTWYLUdWnE1iSw82Lmai9xHDAfQJDpq2aSOuDcIobin0420I
RIti10i11uwsVv+/zsjqlwYQJOs5ivzMcvaP9g5CeX7NH0m0jDTYGYjGwYtqI2PSxSlJBXvHBYbI
dI6YP+qubS/uRJlo5QGKTJgA2RUbTiBEXdPykCtcyYNE8w58nli70y3qCXRqT3LolHmIUsVgkOGY
JD9ojuaIsXb8BjVm16diwqGXsmA3PM98l7etl8EUXyuh9iRUH28Njl/XMiMula4K4k2GpcqvoEbx
zBHvaFqsW751mjiK9DHW8thHVLEJA4K2OL2X8uZcQ9dxj0PB3G6/99K0Hd4rX0Z5jNIA219QlA+p
czuGqriAipmrTd23tcZJVmjpsuh2X7w0EDqF5IMo5VfrEITwIqC/5YVxSSfz7PRpI7ljVruXXfE8
q146reZusYLzlXC13wrH49wdOPveIy37oTL1nWa9jQYRXcec4QZG1QrMkaUb9BxiSKcADwTHxhTo
q9s4ysoooMqeFG0ZN1AZV/RCwff5RuomjsxJhfURVIA7qTRyV+5UYPkCakVZQR3PCQbAbWIKgZAU
BdcgabrFlUsaLdBfBn3OMr77uarjL6HWzaCMgX98XPTEv5dqR5HOsfqwsLEdhMnmrr9R+frWVUkO
KvulUlfQE7b0MDlQlBGnDvOPYYkktVktXxXJkQS/WG/U3Ly+DpoJ4gjijW8qQqC8pUjHmBlCHBIK
s3lEFzRON3N/6NMDC5KzlbKEeq2SOmAnc+NzRLyW8f6Umi6R1nxjlihMzZOH0inzv6yeW2MItfIn
6eCTd/23QM2rBvCwuDvOJZFhR1bgk+Go6TAmCRTtEK9AxoFkAOEs4wkCXC2OqG6a7mfx4nBcvM3m
7PhLuK0ah9O3+GEMAomC9mE033Hft/OzNQixRkis2eIqd9y9lJ/kMcHjL+OwrW7rEPjH6OcMVa6n
qBFfT+I5t1tvHapaNnwrLfcw3i0iiqYqXICHC5nyEWcC56S2byR6PPCfeSBkDInLtP5lwwVeqOwH
20FM0D8245uNlbGOONfYUE0HkYS83OoMR7UHvVn3yS5MhjablQ55x3aU1e7Wgk2ygdh1Aq+iUHt+
HKAhzq4lyWw7D8AGuOUoVYg6iZa/yEf0g1w+HYDKPgVfMHMluClJN6uohugbDICNuSRQAaK33S2o
ZFjwdfhTfSD9COZi5AEn/lTp4hyuzR5VzBco/w//pjOVKXdhP2d2LehP2aAlm46r2EEmiq2P972z
kCk70kvidE4O9DNSvZazZX6xgRuyi/4FfvLCpAYmLLeHryDSxuIABgNzY5Sv9K3fIwPQVXVGI64x
17puGy3h9/2uu/ukHO6k2awX1t+jUV/Acw8dDlXmtt1O/TdE5Yoin9NIom6HgXuxBO5mByYHAj40
e4a1yupjDY8YSnCSC/UX/ZkN8TPRNGOUuEMUZfIGf3xlAf0TCcQqq/qGWi2vzAfMe3/+t+HZCm1+
51IloZ+xuR7vQELIUQrsxs7cS4f1gdKSgoEfaqEpp8I60UBVX7OiXjg242BF40IbQD93yukyHjlV
GA3ONmee5lCadJKIBYsYZ/cKIqXLAY4s46zRZk8X9w62r/UtBAUsiMjIKtlZl//dgu+ocZiLG7Su
2LHgcQBgFpR7/KntsfQpbKMb1Yj409TpDDZxFJ0wDZeueMgQAiPeQTaxvzgkRa4NAXDmhNcTON8m
1/cq4UkDgEGxXR7SGoxhXszt02zGdYvM5z0YsNmsHS92PMeBbHtpJwPf/vTkQdCyUzC9kthKNzNa
lJvxN23xkMQAWTtvagrID0YZ4Hqk9Niu7+/SEJHXoys12g07re5JpvmBwVTUdvGuk0rg3hYN2K0H
OeX7IVsSbiLA1zcbzmXNH0C6wMgR7EPcyc2Ox8AdpuuGqYxmRqqihfG5G6Lx5j5tWwxArPPN1SDU
HTUlnN2RsKX/IXxMbGgIHIxOiVcI02a6O6MG+zFcGXs11Zsh6R1q4DarWGk+IzZa2quPOXcAZqC7
uPpe7/rBfc4i+5rhOwpK9+K3MCUk9K3M1XvtWyz8FbzeuHr2vTkNCuay9olpkJHpaKP6UNuUCYDf
e7y52CnzN89+98k+USx8TtCVzaWaekcQQ/irL6YNj9dlIywI+O9J+C9SEgw5M0C/387zd1oZ5Jyz
/l3T3pJp5+sPiSa75T8Xq8zdZh7/RqCsmm91HxuFXIoxRFEDrpKfsh7CzAdMVvGNr4LTaHLpMWLz
KymrDyzvWls83u/0KK3PNlWYl5dPemh3MsjJKSMJyyWe2hBSlwmRa21va1vLLM9QRDQFLM72Jc6v
CbiIubRjygnJJYQtKSo1AtNWwnPmJqMjv0KMdwILpCGKBblni69jGO+RVYxgWG5HU+P8iLzC4M7s
m47xSS/PBfuccyWTg2zQLt0T/f98Jd/OODVRM1ADjvnVOV/45EXtBbMB5S/uV+TDRzvq65Uxsi94
U/ZpkAy5Bu0NU9OnpBYQJ/7y+9p0fJ5LBdnjCJXj1ewp0tGggrlDQG6xph8bfuAtncCkNQ5uxfuE
7CaByfWGG1xuH7LKpgrPrjFz95Ly/ZWPn/Jp8lt31Zm5oe/SuZ4URpCnkThRZg+D150kKA9fnlCd
8/axKXuvcsOw+KusyzKhC+hPk9xllcY0PPCsaSIlRTrdqHv1rKsdlWLOh8FbxrHZ5jtzqe8DqEaa
dlLWfGG1klhFpbwG7qdSuLrTOmtrbcAi/kdU+h+lhhcmrqYDxux9LBzrY+6IZb0vKz76UXzNdn3c
HnRMzU779L1NcpW+vsJEKROqPfi5P68udgn1KAsuc4FeST+qTNOrNpPYDZEkbmX6e3bSdBJEmfkJ
UtGT10ZvKcalqBDfnT0EW/+blHzkwHD7e1X3XB6cxGX5MStBlhpCJTd/o9VZElf58rG9lRdhIj8d
erzW3f2O9ompHIFIJN+M0TEq5dNs6n/K8DICc06j0XjCA0RAtGHmogvpZ3nWP5lp5o7xqvRl/JV1
zQwlVRIE66iaAXryn0l8OWXoEPiWNiTDi0POApHrVZgs3B7RahVUFo8bg8uQ1ryJ+ZINixgbfgjp
0n8xTIoQh1l1sm5TQn/7RdPLYPg84yPk5Th9uL/oeFfwqj/K2Lwd/Q9uCT70Wfp2YEgltXQD9KXJ
o84tMZGimpvrrsicWi9+cz4q2QV/8xicOtZlS1qy/oTqU/7JIQz1kEaQQAUtQer7++y4zflIqxUu
X/6hym0xNO4wCh8alqK4z8p/AnQtrKXx8PPgkewEF60Wr04UmBjIiDUmTZ7QRWW3E9SHRXBBZKYD
wn0z3cwdR0jW9GNhKRKr82Mbx+nSsKoFfp7NEC9LA8GFWU2l096tlSJUhDGXuE7IcpR4NfCaqYll
z9HRosSw9Op9MJ45h8r4yvsrnnReGLLqanEzNOAOtTi2PE1RAW5N7fT8U4BqlFyIin5XGfl8udRm
etKAci72WEjiPYId8yjGao/mrNXmRn64z7XOK165ix87oT82LG0RWqmd0jCB23z4oY2eox64pNO4
oVyLV84WYaDu6YyFPVNmNSDVHrdQTD36Wes4WD27ryMpDSlDNS09ktqsetwQv8m+FQCt8tFbmokU
afx2F5he0J/E10dTsYjDYwkMXeFDUl398DoRw4+QSdkmXs8SNLY0IlNsqPJFMi4scwaG7wX3g1Zb
ZJvJkDUTfAiFBeMIMJ1S4X2W9mEjXShKCnwtDp8PmZKqOpMTzgkkA15hJeQxo+nMsEDbLGUEU/I3
kS5ag/G8HE4r5rt47wXipqBuea4zU1LC7nZp+0/Ow42TzKW2ETXVF03pxsPxpSAVw6EbSbNsJAm5
mkU61tvfiVvZ4uCUj4tNiptZeNbuD4gkPa4mi7/HfqAaKx4kdztaUYkMR+DV8GtciaocPYlnDKnz
5JkHDrXPB30dE5w+uxagNxylnz/51skH7HjnPwXMdNgb61D8qhknnm7rfkFosB4FrAZqT22WKOW9
ABUa8+R32jg061UV/COe6/DkI/Rr32P2cIESB4jHlXN+se5FKF9MQdAZ3DwTjXWO35aMiVe67NQj
Dakw6VtDJNAOM7gHmCkMUl++Ho+SewaZ31px0lLW0h5eRFVrkQ/sRUYKwZu1tNivfVK4XcP4Y7ek
yF/hU8rfOsMbLzKJs5zhUkHMXwkSn9VStjtBH08w1n3umSKuhgMZWQkE5htMlp+N1NVQf/kTdw4C
yzIYe1f3w2+/54nVga0lV7+70si9gsWkcchfxPfyIoYCITpNdO1CXQIS+x8sOQJYiZAVkXcoHBkL
wRl0D2ScuB0e5vAhxUyM1J6H02i9mC3TzjcG/Q7DXdRmicQveGZTMMHXNBcQ+4rS7l18csY0xkzv
lsGOG6sbwkXjh4ujStHCrUM3xnVHtKodoLUvjF2IeEUFfy/U4pBwyzE4BKGvc2xBBKmYiBKPqs6v
MUqkKLyd/sB9i5Ris7kppiz25s8EBKLeNDhqJQ/n9S3nRAvpP58ehLTS8VH5pE6iesd84tm9gT0+
TZuS7kBr5rIRvovoWhl08HA0MJNcOhcX8xQGyN9o67tB/VlvcXrRGXbCWhl8hsac6ljmkmqSM/br
iS/uQRJWkIw4wUDc3qIKZO0iCukGtWP16Z2VsaWZosE8jATYcFr1jUDG4gx1Cra8lDZf2XAlfJR/
j7ahQ7YcWJoyiMLrNsRJI5LOjlJbNF4dAvFHaMXgtZFVOpN+uQuAiPqUJyf7D2cE+FApRsqJZxtU
HiO654VLepMV8bkb1SSyyej0dSJqp2TKf1g8a7dfkkNwClyr/Yzez8uMMPe7qCqQVGVybtJxLnyR
+uWAJtESlBwUVt2MRgi8wvFBjFuxnc5YbC9GKUk4id6iX8wiWd2h8Q47VS6S6jVJWj3yoaGw+vr+
OUkBblbdho8rpERxBZeNNvVrmVzxnnkSUwKPJie2t+4MsNT5z9erWvgqM5qUpoOEq4j7oOPDmkc4
OfrUgWROtAKrM/alhVfWCLuYhHDZHFGGyont7rgfk90kj7J0P7JH/0uOxwe7iqUlCTh19aHCYBls
Qhzu11K5EMvCF8WH4uFH7J3/+elI34/qy6HwcRPAGMf9i28UaLZo4BD2XWgh+a8PPHAw7A9qOctv
m1UlgHXHRweC6Atk7Nk/VZUOZxicCM3n+r+9PM3oA+JAPKK2RiyY8Cgtzrry588MQHLpKkMwCtNK
8KmK2KEqx396/8wTb4fLgocGNvOsqbghDeUdlWaPi7xn0pkgt7mIaz4BtbVmWpUcu0Lg8MOgMibi
pwiXIX7g6cP5Vw9BO+Mt+z8uxQY3F80NftqWG/JtH59syvUFNfTCIU2oHdGYXmyNyuPGyWNXsI3q
vMx3oY2TK1UI52rjeBeIYWNaL5o6yWRINCCjUY5+RBQqmcoTKGiufDbYAzN9on7pKqaXS0TKJiTm
6CF1yDWDa1yvsK97qKnzqAXNFYR4xvVEHtSRpBTtWMcN1j9EZBjwb5IYuWENEQwpSWL83h+buBw0
TmNg8fUaz2t0mToUr65mzkrUNOclLmLJBQoMibYU+CsU78/kapIvpD1QKtf6ctHqwO9C+xXsQlQH
3j/xogI7xq4qptmiKjqGOD9e02DTKHBGCaJUWUpXgRKmF0pVpfYHyMgIM8GCQDQrGMyN8LgDwqTu
E2rUsFGB6h/M5XCr+xzuSHj8lEDFqsXlds7rgrJHSsOHbufp6s/UkQWxqp/RxWOgsICohQo0CS+4
Mi3CyrzbaRMdYouXaUElktpTsEnAYseyrUTFpaAfIIG0zzA/a2+m68feOCD/H3lKIJRQeJWuG6lT
N147shMpH3jAls4pp+KCntSSSWbn90vsT0W2ij5d2g3oEK0IRAPh4HV8TxTt3Pm7LLCl//GarP82
CryIxVhMZ5y2zDDI6ybbgclprfeybhsxj3pWKdaPzg6puGFZ8IuhxXpXPOHsqbwFoC3pGNm87gjw
/wMgW/IktRIfmBRkMGh2jzgVczi+ygqIeCsd1A90wKV6VrxFNEZk8QEGo0iAN/dX1GVAdvrOyViy
j/YS8lwzvymoIJ3ok1HN7+4bh7ZcFZkFU2HusDnsDViIS4NBCbctuaKRMItHcelQYw1poXfu6mKA
VUWDpsW+l0KkVovVu9wM746fASMtXe0nHHzeaSTkG8rc1dGoAsCwIuXkf1nxpcE+PuA05i3yD6Vb
FjnkfK4tuFQBmtwyGzVlWbmH8/nix6OYvuBOBmv9JCYqwD/TQ7LLCBbrhcCxlhSSYxcVaBDSTBqW
5AS9Rp7atv0CQTLGz+gEUNaNWoQupAtdIK+QeWVku84joXs6oTY/MqJUbWpQcNyPj1jq1Za1QQpO
4GUmtD0wBZ2Usy7Z147rYZorqDLZBGMEW4bEFrTL/2e445IE6ShnKbbUhV0vMTsucbNCOCmDv6+H
zXzMgiTPC0u0bmes1P9E8hW58X8Dr0Ynd2Wg2QrwQZ+jN6b34ZIu+EbuFgAIwAYXLZhnwroz9KL4
RQvpGUUkDTf0KZfeNdv9e4PwT4xz8kLAheeuuvHWDEuoNL6IIC53DOWIUFxw5QocPmKpqWpR8+rW
0ajTOpwDUeQuLpGAMIdPq5aZPUIOSwbgw3wGJ2k88zThMPWZ21NjRJW+l+j8ikX3O4NNI0wrTKNn
6C/Q6pba0FzcolwyePCR9YwoW++cLXj2ZxV5313fHQDtcd5Nh2bc0xq4Olkh8RlXGJLOOcZyXYW4
fKmPnZLuFr5vyuHVav2EOm9OAn7etkWpOvIp9dRMgnUlZLUSx3fZEbM2Nbpwpc8PsB/untNfSo+g
h5bFTGks6OHzmDTQIuul3O6VYSWaZsiG0PzCTGveMMpnV8Bo/8R2+fVo2J4tS3FVH86tYJuOjazO
j9U03Y5cUAzS69If2v/nfzPL8y4h8GDgSpeGvmW9ar8eMvkzHqdlm9VlJJizRSPlWIrXK4QNjv6X
CGkDNDXAnYGv1+/7ziDwwLIhnqpjNjl7opuIOItq9egjeK+6rm4T83Eiu6R75UpTqf3VKIpefGVm
JlHmAuCnf1ebrf5c/uhFlsSEbv+4V4J0pPy8z3vPlX5sHCDe6u6WFtZxb/3dtlF1A6fBWxBp3qIW
LZgkJh+TXC583JR+iWc6vSzJr7rdIPK7orETtqwlltnBQphSmHRruan8vS7yKHNPy9uUBHjx9Rn+
poX07TUiB1zfZnXgA4noeZ2nnMaktQNZn9Cve7fAWAXvPjwtCrYxXPaPrlypiR86Cz9dt4BJDC7l
De9QPq0i96C6mX/dtLULtqPwc12uLTAi2cC2Fxc2dOchjakYIR4ghxDQ5oHMN+nI1C06u6j2oryD
rL6noKxWK2Ae8IBDu4y+ZVbLvvUcVPEBWMMdAI90i+MIoOrGuG8+qdg1YGeSfK6l+lD+yfGX4z8k
wf+AtninQncKgxdN6lxT/iM1vRqdYnOlnzGUeluZ2kN0va2/3RTMVC8QKaDny/xC0xQpB6i8fUz0
VVKAudJ+SSUEycM5vsDGck93MgplZZDn4+w8+oWNZqiaGfhY1+0K5JSxuCBVEJOE5pY+ZkGf6Dai
glnR8K+/0mkID9DiYTG3yz2rioPMfAzowJM/vqX4GQzOZj3IJhw+I5XgqDXBM2w2lXRXBi2g7Pb9
lEyJpT+nC9A2wAAVwemsoFQENjKiJfrCwg9CWd/MfQgZm/6DNB5MCfGNw0/R50XgUmvvqvpS+qtP
MnbJKCKsIymNsj7a4NYbc4Y+JYjzy5PuYpcaLQY0OlMJcQYZFyhhy/eowzAb4sq0pXJBbx9FZPSi
UBU7+utuVg5dhz6WpHaC+0ZKrIG3pRpwq93oE4u89sttxt9Ul+od9vUHHlj3LKi0nE6Rq6qG9mCj
Yzdd4lg8PPU28pxWBhqbvmudtw5wRPKkjgYHDLyPGwuP/FDjPj8IXfpfUlAZWuujFKetDKkRdIdd
hnRUuxvY9hwNxqRgFapeLc2JtNqcNvKJjQELnWSwkpLfaB1X2SWIEZg7EAXOChGqQAOLfhvCNxhC
ZhaExUIG9u9okzrSrt0vwQxGkQErsgRUosr7tUxnZ1BG79hXIMGWOXY3+lf8NcbMXxzbB/4NJOmG
d6vTN7m493/KSr5yE/pNg/ghCF/mQ9WDdUH6Q/AdNlKhRqhBs4yqgORx1Xo22yKYtHc1x+iqqYW+
SmMElUJJQwt47HaA9XKY0QDJFGHXVdPkJen6gijFkfomc+dakCjTO5gVra5qce3/B1n7kkw5EnnB
XG/+VEU7IkjHkO7bkx/TkOxJqzXJ7lVOa8dvABkeO+egQX//ASjVz3R9qk7i4NcCtOZ42K+fuAyV
bb0RRnJa5fICxO1CAGxDVB5pSx2rvSLwDi9hzBcTHVQjYD//q41F1DruruyRcOaQWFUjp7bD3pyc
Z2jPzkIgBMkmQiKOCSXXiBAqeQrQb+eFFeiPi4sZGNndm4y5AtNM1vHKjQLSMx7wSuTwAbuQX/0v
XrRn7tKQ/Lih1LgWPCwJU0VcXHx085/JcUVewTmclLCdgCRi7DenFzpdHpSUS7WMxJ0rLj14zrxy
iG8PfNoSVs5G7eW8JEpvvxuMWIX6FJ6dbpmBwtmYJwmVRgK/Dr0jy2SOCVziNHomhjdEzZ/ok+ia
svmNl1nsqZXFom4WV8P10SMqF7ebh85oXdvZT4lquxwyclER+IDBy1ungayB/LyD+3VVEskYj5zO
EMTxwoMJBpT4zloPM3NB/j12bTaA2ZK5nQJXREn6JdyTX3lqYlzaOvafTX1vmG2TOSPkjEGzSEb8
ZtREHnzrlRjFURmuyByXay7wAjNmwYuKn0UBqnlEA7Fzm1uCI9Bb06p+BLuDD8t9x1iHewow6WYw
iAZfdaZuXi/uMru0cOpwb2r2WNKIU9qsFVGPVL30ztf6eCpa/EjzXT+vVooYGzqJJl7bIKu09W2H
FVSFlMHZYv4AouWKfTBJTdC9N1JlhksOllaHI+cRV4eXPfA+CeoyG4qVjovMAdAz80y75uqy6L7l
IT5Y7T7KkFHmjhZ3cm2A7/sZn7mnqniGThrhRHMxb0Yo/0UCteZcr9hOKQGG9wUoIpWaxj+JA66/
JIMtFoOq0SIqJA2FBTB1S0TLC8GJcxRvay+kL5Fer/bouyxgYRuzlDvLchq6LVcYQFzVlDVH/Rfy
mRFSIydCfpKr/pnyRYOJ8+Rg65Nr0iwkoMS7ZEwR+E8LbiES2l/tJAYzV88dANXh497SEnGBiWmc
qBoFL5HHnexHhJ5uhvYKqnIohoed817ICht/6+s0aCmN4ilP18txTU3SrpGnAXYOh2V/WXnER9jj
YoiUfTc2IY74vTRYOvUij+WSfc0yKHKHRetCZPvkoHqF0q6GqmiLb6MrfDhTU26SJW7cuXSXTDC3
qIu4kGt5u7IQKgXGIc8Tg4yH+aZopEFpChuhElcXcL2varGNdO9xD+iQV5j0WROiMhrl7TnzeCXN
QRAM5imxaAAmWoh0tKl+2kKljx8gHO1PMk+aAvzhizUm/nyjf4vvth4rcqkFZCDd7elP5mBkHfQp
NOMCsdFblcM2X+a7iuEbuj7lkeY8t2E+emnPivi0P8dtlqzkLLM7km4D/v5+Lx5t0bBiDoT5DgOC
sMhh7jeV/hW/qsPD0xeF8JNRcvMl2kuLbadT2jkWySegtG0IaN6Xe2JulLqlISseDggRpSMqV4tx
HcTLtLrbs5dsjgSozCFKlI2RNBMd1O9wgtSUdD++v00N29mVv6VOkaSjugMD95GViUDmZJKSWj8P
f3u/rK7IhSEkcLvscMXstEpXUoCrwT4EwlXJf7RbSiycjxuHlThkpeUJUshg5MQZXIrr2Zyp5n7K
Nbxe/hhujAISrFWX+8rmEWAljV1qPnQ53C3xDPU/oDSlnVBC5bXsUWCoqbqWKx9NnwpL7vh93Nbj
OkpuniWecGC0UhEY8WwHWwgm5ad6aFv6mhd5/wANN0FX4z7BJVAI8QvoM5rnljm9x+sUAA1gpxzf
7mwWmOjdk7+l+Ag58va262dgoTlW2q14J3eaZ4+RfwqqtlmkgprQH+s/A9pfGmT2LLbLpNhQBD27
Gk/fs1c6sts1RW0IuPzBXQUOZlSx7iFCZu8q3AVb8UGRcpllCscLbIBia/cIcKypr0nUC7D1xkZN
hPzpbb4ewVe6mzHt+fNWtVOYWnawAf1MB8ZD0DncjwI0uH3O7mN8oAHBz8hd72kyK079SAnHZVTu
eshr+HNYSMLYCS1TP93FWDxhrP0oE4+ilqr36+Umnn/yNgcLyJntXwewohzvMzZQs7hucuazAJ9d
ZTJASSFm3eakZ+GKhWXsHlMmijymvChkqfI8QzOS1VWdqGJHBgCdjdXFFzZ2tESrnJdaKsF/T04A
NOVridCc0z18U3HcxdXTy7uBvgnnuNO4GtAMqX8+AUhK/BDYBc90a5t4OZsYzAZcqPfnSQfftoy7
blhXLtU3sM6+8yBGPbEXtW/TK1mAK9DXOKflOVcGX0j8ZIlat6cM81bWrOJAbIR58DG8G32pGRgj
IcIqryDH0L4bwKrTM7q/w8XBtMeEe+rSl4qlG6fPXJ2hNuw2fdlFFOSmBGHcL+G8d76fLtcAUKTm
m59EE+0KPxT0uIDwIihembdCYsvinc0sEqrXSHnXEOJ+qZrNgLd8RLoLrhuQYHj2HrZ7Q409MAXj
nkCNvrZO8InMjLEoMIg81HUfAu/IZP1nUP5kgTpfPRPxuOhw/p9FY2HHQTvQVvIdHnHXOjB9/5w7
qcBNm2s6FHwc4Dyh7BW5SCnPH/cU1mC4vAwPA+iJlUKwkbHNrSCslE/z5o8LtNW5pGcSXyTRfzll
Jrnb/RBp0U7loXLc7xTY1D1z9eOiuN1iGmi6I44/I6QoMFaIPHe76juxZq5jlVArtcrDkG/pu8SX
UYjVvbmjWRzf1o+YAGHzLzJlbmfMi65hhV4kbEq5w5upd/Y5fquION54eo9VKDi5aYAdWpfhXVbp
mJPff6AkBvTybED7XwUlc7rn7MI6VjX3/NJpIhL4f9/4Ka2E36m2yDueCW4lZfjuKTGl+AK+N/3S
hqBo4lRlsirZM7/Rb+MRuES/HsrdSppB8K8poHBB8njDbCiNZtg8b6G6UxHcSBg4VGUOoQCbiz1t
UlEkbTmROa0AqdboF7xzhOYMZ6lzmKe9u/9K283guJO+b2eSEbxSKgH3li3hJpfxcJyelSDM3qnG
MVOOn0StDKupUKsQsm0RMRky5LosuJDTJxCJMR/0wgzFtOWKHpcEhFdWj09pOskTQBTvzDBnqUAY
cbjT2L/AwvZwJKkBmv2iu3kED3IsI092lb2pQXLohM7xuT7YQ5QZihhlGTdFZn0bfZYMqLWCeRiS
TU66EN8rQBm5ntuhK0OE9+bd5c4h0vknjLpu0+44vNTOGQphQ6H11A63ycMQgYPeq4vENN3YKDWt
eGwDGcitYnXWXofKcUwJ78ZJ01Lbiu6Tvv3LIL+XV1okqGK5G7co21lo7R+P3CQhvRiVpNTMIRUg
xSSy24f/joyXIeVgoDcmYLkPdiblDZMGtjY2MGjuRfBQ5vMGnM9R67jBfGVLf86/YfhPAnPWOvEl
icY+lN7aZd6fUuHRRWPUO9mkvZsTZyY2HH7oBMg+xr3hj3ul3TSirjD8JHlYFTyDQO+jZ7KGgddn
MNz4anAMmG+T1JIIjLwLzPOz9PDvxVkoOr2WyZVQPMTUMnTvD0P05Vu83CqJZ8z+jz650lgFWlWJ
PJG6f/sIeJ3jJ5L4H2JZkNOn/hnggFYisSwS5KsOaQeUf2tIY9yfaPJDLQe5m/RzDvK9XPin7wHI
4espVQDS7MhFCfRCyUrco6kPs/trPfNZXM7LJVG39/FFd4LgP948veaNMhNAM+9F5yn0JS5eqeo4
YscZrOQMrIn5xIV9kjUnPsWiGuZXWL8pDwrR+GdQcQq//+r/8PWCS8isFUjt2mHMgh2WFXmwdYsD
tEvxR8/aTbAaj5drSRa0S7pJUjwL+25MYL35VxRdf+MGrHnXJVVl5KaCJTpq8yLLLeQ8BMtj27gm
oTp2E1riZgUoZYSmy6/RduRRlkEpDBTbngcuqNt4EjheGVUmktVQ0WcgD9NwqcEB51YQIhM+cfTR
vvW1PN/x6RVTPB5nrh3YZswfvnid3xaDur5pOifvVZX48CCBaLiztIU3Q50kkeJWlAqo6Pcj7ZMB
WAaAkOxrAZa4VcqZJdG8XRE9nR3OM9FwwH49sPs547/Xa2wXm39FtK/Kk9Ypz2demY3XFD/whS7F
PbwEGSwiWiD+bSmsgs1I5qrFTwWhxF6Hb37qFwvDZtkOnYB5TKQYknyk2sXP6hw6/mOJFb+bGWCw
d62eR21KNS4gXY1dUzdITzO4mWuj9soKFaDA4H2Z9QKgBIvJOf2d9i7dfC6yBnG8+Rz05s4MU5Z0
1Sgw2+j6BJ0THr9mLOmRQSYTfNx9Dohm9UY2Khg9QIHkMMFPea0RnKABzx5PQd1eaUmMaIWCJAp7
xql6v90bzwJITVDYEXOtU+vQr+u9iFxEauH+gP5dyYG0+7CqcH3EyhXSTeDP4+NvQCbFsITzJ6vK
EmKTAanbeJyAfGQ0rv8GVT4UNffergSD/jblM6/KoobQRjx0YV34So0fMPlFzHnWVzSindoxnWUO
rbkUD5Il/VimCZuSkAbxXvoxQTogB5dtdPtzxI6qvmtSo4OXQQMDMlnr2Azfiq36K7i6TDNluUfh
BkFr88e/7CxhwTjr3YoveW8JDTO/PeR51kij+I0xf6xCpyMDov8yaf/UQ7R71e9GKKhaQIiIg0oG
JWRTzMQyPlCk4j79IlLfww1bFJmkujxHIgNM1lFXRJnU+EgEow9K/stYZuBhOUyIVt9YXyss6mNa
iW9t7wous0yyRQkjM2PwgvRbZOqKuLmN+G28U8fKHPcabRjucN9mW6McAH3xVSe2GqS+60xrjYr4
lWisj8HpMaL33qfOj1PsyNpUGQjQ9AQuMZm+FtvGAA+iqPoHQeoHojL0AIGUTzD7heFyRLzvQ/Ai
or1PC8vEh5EfjEDlbP7VLRxWJ2YDtADK2u3o5yza7TCjO88SjDkLLNmrZ9LaY11sAb5Czi8bTHDt
ALA7wbxT9B4/sobgZCydFf2BU7AyW7JaK0kaHqRZWqXArvIEq345MnKnzrFmTFDgn1jEE7k90kGK
JmjTPt9EaEwBydW7tj+ZI64s3kWE7gQAH6rI/thdlmfyMj9qS4dkczTj2+n4faaXLmbjNTOHNU9Y
v051GcTHcCL9P/E09FAzU9s+M159GYIcMHpTWLElKHHMPEVsr7a1+nTcFgP1d9pRVP79LhdXcY2u
xB7XbE7MWUhUMrXOGGWXgU4+y7ZT5KKWNudXkrg/qmjMu9tZcL8naZUsOVR4H7/S9QRnLx83alRD
2texfoDC/tktPdE7u9vUdQTAFGiYYbRX0lFu5rpX/gPNgeGrxpmkBaIlg3RoyyhEz32bFCRQC/Ku
qHAEBDDmFksN8rpPTID9qQy0eZnhOd+zCDiRfGkpaPzofEn/j7b9UkrOU+eFC3APeijF6Zye0Kl6
FvqtBdFZEgEt4KFz19FTCokaJdHZl0dPwOveukRQg7Z/P1iwM9+Fv6ADTxDBc2w2IaLzZIe+3iJY
z6kT9uATBp9diPltT0h8vRl2ahgXh41n0b9sXP3TjH0zbK9RqJgi/Gy6Af4TKTTsLgYvRXNOJYeK
05TDWBh5nI4eu8/6xcFAWpYx9m+d6LpaTKtv7bmUyIyNE7lWXb6htFCgIH2tcukn+RFLFSP+Fxsh
p7Qh53wPEzGxtthAFy7+SQ1JKQGcU1URN5XXRiRYCIURtdajRvuHLyymx1z/eiPAe/JUSjOW/CAw
YzT6kw5e0BRE5SA08QbKTcI7PenBtnSsQODoyBtvSlfnz7iy/dQ2GZdU9192zJOdl8NN/Uu64/Af
eMb8QYdvU8Pcgi+YcZKF5FFsK8nveCJ4Fz8HzsVKQQ/mmv/eQhIIfCwzTIUmWGPB/6orURJuP40M
wX7C8OdjreqvuzTwcGeoKFpNOl39HEsRHqN2gd6/q0a9pU+qfuxhBGgPdLc9vT5olYrqq88f6kNS
Fic1jYiij6sbw6j2gTh/E0xo3xS1F+JfVZcOUt6aTiVBV3MyGsRkHswXHxavBi1PsCIEHhFyfwTf
tCHBZwK/2RfWtSosRPBq2Cwb9FdW82w3j/oxtAvtfG9kRsdgyM0giDsmXcJjr1tkFKro+2mes+pl
KO/95tYfVFgDJRbTj9ksnuTLnE1N1EYO6D+SXjMqDsL1d4dfVYZMBvGm2uRxmzsYSJZ5H5cIvQUs
KJF6jDpYOwXTvt1wC57n7/cHplnvpPXZVi8MGnGRIyRn7Dy2ESdBPuRh6NC5tsla0Du739Mk+z9v
tP9wKpHDnn6uo6Q9lXfsekpqS/j0nWjNcn9AZH3OhtsXDTE97zhofEfKFmB9SjiY2cxx/qNMJBa8
zlLtsiJ0YBuflpZFktHPWo0erZIBqptxwBtpmD2tIjuaa1/7m/WpFTpTBoR8jE3YaWi5NCWsZndI
o/w1y5hEh+zhpYQxc+59e7FCt8r299XOOgxHHfdjLPE1pLs2E6S93ezJc1dZkd1VaDZn/L25F40J
Fjm+EmF/zP0Lcue0qUtPZoUme/3vKbUtHWJrXvVs5AAy/f81TXxr2jQ+sb5dZjAjSi8nVD6z2Aze
UyBe79vTBDpIYllW2VYm8nB/FdXVS6E5rlSZzWJYfK+flkvWbiJp64lQjGnVk1Raqa2CwOhMYcX2
/8rYzCFGj+V9vu2n71umSkoogcm6gGuPSCnSmfcGvkguuVGORpMHSc4FD2JbCWu3ybkncfetESYR
PUJv5ZRP3n3bgIqdylHaB78LZw0dGWuI4kN8pSUEbH4RHQyDFfjvDpekTJ+Q/zNFs4gGANfKM13N
p7AOgS88S3DXJrFZdhamzArYhh8vuynFG/F3kbcIeHKXHP5QOqk34Wx7e2+G/v0A14U7cHJe/2ep
4L7zi149i9b12nuFhqX/euYH32UCG+X67Epvtk948dsz5F+UXGpo0As83DL+ArZlOJaQaeaLf7DW
QA5Mk8LESEOsPUCrGkZf/L2orEnIv/BY+lt/GXgoGea+N5/iePYsl8Udr02n4y5PAzZPf1Ns5AZz
ClcOeJY82J4Ad/Rs1gk9ruu+nLu7+7t7NGrXbt7r1PqBqzgRXxmx5wSl/7HQDc5BJnpPqn15Xlwj
njJtLmnadsdy1R29LpLsLnWWl9fk7uriHao7U1EqpjAMyF6EtwW+lcsQyfs1hV0jLkDqBgcdi4Iy
DBbG8A6v4D71VtyhLs8haVjpFs7T5F9oSyzf8SO9dED4cTicVEPxImrzTegLZshoJKZG1PQmcCEq
Yoqe9L84hcOoVER5BvZgYoL7UoZUn4TBb+ccFxLHwxKcoY2HaeaPRXSqSgSUyKYq5xWpMWmJC/3X
wZHR973hr6v+sTFax9QewIh/J1GA7qt0S77u349HBg0pzVQ3AgUIzOpDWzUZ7KElO2AGhYEkmuHb
KVNjYqjzcMXGzL6Kra2OQ5RmCiCglhcIFbFuL5DagLyE4B9duSYTCoLOMzTP4Ykfpl6bU+GxLI/R
lIzhW3RUMk1HJLiHM/+c3JHNhiTmiZTAYUhNNgqSXOJgza7fGpKDr3wIzGWwP6CikDf/53Wh+LzX
T3+/TO4KYi/yomAOmwmoEP4AarYKq1qLhErAH3q6f4aKcZi3q9PKrDoGBsEOgzLi07He28pbVOUe
FKWJfzKOK+ntzxrFpCfXAktR6fmYrCc35fG9by3ztmzTCjEFIGaG22Ls7gUEzJnmUxwWykd9Mb4o
fxme6XMua4S+fHYlncKXCJvx4bRxLx3X29hl2DgourQLJaKpRbORSn+hoahiLuYVsP2qVAm8veTr
4+NK6KAWBYDoaPjC/lmkdOvzeIDivgBH7oiVAX6xOi/2zvvw7xDwGN7CX+46ymbGe4BsJ2JoYCHU
ePuTKFuoP9HirJRmq0mZauuPIhYjF0b6XugYtYnysvx8gdX0FJKtD53Sr9lraDe2E0wJmyj0SMqX
AWI1WOG0Vl9QQyWD10HPprrEkbVUYsNipPjr1J+qW2qCt9pxze2o0NClHBO3CBJERf6etu35ZwoA
DFu7WvzJatTsQ7Wmhm76RrVCSVrbQeBTZdnW9dP/U/zVCQrpM384UbNKUt/FpX7xbAcHUnLaOWoM
6wKfHNN4Y1onY3qWtJGN2hgtRMos5MSczqdngzOSJ6DSCaAK21x1353d+v3qDfoIglfRzDBJAqyr
vN5wuGd+NaKdzn0JbY+qhGg5XLekhJOpnnsbEuS5Ez/qLPAfIKoeEi7Zi4wWuWO16WpjOBBkdvxd
V4vMMuGhO9RClSp++kx4u4JQ3hNC1tZFMFHAw64PVJo6inV3DC0/+LmLDZtZtG8scP8LKmmw1wU/
/oE4J2jPewU5OfoUXvhR2SwNrfMvLFrUU+9GsAgTwxEkmjlZqhHR3WeKElypQbsAEV2iAyve3xoB
J2BMzCeCQJ5m5Iud4ZUf3HGiKqDpxbT7KdUFfPLXX4ZPVp6nPhdkYnlCsHwsVMT4vNvUpeD4SJJJ
knKf8hdAOeLQMWtcmGxYMA8jAByfvTqGxN7R5k7WDbRNaEdyz5A1pn6rYdpRb6B93YL7pMNiQ7NM
6ouCTDtK4I/bcHGy82Q8YIAJ47eNVN/aKaa5sehvWo8td9kIfkAVb4CZKHL7b9vyxLmjdPTsRhct
a6dcJiAERlIW+/sm9ZShRhCRx5ZTvSD7x4bEv/kgvhOZiSF4ZdovN3jEAEziumHEh5Wul85J04At
IQ3xscSOkG74t2puq+1dHAXLvSIW9XrJt3EbBHM1kcpux7AfWKGqUBJLQCWmNSB1qDbAVbMBQPSP
z/hWfm+5u4Hf8zmCuGRy/3uKRL6GmiFsOpnRIcuLay26T3FYrfRTeZqbCSOamoI5GiCBV8YYri0X
x+glfHaU8BIoOpziIdC0XMdJJRCeolgXLLWHyE2QvLPYFM17vvf+z5VDijYy0DEZeFbNqABFw7+3
N1ucaE/WQxXx75sq6UIqYV2h5vnHrQoaXD6BRy0jnH8pFHKEhdhYIrV6FvgefGdeNfRXmh1uZM64
we9V1LrYInbR52gbvhnjg1g836GQqpcnJ1IZk01DOixKaTO15S2ZzRnRvdY4T2rncA13aBP6fBTv
OIRoK4774Cf0gXIoShaTh6J5ZoQRNC3DluJO5nlMjdXwVJY+D3TkRQS9G5Mdj/nrElAyYATTHVu7
2lW8p1wJOWqWg+WkbN3/JloN5Eh2YEyMUNRKVthkEe7nK+kJcfcreuANPs3txfZPUu4dih9QroNc
O0xw1CnJS+i032FyOalnSxktCZBcTh1v9lT+vh/0YbmnrCiVXoJrR43eFSEJPmeHn87RBiyv4HEI
C0K9yL/l/dT8bEqE4ewkTv0IhVCG30/hvhmJdTcQAuSp3QdRm+UAHTNCk3obbN1xQs6EyJhR78tM
6F3APo0vAqtBRiRIctB1l/zad1pUTC49o4ocyFdeC7/mQqfjgVbm25yA5CM8G8OTAPnLaT9F/qPQ
Z7XGhRs+cbm4AMeKcJRGQGW8l9tOag/VS5/7YsYscHKksa1qCStsrVR8UGa8DMlDZNU/0+XHuGZA
Ms9yKo3/taySG/R52iTUki7FIl3ntTB4yuRF9EhR/cF9g3VHZk0sr9rhIkEXCobV2gd9PUweZmks
ECrIDgGSA+Lv9T4wWER1z0eIzuLiNt0C3f05FEKKlJtjAfyeLwVdjwF7eIVYc4SxoJpkLeJ5arDF
TSteEPp3IPeuH6nQDMKOTpPkcX6nH8qzL5hfqayqHdFOFPFBC9IQf9Gv9lsavenhmuWtDq4ie390
WF+TjlWH2I/ekT1l57oli4lf5mpEmwmbI719U2DcLwAgAXUANyMHk6RWlBSj2OSbDq5ts1y1D1UK
pZwozBcIERcAPttR70Em8pxEY3yu7b4JwJUhPPG+ZnbGoRlNU2jqMWxuxDsDzqSZwi+AdGxbhlNs
N3Y1vhBOi9/nQk3JaQ5cU6vShrpFEADxa9Om1d3plpxo5AoNXNslz22uglip+vkgJ/kixuFXwrff
V6WtEUQZIvB4pVtIfdywh4DWQayJPD7QIgweUeac7Bx0n8KapNWJGPBvH9FHMTinGqp1Ax3c4Ugv
Xss70DWxhWHN5qeSnTNmo0WY4/tdXMYYx9lpl3rzJbsdN87AgHSxNv20P5aJvMLNvDPqR4QPLD3Q
Pa7nValR22UIXh4sc1AJuEOtY4IJzdiZS3usxbvQMopq91ydY1F70BBWhaOaj6dDopnoSpbkUlv6
pGiCtF353d3gZyj6Q7Fbmkp8VcGLQoCIr6RMpi2mthwlWRJI9vsnu0PTgR1k4ONrJtIkefFMQ6OM
etUn06UY+V7mpzi1lVYcbPsRNjZ9/3OvTxOO51MA7k5+8Z7f5hjLRQl+YvHR/jB8Qxx6T0UgY5g7
PSvxMX4TCktT3Zo4208YImJwIWyk/OTYEr4i6L4V+S2lWtBSIHOhgsc4Izbz42gzLmDLfkesEqUb
oKTNZvRds86l3Ca7vhOLCvi1N3w9n2OXKkFuEazjf4ekGZAc3hLibNz+mM+iZjJdmKeqg2dEL/q6
2SOXOV6ekXdGLERIEA5uiQfMWR1dd72uqM8U3xXW/4xuBEu3+/WyM4RkxQVpP170Z0h+fqZ2YBKy
86e5hH79lYSe+AUUhAXsxy3DAFX0X14mDoVScFdMBGQny5Ef80+e2CP5O0ML8MFuEigjdCWCLqWe
FEvq+qnmhrQMawcRt75JSXjVbxQx5MYHem8J8YgJ8UeRbJ6rQnMpWUNLyBddnswx6x+nCgbJjoVa
SVJFVlhn0PFkwyrOGyJKMd0k89LpkGUAZHnH9Znh9fG4glKDjQHcjV3E+aiUemfsWtqWag7oNnJG
lHNpqju3Bvo359hnecHmcQHjfkpgwqZMDAHKmiOrYoj3HVmUM44WiF67Htiq8VXjoaaX3S4iMhaL
HQgvbHCz6skgmh3WqvqtYBlOi18wBSZbf5788GIxu5gq2t6zHRWq4Lgm9VM/IzRiN+Mk4UY58jyn
C/jJ0j/qwE8ixIVIlKButSvBdvM8VdNN9dsiV5MJX8b8fg1lRs9JnZGKlXSor6T2GSJ0UOMqRPB8
IYXTOocqpd7u2KC91Z88DtOv6H+11ndCinMiQpcbg+1cWtvP0IiPS1B+QuJTkSAizmTHT+dzaYm7
Q/IRfdzeU73vnfEhGd/bdL+eXAjhfsrSA8RPpANwo3fmbmY0iDOIv7wy2v2krN0IfKba/na0tKb6
3+LKumt18eZK6SKz1plqjZrLFZMum3WDHwZjorTBLWnE04JBD0xkgy8WltqisqayYPmU4rr63RXo
smOzWf+CgIcBML0x7WnlKrWPq/niU8d+xbO+KBZWVn++FzYd8r4WNyADIk+NIAYQologZ8FpuNzx
uF5qphlAu0Gd1Oz1n2RVjPYHi2iWb0W4AV/rHuGAGWto6lGfhE/EnQPcc+V/PORMr8rAcD6b4H8l
GWREoj4ceS71oAu9GDVIYe9x0I9AnAJmTyfav+otqiixBjEivwBuUaqycU72Tv730BjV6xXXSLBW
E3AY2XFHNd7VQxOzUn+4i+H32FLtVEg1b4Ru/BVzE8anbZSzy0wcVH+BVPjUqNCY+u6Gy78EM56s
2owVlmLC2HGfLLspk+/YiLTDhqq5A66xqarrnydShq+Ip1FUk19riz8QUdGjZIR7rFhZnQleGHqP
XDih/Q2EPWMntR7q9oekrX/hORDv9qejNnBbHODe4Ojq3nb6QUZnKkgKP368l82e2t0a4bnqB4OA
mQyiND97fXeDfv9FAOFsa/yHR/dAW20WrTRlNCb4wTL+T4nHHQO3m5hIeNGshTvHPrc49pAhAIuO
mpYXtDGP2HlNaGk0WBKyiRf9mvOw5ts1u2ekP0O2v9lvXHUY1etXC0az9aKaJaxIJOVHAVDdz6t+
8hFHuYad1z23l+3lm+K/7nBiMFgCc7UuFbdE9x7Xpz6V4A3g6fbmuy1XfgobGXRjTWdgH/aVIUMH
NJjHv6JjKU78waGvEjHVXPtAk1z9x148n6KrawC2mzK54y01v4cei2xNif+AUcPbzhK0IxgdcXzS
CceAasJ7mnf4+524bw/eNhM2UwYEMF5gcXe4HQhTRNEA/v3qabu21tE567sv7ZbWV2ayd1ZlH6gb
ZisRpdfhdf0TW42nHGnSri0UTX9M169yahLw7r9ed+/Qnxi5I7Pyb7KP+3rRNVxuZsilcp3+zWUR
CMQ10RvfeelgBXT4TOlCEy4hDg7OENT0H+uJn4hqmdoAOlyvVp0+/Rm3D6BBcXyoExxBXB1y384J
g5fiKJtORrqY9nTNDX8MPeg/LUA2GutqXGwDWl/hXp1PFiLfrbkqBDQkm3/8MBPwanAay9A1iN7/
w17etS5lD1ZSQvVxwazi4KzodSj0h2lXUBXz1xzqrSUD7D/clqsO7zdWc3rWzVm17TH3HIlAfDiv
vJLGTeW6VnJ2ILV4IZNExqyIrYiu5Ex75XRuHA/oL2ngdL6qynNtsi4Jo9Kt5zYCBu1OPDHvGIIB
QmfspSAkZJGfQzUu1kN388mCm59oB5YLrOeccTHPJedP6FylLf05qDH95xbZLMn62RrK7BEZrqoc
6jXnyQGPlx/HhirnL/ipiKrPBzlwXInBrwi3wgW4NkR5iptZf6Uc8kBFff5ciIuQmc363B7S6wEf
0OmaPlXLxTTqEPmIGprlY2X3PZtbZewrDyBs2/DIlpHIJeNzfKnxqX4i797HYrpnByLFrC5ru0Sw
yeOjXHe+lkeL1rPfu2VfVuWWWKvgKmsZ5p3T3Tn+0J1NxVVnJ5bCiVLaTw0FhwxhyCte9PsPgPJp
bytIg560CcycopxVH5wdjgdkz4nfR1jS3HLlIVDHmw5f0fAWbfwovm6z0idc3TPA4sdVAnWFQo/k
M6HEG7O5fl4YFVcyBtz6uPBDT7DnsT/gRto4vImlk/qzq8eF/gQm8+8YUgnbIQPzuzAS3fvVqKN2
DiIxOsrhvtl004+ZIz0GcqWztQc6PMvxUThh3Nfx90BZSxL3beEelpuD4U+hS8DeC1KwAdK+lFPM
kpiM96MqFFPX7aKUBTzx77byvtFJt/AktMyACCpYddcxALRrHOKIMnf8f0g4+0NywhK87jJy9VDG
mNqbCa/+Z4vpE3Rw6AdX9hVgdbmQOtxtCNJL6dSeyhql4TLKFcEr4I2F3IlsO2ks+0/g/ijTwcoV
TUFxXPQk0Saa9uM0WteBTnXffPxC2N5A/c+UfmD1+4s4aCftz5LPSrLNfuJOzC+lVKo4iytlzyFh
ly7J5rJHK+2pDP7cIeU+xcmc3lAEYKwMZpWSXrfB2p4pgC2DSXiv7UYQc2qlEHb76rwmSY8JWH8o
xO9hWiUb5msOcqA0luW7lBonFZv/ZbCWW/FCJyHDorL8+pLHRoDTqmYp7BhelOTvFcXQ1DTitZ+x
1oemwp33rifp9UXItmtl0P5ASPVYoHd8rkLGuzxO5HlD/SDW4PRO1fctU8JJdW1LuF6p/u/cElK5
DrlCJ26QpocdRI16yMEsDWaRGeQwVo05cCacigoQgH8EXjWF6d48mvm2jdGVFOMxN8PD/F4TkAvM
8di7NwZd2dUn7/2FtouwXIWP5YSQyiiuh9QyzHEwuN9moirBYbBXXLv1Ce0Q4QKKdZv/HUTA7UfI
3lgD/DjWZE/acypE79I40LYu70BNsT3MQADgyuWhsb3/uNJhOCq6bWSShsQF/FgVbWaC/aPiJtZb
ejqQKdCk/BffWZVG6dyGtMAFsE0GUtZVHZlZdt2kMHk9lJ69XrKMwTtgaRI58DOJKNRKjdRX/UJ8
rnv7Pq2jpn9oVm1Ola9Cbl6pt2iFTzMQq7f5XVp4SOUcjVI1zTeW6UqCCslmN76/H0WQBzXK8sZr
0vCyALrKscfaUD2WuegYYhOjUrXQ095oEq9lJk1MRgfzshMhx753zKqb6lt55cDyKgaEWPgFXW1W
HwjFTB2P08yHQNKa7PEBPPR0XqaarC6Pl2D+ksYlQs0ue9Rd7P2n4NjHYU6atzalTxhKlXg89c9i
nQVej4Ww1LI6ue3oCEOGh+DtxymVg3TQfliaeCN9gb7CHCDhpRd+bRLGP9XWRxbaXEdJ3s0OCotB
nB2R8L7b+e0oJ/7cdsx/GpeJ0fpJIV/IpBGcWrH0v9JBUop2sPS5TtBEbWoeOpakuTFAqTFT8G7+
svMmthwbJJUovF8o4193VX7CLhcwx5+6FE/WUc2vaGgxkzEZP8v6taQJVZkoFkAfgVSCXi4r+EV0
VFt5Wz9s32oaW/X1VleAYLMbUiKRCmtWdsPXCJF4mdwzwBVcTe0RyGaigbdB173guTLuhyymIzCC
vuyoAVa0+P+dPoyF5Yan7xtNItH9nVKofLn+FmdxrJv0mb7JRGqeRotBb1DBsbuD48JwEwZuoK6V
NElYKeMxtVrUYNJJanTtMLAqvMjEOLWmqevVIyeuwLDo4pgj55Px8weEUNfjFQtkGjjHD1a5HqAt
cYp+49saD09tLpQyvl9ScxqbdMZIxx5RBsmJSz16ZQQwJ6zIEEJ99eIblePwV4/XwVJHaeKzt9eW
DXd2MIlexvXCLNNx93Ooh3XE3gVaulrlfnFc9or303LR7Wpti/k+O84nqZ9AlLSp27Tm9sjlfSG7
+86oQkcPR/GxzoVVKrGrCffzUSu94tqaHCyGOW/RGG0iuPTFovRmX8r+4KMYCFHH0RBpofcntUon
ymwQedA2DVz4CaJPuPF5g63KkUXJ3dHn2opMMmGdgHR01Qm7p+DQnpUBLtf6qKGnWpTPl7/w/G7u
jSo1pN+PAdbBEJ+mR8bkdB8NbS21xyCfO9watolZO/1Ik7nd48Ho42RK1fo8HoZlWS4EqEjTI2lk
cNQF6S4CsV8aH02ISRRDd0YK+nUFga6jG4+zRJ/blIxegmT/gPY0qNqijfY6QthGA/cO4FqhCuKi
d2sqMX28pgBe3mXsDDDWY468DRwkzx18fj57nA/uZLxiWCKxPFZyaUjSNzJ6O4Hz5MGFoYBYTKEE
KSlM4vIZrnwf6Rxv15Y6abmZrESET3piSQ0+iqlx0Tv+sn1PjYeBSPKpHitQWTOdK0GxTByJOiV9
/9UXQjAGrP8gDtKen/RJzx+xrUFTbdeomTuE8iVeL00EyS+6jf8SXtUayCbeaHv1NPHpaAmRkDzC
p7gPQdGnD6u/7JWgIhLL/QGISzyJ7SW7367uoH6vcRYt52ajXIefhQhcCYrgNr/JfHzLCklYlYKW
GKm3x5n/NQbGICfoEibl8UxIRVkYMe11++2vm6eODKGULiOYWuDBfR374yo1kuPpojO9n6y1hRJ8
6S2ghmsy8frb+H4U6f4/EUhYrt8MlymMUGCcSWYVkD7RPE/9Um+KKNj6lJhWarrbmwiTDdtjW3QR
GZTbmJz2i3PzEfB7reM9PwoGLGUni81XeqVYSn+XvhXjxiBrsVWbaoyN1L7bIPQD8YN0XauMn9uz
+bpgH9fIjZ6HEgTSG57QVS/SCLohODTDD4H/wS2shD4bF7CS/P60t3To9SZiyd3twi96PSaP1EBX
8xBwmxu9TcMg96zwGl/TzP/Edfa/cpxzPMbtFk1PYdhFQoW2DycQqosOf8ZoQFth2XWVMuFwXdxU
AErPfErv9JVmT4BDZ9r/wZz4rZwzK69a28VL/DSNaar63aVkEwTAiECp7rMDnvEmhbak+1vVVtS7
vFCcW/G1wNui28BbBTneWYsn+sVqxXKl5YE2zkqU2DhQfcO6aGqOGleamRoqfrX9szfwCbkWVbPE
l5Fdxcq+YwJuSbufBaPBKZZpHbxy28n9zTMctdQWUC6a3Mo6YrCitCsu5FMdyaTjiGGxCVO8UfH2
a9JNRzouHQRbZoJdShc7jmTEzzmntAT6u1HfIltO3AoplqSEonu5IpPdho5Vqkeix4Ic8QCcWY8e
VgzaPrBVDZbAqNQDkKPPRyD36pGeVr9MhQgTNcjuYkddnl/QhYEhjo0DDsmAAxEvoBYqMPkKpGFQ
79Sa7qLh+gY1NY26MSmFuNqpweWl8hrea2VniOBoFbFwS9EfrLPL2A5GHyKTXAYHuE5dfJpZPL0/
xnUXcex+1U/68CiMDtcDJajWumExjR+4uWRoP9tkGDLRTBvsNTtz4VtmfGAN2yBZhkhIQJRh+g3g
ncQ/zEDx1kvKzxGwBPNwxCQB9PFU0Ek5wKnyPvekhk4Zmyzc4DoZNlmdUKP5opi2N4nOC9tvdPKn
3xOOKUhF9ohQHF6+JgEth9J3VI5WaRXZksVhyNUMBPCkZldJaapY1b79jzpOd3jlC08wgdTjqUOh
5r3lRR3TO2YX0tS01s1jpVIZQDIkKSV/XFhMs/6BoJBn2/D9qFalk7Qi2TTDoNPmh7ZdgACYhsaO
iSz4VttomRPhHJOygQSY23YvRrZyXucxnw87VQEdZPCDaojJKIf2Q4BRtll1PSVEQTK2ppUnW5eD
TzBu5SfSe9EmIe6kv1Y5F20CBjiDkPmDBSc69bxpbysXSRj0yCRHJ9KoDCDhJshPaTUuZNCJZWZe
NxQqX1RAwyYX1etQiFlNtLdbQAURiCn/euBVxlWsGZpYZ2SmXQTgNSR85oxx9tDYvuNRD0GI8obf
yqxk+33YbTMbl8M0Mo2n4zfGpr6PoxDs93GIlWQ2MXh1NSK7Vrj0C7KcSh0NrvYyvVMjXXyzlZBC
47KLyf7AQ7oYXkhYZZczWn4gA1h8puq7/i7wpcfTYYPhzDtmBjHcTYEGRYI+6PvfdCyqUZ7Zvg7J
fZfoYn0ObCsM2y+OHlGcZwmVAc9Nj06wV6CM1StsaMctnDIgIFITBVO4Gi147B6oAJckvQCnbJCb
D66Ve0N9NCmvkuHipeICS5kWZ/eswKoD0HJ5SM9q0QM6jmzG8ndkzjEXfB1sm3/DXJ7/Rl7KWRU5
ChkPWvQT/gD6vZ/4p+llChrBGh+dpPrs3RUdYlZm0CTIgb5R+7RJNLt5jHGhQAHFu/nkcTZzD1Cu
EpFJyhZ79T2UECZQLVXo6nJW7iSKR9sP7RAEH9URUGXyQZnrt+TNHkkzbcq4dyu3mLwCOiP1lodU
GbY3VE7aPLntg0uZ485WIq3hOZww/QBNjB5ZnRzpJSgrx3dX/nTjMNukeiYyULOcdr5rhgnAVIwq
MSsBQUHc7zqNPRHQXLLKgQDPjREg8b8cgHNzbZBPQoAaVWGzybCGgFa9ekMBfz4RMjtGDXdYhRwu
n918IwOiFAa9DaCXIQizBX/Uov+c17LOWBlB9KsPW+fqFGyt22D7b+nRj2TIFS84NK2dCNVvSz7x
dTUQVNrJeyCB0Yj+LdfON3c1MKa1e2xJVjBb8oKejrSKjga+/FvtWodUg48erWeNEacmE30p/M8a
TJJit2DncKbvTQSZF59LkG/74VnS5oSc4oYea1ygujauBIw8qYO1ta6Z00Uh/rg7972GSOJEj2jz
O+4qsx5Gt1x1On3VNIMi4ykw0p0/VfTz7sMFUVK7dPd1lGzJJEyFH2cBUVi+HRyiaccqGgHgnDtY
39KxcPdHrWA2q/qeu4ZPKqV7KkoWg7T0rUtTtWWZsh9HxIl80/vL3jyGXRek0bY3PPJJ8knNzi0j
a+01EM8rh4tEgpv5VXOU6EvgKBDkOwvoiHLZ54d8LBZfXla7en5+rwFpMASseXqyNMtHrbSbrZYY
w67DiVE+N+gPsv0GDAtwiuwyCUSUkVyZPrMXNKdzTBsQ0s087bFTKaBSZ0MSjLD5KlPe7Cvy6XFj
DmRS+GbnZFR/xwO9JhzN57t2Eu5OB3Ljx1jc/MEko/l0CkzjDkwhHqvz8Ftor9OQn88nIANWC9Co
4Fg7gdl3Rrvk+cu00TpiqprKIK1KDMbZLp/l7YhUFkNwOP7QEHP6mtnVfvUWaljwserd3/5YkMc6
x4w249XAL4sgvnkn2GAC7USpq8YtoqOiMvkoHtk82typyrwBmhWrrz05b3fMH8Jiw5D/oCw6uQbZ
s7yAYLO86DsDFwfq5YOeXfReHOf1V+1p0eg5X1/5iuWjzQRuXHelNA6WpWxVH/iIJGS5T8MRveni
KSfgeVUh646+vb2/GluIUjyCHcGi8MOf0vaf1BXAAF2mUOgvvn5CM7/2N3pu2vZEOjtTVkBljEIq
PnS4cJICjOII8wF+JAubp605TWzmM/JVpLEUNTz8r1Y7fgKt900pfFAY3492Fk/4fdJBlkYeiiES
gZ2lPF30Rymp0ftbI+jSorE6bsRi+mPrBpA35SsLzc4JNdEgLtT4Vfdte5Dvs24RomxvL89xp6CX
te9MvnOKOQlVVqyf22QRnGVoZEfGriVmsHO7K7Yzabh478u+SleJAtnoKtSKSV9hCLSpvWfYR9Cj
3hq4HO8m9+uFOlX0jh11IkMIUA5geXTp+pK/iZy7Z0uDFJs8Ger6bsiDnET6haA4n4A+oN2h96vg
AtNxxr9xFPDiUFD31CMqMdXT3HmD8aGNus8Af8rv0XoZgk3AM8m7BvmgU49Kqg49FUECwa+Ptn8P
NuUIujA0TqQn8pIEgN3TNZ+nZUHTc0P22XWhegJwvd41hLuH9JlqwIreveRMtYvoX51dRmINriq5
vk/5GkVMp/lJfp4mL5b9zqvtu5OPnYCG3xUykIgJBhVbuJ6QVPcbIt3Fql62vpDbOgA9NjmcQmA3
I47ta7A8l5qZcl/SHkYs4hmqLefbF06blGmxQXdP5b3A5rLy3kNW8JUhTHGBI70ZxNUoWZnC0VhV
qHpRAYHemCVH0DHYqfxAtL48YtT1Hnlh0RDRXeDqDCSnu6kH5/tNLh44S1xugMHEOMnMRmDkzlGB
0CCrM4QDjcB92fiWetyf18mg8dC+A28GOOPwXLWRUpx0SvWEUzHvvh0S3SN2ES+p+lJoHuGzjexo
yuhfXOP65CSxkjcECrAOacuHpsaOHjGWKfgWydVwD7iQ49pxGlFqD5dtfaKmg6RuIjyX3ALBcQTa
Pd8RgSFMQTh51poZWhQc+WRTsEa026ifK1N3UzxGYM1s81ZYwmt65AkWmUkjrNhfHgdg4VSHKUmM
6bQHhvNM4bEJRbAi624bcfw7VylrjM+oKWFDoxERwS/GG3ZWGe9FS0n5kgRJ7XGhpgmQ3zYI372M
TbpoL8pUdBz2QNRp91SzQvNOY1OAVw6e9ol22FqAKXoZNDLhxi/m6ht+Dq4LlWwmtRmUxVwRTBgN
IFQVEMXhClao2WtIhG56xBNYsCN5rz5c5UtBP6m008rnIErQ/Cp1Y0CRi55SAAN9KYD/mGc68Gxy
yrdKKWT6oCOCPIs0a8Q3h8LM+4ja0MXObNa8U/hhhOKGib0eB6UKfxIIcR0amml+p8RQ3K/rU9pO
WFpHBHrooltG/SjIyOO02koKE+mJVaIhn6EXmNE+XR98ZVPs8erc4FCR0XI43xVhuIOaItZ8sH2S
LN8uxyYEPeM3/r/IyOS5Ab+eMig4W1e9O9gNUlRfdFpZVkpTjiN+7RCN2Y5TZmCoBUX/xyw41QQx
47IMo8fRgELrKIWDa6BcGiizM5QjE8XDhk7BtNB0gdG2WosFGg7gPZU0QX1uCHbnO2mZHOwZlkz7
O1g5zk5xSUmSeTaKWZCjjWj/X5EM4Pht98XwES0+CSdLbc8q/oTu0damFAOZnCb/ftimpih8fv8d
aQ0T0xiN+P6Sa0CqKUqlLBAG42SIaWiY0VlfFIOBMvpYcA6+OjtncUOths64LcKJUCfpxvJpWTvc
HuXVFpz2st+URw3cTPqVEvhpfzDB/7XHo9xfeXSDjuzj4NRaFORHB9gCvF8JAPCXmOyo6tENCUuR
ol+93eV2u6Rm1Gz9LFz868uiLUKNvNxjF/XQqBQ7gNjLnzUYHlMUpWMj4dR7CfAtJa77zsjBeQPE
AWiPFkwrLnhe/FwJEnY5RDhMUoelclPTrgq6uD0/THp3zvT0GaehwbvVVvED+juK5hMnJ3fvezyD
c6c8z6HVdOzMEhkTo2tusd/uqo70zE/8E/WSOj/Osr48Ncjez93ajN6p6RlEOV0Gpg6cV/Yz6M0l
e43AWzVl5XLDS2u/h9tqLr2hFMMTq8UH1e29E68o/lHb01D6jaknA8s5z9pvfKXcZ+JDJWTD4OfF
UXNQ096ukuXoDfR2IWM0oKOT/AEGjgu9v0uL9Icdo+AFJFqCmTUumfBRwgKaQFyuOpIQRbaNwXqX
y6IfgzBz9wS/8nq22uGu5JXCcc0fr4VDJjlWd6OZZit3DelYy99dAdSgU711qOnKoItEziyQjI3O
/z0lwqdzZmOoXpBa1a/PV2yVajJkc8rG17xp1/xUJq0/TiI2H4q/haVqCNcgzFBOOjXgWSBVr7pN
i21HB1hlvwwa6tdU9sKQ8xt6dSismM92vDJ0oakINkqZUTpSK+dzk7bpoVlSbffme/N2z+V4FkKL
Erha+ikmlLlVQckkHjJ4PhyqxsyoyofJd1tjFB5sPsEsCMQpdX/hZvLh3wIspyTkEtVk8PUgP/XT
sN+vo18q/P3JPmC/04bDZh0y2NAYNyi/Bx/mgQEAIfZkyojdY/kvPxHC0dl4dcIviMAMmGXOjfnT
o71g+VYtFV+13onfaqeAcxGD4BJ57Ye5B3OqehvPg2PWC1hUz2nRzAT+u1I749PESvZNJuhc69qW
PgcRHftUwANXzJncHvulH3joRo0ZXBlpfV9BCmcNLb7rHGqVyoVrylPZAWr1YEPAXYaQRiXNUDNq
wMuXclw/+y6phVYMBg3h68onTySj9H7PmN2lBD0TsM4BIue9eA9XOBhmjsrjamx40ZNs8gx5Lwnp
vmzH4yROyFphfLMM/UjTzMj1Sb3ynsIUiFx3WLH9gmtzz6k0A5s87+pmAPez8YbGmZagS1tnus6m
nY/1WWopqfGRCTuGyjnn9BM1hf7Ay9JgyP7GUlKC9+ESc6SHldvQ2ym1+JtpyYynQuuC7wwPsxz7
HrpeBmJ16lG5+alVYFBv39ktO6eJbyq8UcARouQ+3CvKCD5vxdYWBeEFEc77t5TKfNlAS0JOzi/s
U7bkNoudgf84HsZR+EJJqArDLevvFdjAkFajPBSFvRg3hkRM0VNpzBHq3XTr+pMMesJveeDSy4fL
bkr0kIYTDTlKgLpFZn+gm2jo1djrtdMIUsT/9u+3ATR3Td/WGo2mRKQJwSBtgsiLumrjdujOtVnV
MW3YXIG54al3nRmBM8B9og5hEuUb7OB+8VpjlyhATrTcjFU/GQ0J6FkKaYFwAkRwRZh0mRFVulWw
+C3/34ftX0bBJU+P7X/vKgH/0EmXVNzFrzKk+umCR/PeCF7CXMPMC8kncAHnxDRp8bnFn8VO8lwO
chu3N7gCiHlAT/yfH52hZxPvxoIxuQdv+mGNifP1f81CuFU8KHRb5OPTNAiOvpt4vjxvf5O/e7il
GsygG+9e7AVUkX2oyBb5ycpMb7hzmRVKYURaFEv76Tk7v1RIJQzdJLIRrAUchoN/2PMh1hcMePXH
HxnS5kdXpB1B8qOsrPaD9QLA9/aSrY90Z6orGPcj2hpB0Ex50lYzJOyZeZF9UJhRIv0o3wyZLtkC
4HQAc6BoRXdJVlbtAnMfAK0/rq6tW9TNh5YJfEM7si4eN1Aws72sVCJHvlSeQ/D/FyjFfDojfK9k
kncb/oO8Rr8SW5bpOrZBBR/8irowNAPw4kwLrrerOoQBXbpeAaQQvJ3Pe450KojbvV7vmLUEslM+
yzEbvE3Kr8YncNm1AiWQg7f2btiouJmcEprgttnf+vybdvsH95OaX2oXLkLs3Q7enVbxIV9cpiSt
jTIYmoXZsOZiMv7zbo7dD9ArGLOTSZe/KwsLAf5fg4u1vMbSUtIB/0W9+0lW1P1gImQJAqdAvYbR
RQGpoM/phUxqnPv81gPtwM5krhUqFeYVKL6fZXfTgirvIJRgTbziCx+VTqOzbrNWl521sMqVIhF8
86c1yE19CsA0FbjQYLS2tDIL8F8MHyMHpo+LhTdg6s8dJam6PTxPAz7Ny+mEO02d/BRcOBGyD+sA
DBJQBayJRIg1Y4CwHQDIV7SIZNO9QTLBr7V29xWhx9wedlZUlsHAXmZGRKSpYQo58H3tKJvbSTwP
byjX/cxtMt3jbAwtBvWiq3335LN3pKhNm8tB/CrYOkc/OUXGbcQtVFLsCfTWFAJ0ivQzNVQgq8ue
yln+myVgD/N6HmE5rTKmHgQulC4Aerp1FfL5cGbXHSBqcHj+jltYBRDAWYbT7NC4hqJ8HvrS4kUj
qmh3vkF7NQPnCMch1CmUzYH9cEGokn1MfU+Bp2uLaqSApE/sItUTjIylaujHQ5WswPvJRc7hyfSp
fNHvRfcRKwGYjZb3gpFqX4V2d/yBFKHOwWYuGh9zvShNT91lLUYaTkrkMdMb/P+ymCseNb44gDwD
gW4TzCvULM9WL0xNJVqIsi7cvGdtl2L8Y7accAlrUA6d3k7usEpHQZAlC+vfhsJq1w/cqQ3AAWq5
TQKoaGyhAFNavbfkqTyGczdcoeql0DXwVAQmf8uIdpvZBNNYG3vNi/faz0ahbGmyWN/yjIq9A/Je
49nAtwqWIxBqhhOXsEVttpUX30Z2EAKlb8n04XYRU9E9YLlClUQE8Tvk/YJhkthFwBV7BeOywvi6
jokRBB+3GwBKVAjfeBUAaHWVXJI7dBe15+JB3ljWLcQNpxxmgve4ObpHF/BfTJNQGybxr2gczBXi
eFCnfnuWjEfuM/IZtWRTmFr1SXhCWmfQV0/wxd3Y0ZB6Mt6ZwlMiMjMTqhCx1PuoiWWSOtt3Y+/J
kS9zOlnrgQWOwsL5v1w7gE/uqF6hAQvCRpA6VgcucCUBz9TecKHYJK6DLpr8/ygPgSCh5xwiS41j
706diZRpTSQ7zn3aIPKjOsShhxXlfcRVfDWpSmwi2fciq8Shde0HJ3/0HJLg3NxbTcrswEZPSrnR
E0s2Qqvw2jQHHKLObrOCPB7mKsLRs8uCM8OWbqmuogfBVm3jHztvrfzfetDews5mEGsY5+KdrFrj
5Gfc6sC/WhMszM14D8Ove+LKJDqOCWpl+vok793MsPzQwQcO3G7ENYj3PUAZW2cT623E0kKUxKWA
5Ap7HXDsaLZkl+QmQnNbvgjHlb5WQpbvno6BNDhNYDhPlEC6vFt+02/b1cfLpWvHxnILxe8XQ+0f
oHtPDFS5+89FF9A2YR6bKPNKehRY2qlLdSOwjsDxJ+fmloApdJ2h9I5XaAp+GWjIGW1XwMWOYip3
qx7/Eoi5mJ/wD6OdHZeRsC3EufQ4etu6FzOFzMWpXfldzNnx6jvATWxd4kR8J1oIB8cxOzsxR0M4
XrMpWCryWlk13wp5/hXTZJtRan4sqpoOiNXXT+APjwEq00Ay24f5SUBTh5LahPY4/iH9Rp9nueHL
BJF2q3o85swY07g812lRN3d87mRwCABwvH7pjzpZzhQnhFfMVhIrvx/swsHhp7N75tsAnV4DZlEc
1CGGbVlqFTGTa37LhnVPhm9uya7fIrSbj5SnbbX+VmW2K1+tF2XB64H0MZeeZ+GmiHr3lCGMpBPn
fHW2Al4pvratcTit+MyMvRF8ECfjZmlLwr5zk/6KaB8wmMb4ZlVlgpF415JaDHmiYqk9DTutXZqp
qo7iw2hCCSXKXRELvTKge4sMy7SFeJ9V0Yv/trsPxvua0XINA2ytlHpFORNGTwKBXrOoqlhR/FaF
NUuQoYiegCpVV7IdPemhDcrtZvbzky4zGTjR93Z64TiBTDDDvmdUX1sqoULCCD4rQnKd+zNvvIZD
zwuFiwHhzlU0JbXP7DtccL/4CUFpdjmrlpwLXpTaXOz5ZV9iwU11mu4mIhczMfsxnQkhvt1OUriv
gOVq58y0ZbW7r8CXF7vN3yg1j31iIzVoqTbwHsTM6CcXublOq2nleckwyev8GZ7V3GvYp7KRy+Ql
whQx6yZElY6JafNvaVv+p6zmeg2GIjaxH+rNa8OemaCxwgKaiLXZr9t10/cY+gFoqzh3lqk7ysmY
4nePaPRzI2r+h5VIJFbcUk70Om7NCdufVRT0k1FMgS361F2YaGDP/Yfil+MAgFkEoND3WQ1og5CK
WwAwPo+SCN+TKjCVW8gVpRTCk1zZAktukwuNA66+mZ8RlDVkKc5WP0nlJLLHjw7HwzmwcaGT0/XF
KgvB6gUubDUlxz05MFcTOV4Wp2iKG9alEA4d6E4V5DGrjh53xS85RavY4dw+kK823PJI39hmU56x
gDXhH5yt6nV7MTQQ3mgkO3X+6zFad8oWMwegYWnhcKjikYmf5FuR8ofAjMR/YL21nTIYoE6UTnBB
F8wT6RwMmSF9NppNGgnh/1fSA1mAMqG6flWkiQpn/vPfme2yETf1v2J7ZQ3x/SdycGizPBNiHpB8
acEkYXKHkOLITw9nBk4vn0+iIyjXQznGAydHhya+twklKVE67yrh2PvBK0w35TYVE0k4gwY1yd5v
oE1VMzSwX0lQJ+mm7nUQaMhF/0e0u4dVw4yyBqA1HqLuOPvLUyZ+qDXPgBRlsQcNkw9rSSsrOI4N
fErf33LvoR5JB08Ycps4aR2IXK+tkat3AdtIN36CjRyzDgyRW0tsYR99+4Gj812AgmSV/9d+Y0Vb
SFZTq7Es93DKU9fxIMcKoseTouZGX5v8+SrvgvTq/Jp/Ko6tt0EUQiimxe8BCmzQErC5Ylhs61Xb
DZBcfj6L9yrjcM5Yr5VYKX3nBK4AzybjcW6RCm8DkLzYWzhXNxb2nPKobzElGcfXQZj0yLuNiLEy
CoSvXX4haVIvPDoVsVrrPmrslv6wEFluH4mgsyE0MjPbi0sbwGz/jWmXjw7j3I91uPslgEhuBcmZ
L183k6nvAHWyU1jo6eiPg/g1YQBsw2h5plt2ukYtpP0nJwn8kDwFiFlu8jz0YqJ3J894W94WyWK1
QCgVVAG19Oerp+2kM5KK4FeA4EthlbZ8DP3pg8Nbuxmen/HiMlShuTEm9CKbbUm7voVlvSjxdOyc
FZ18oHUtuAkg8Riy5jOPnNfUthL2db347ShlfsRHCkh0G++yRjc7iAL4Av6dQgurZgnuH+DEkii7
e5W2Mi7Mpaxkt0E4AiYcUzYTW4RC2geEDCIAH2mtHNCKsaz2GTPWMI7Fyg6NxzEzq6aobbY48Z4u
9fW2XMZ4WFuCcu8ea/Wzhcej88GMVVxECmLHY6VH/veBPX6c/zmkn1FE1hx3ELT5FNg+jdjX8W51
Rm49yfJiJ/PN+cnI0TYAWwSaniqMx7auyTf8/jUju8whXrUAY8ilkAonqzxJetiMuFdhDifmN3tH
ta8Km3XI2fgTgjm/eA9131MmVTdBjwQTBTLRqpAUG0lS+NNYwlJt6yI3Ehg3/SRlIHwN2ZV8bvu3
2rKz2D8bf6JQOoFcg1LCnaYyuFDxLIgpAb/12j4pjxSQaTTcUOaS+nIGZ6d7mNN0o26CtYDXUQrA
jaYdUADYKI4ks6/qSSdy04NvRuolkVIdWNuXrm+asEwwi8jEjI2Sf8rbvgvaM+JXL9L2iekDg/M3
PWQrxo7eteQEPmXpE81Zbq8N10M3g91cAfdU8Vqd+8DBcEHls2RWHCIwTCRtLHAY3O4IdVdrX07E
IapDmkvgZNPR51FqRcj1plszSTi+94oIoDaT+wwTsGRYxDCYdeY4SnuO1Gmj2lYBv92/m70hs5Bw
OHJfW/oxKgRXhjKDVizOQC3d8UkBhptq1sqHaIJqUeXB0VZjtf8AKZCh7BL+ekoBXJuafxjtu8DX
8EHW4v6IpOK6Amuvxe6rxZI5R+kg76Yuq/+MkWdWwBygJUAZz+l2wpJFLGDlbt8HqaunaBw15r3g
G/JD/1J8iOlVuotp5cKN5se7HtO42T3RygEC2bXzi2lzYsJqHpqqOuq54jbk79tAvD9lBQ30lw22
3EfFmQcg5hoMIEBjdZlvQHBb/RSubcEPunkCWTHqNsKngTofguLdvqG9Fs3MfOr1Y7d58VOL0+Qx
ERv5ygjyVz2lRKnyT2a2jevFB+fCkbesoImwFLFfuyFZoShnWS34L56zmmP/keF3yCfA9BIY9vd2
Mr9zLlhP1gkknf0+gvt8Ec21l6cmvfCw17U6nVKyT4Rg4IymMrsU0aobmZk9b+iHbWwN0wteq4Uc
84EZxlNJKAUjiMwnq0DUXolBkmRA6sOclI4eQi2lwEBByA8U2/23hItWLH7VDhMTktqzXsBs4IB2
YIi6IVLkb8ldTdDzcd+kXYzQAs9w9Ul25P3FNw5B/5thxp0b7cd0LYKs2lE0PvqZbn/oELaqrA8r
tDcthFGJ3U4Up8PibxuyWkbgc2mRAy+n5m5Mxulq9aAl5MQsVA7pHsLTE0tjW/M85yq+4wqHgGPx
qmLt2zoXHzAcRSZxR0GkmG1H2FVAw1YnxUNO8n77qRZ6EmTRrVJ6OIAdsk2YIQaiaEJqnFdBwMgU
03PrFiN3Fq2LMzMAb44dsVyHGxCEij5739ITkNPSlSYIyKMnjTSIMjCJ/xyFSst7BJLBoTXmUAQX
5Iv9fbz8QXtlHcLYlAoW09yDmZ2ZFRvfKC/wAgRsuEy5RQchnQ73nxLQrJzmMTvt+RusLsKmyOTk
bl/RJruurBflPbtKEUpRawpFnGbqDcTAIIfYtEis7U1BZ6W6gMRJnj6KDTRwF7b7WrzHVqgv8xZY
C5NEiqnL0WBmql694T+FjMYHUypZfwbuuqgF+lO5HemfTbUK2p5FbVjE1NC03NtX2z1mHowgo/jo
6/MGVe1MapuuBWqrsyGcNp+GZe/k5Pqd9zIW68FYjAk/FunWITqfhiPOnoFaiPux+nRi7KeK0a6Z
bvAW6XAv18epg4DQRciVEKvskHC7WcBhCBSQaeYVfYTElkKCqoAlPBFZN6iQ6S9pR/SX1ciYK2Uv
DJXQI/+Tz1riiFvliQBvkJDHmoDwc47Qhxx0yHX68Mpbx5bQIfboEmZfJkO2psgkm2HVEnQ9uU9P
+d1f+Ivz+yBIjD8ImJY5mn5xIj3v074ekfhrAIex3Th23oiJIjoBiokyqeaA66v1legB/a1grJg6
ZJp8Iw/W/F253nCgg9LweG+XVZ3DcHOrXrYIDkU303dndMxAbaYY1RKTFRIkXATZN9E+Tp+u+K9D
Lg5G+l9rca/e/xGWEzp6APUq1WKQ7QZQRB9EZxDL+8ni4ZbTfpyqf8bP8j55H11chJoLM4TD+Ptj
4adofygRk+yTR8PIrl25kpoJWa5wzZlSsaDK0p+x8zWfUuOfCtOpm1JaCzx+AdcMLZdsHAGWxbBK
9djwlFlKRoJYatjS4rYapetbeyKBsYkb2dBoGbJgLXTlIE75I4HLoFKkXkwNmZcUfR7tHFaxbMkf
oj0YoQimTo1JpHvR0vqgSegzLzDC0WWIHV82xqLFYfWk1QajXZsMJR+s9+TsF0CkeRbnCbWo9BUf
arIjE/mRe+/cFZUchMAkiLfhyhgzNQFk1ZGBl2DKxSHDcvl4ue8KxyJEXDdVoORbr7+CmZ7QJbkc
7b7ACFWGNM+sRyPK7w54BZR+8bMYjMev9TQCHK6Z5Huq2bQfdEKnpcNWHwmj11qxo+fYDfizUDrb
paObIhbAxUzk0mdwIA/8lpoBsMplUiMhqjqAuReEDyaEfIU/vW5NiCRgXvH1ZzSk0/K15Z7m+Li1
uzeQhm3sNNKeIPLpz4bvfl/xOgpDqXtefHcoUUQt828pWzzeRuJN/PqGuhlGQsPI3v6zcJyHCeMg
aLzkMBx2EwExF7+jYeHfU53AsYoumuX9sQ3Bn9QZofLUFkIWFZW7F/4LyaixzQj4KT8V2DZWaL1r
O00MR8rHbXkMuy7cBhu8oJ8VBVxjOYEkE6e/2M/dj5gckcmjpQpTXZRU3olSgaJbMfYUKcLK0POL
Un3hRtE1abMmYrTV2T+Jxz0e1RZcBUXTChKVzu72GRzeqgZyD05AqvxS2iQsWJVgs7kjnflJoxsU
OPPnLjtZHiPUROxgre6aMGPm4LRIgEM2LwMeKgGg0ThAGo7D8T4Q9NR3fDwDTD6/Ibdv2qD1xx66
FLdPsPQ+UXeF2rXJLXWznxgA1RaJPpwyRQX81ak5ZDrd3DeINowA6PbJtsI0zdTBTPbzEwgjSc5a
DYce+aWZzTrsMQfGqO2vFm0O04uWtd8xCZPLD79Y7w+n6PzVlxY2CaAy9V8t83UnY30jyug/m5w4
so4ikgyssdtGqZkk6GmFUjcmG3/MxTnmc40iF5rSUasO0k4lG6WWwUafe3l+8kmvuJmozOxFbRMX
qxrl5InvFaM57cUQsCFeBJC5ksvPmPoBsrNfXstH6+AkaK13r+tvkdwqxR2x/HEbY6iOdPaNgGr5
Myrt9JxumkfjWouFFXLiRmGUJt3WsSPRISgnUDHymoo8UUv1BwOt+RNitScCIDRVJqVAdo9vQqyX
wv+0ossjvvHmcjp0Lp/A1FhFPXud1E4+h66lXbt5WgUpamzvboDlAQVznGQhVRi1Ne/PZXer9tIK
BpTmsSO5dBHutqIZ6uM+JKoSn0w2EbJHUsOyB3QxqPL/vDMiV8GV039jcXx51esQvm/2TuBFAmFm
eRr4qZRVYEmi2ELE3AYvj3nss21qW+jHuPT7AYNEbI9wVgVEOkHWuNgFS7/tr5/7ChToP4uudAHB
VjChrWz0lfDHHXaG1TlJZSTVWx3jK/NpMvFqY3tvj5bYpRm8dorZhCamQ9QH85+Wo/5mY+4PISbx
l5bYroGgJNGJNbrraLKuMRdrDylaBHXMBUXIESO+xpQE2lucfF4rni/CAlm0fxZV3E2gCwo+W95i
Cl2cvCXj/1R5PBZhLp5kNlaWdZrXfrCAAVjq38+urrUoS6A5mB85umVXK17L8j4UMF5ECoAZGCC8
4//4Gd2p+zFZlrKgxzpb6oh4+3IrzPdtvaETObksNluZVctMIwhosT8pjjB6p2FRtiN/SC0h+LZw
c3+jAJhW1Lbsm+1wTeitxAIYDYWszPGBPmr0wYXehmNdVeVqs3SkT9TUvKR8o8gcjFUUUZWClmY3
LazeB5mkoOMiSxi0RuNwdxhn6UWW0kV/9/TRZyze2/oidCicQthEpUzzPeWS5fC7vgVj2hCGn+kO
11dnlj+kzrR3DVlcUof1mI2Szr5c6Tz1vOHrEC/L3n1wxX6B3aCwYQ7dFkZlEhnx7ERSKFBxQZJV
mfpypeaNsSvbtOsX8fg3MonSEh4OPFp4x72f0Nqt+bLpTOkDySoUoB5/HEGFbgh8RtTjMzp19dXL
+3TT+ioGU8kXhnE3gJWnhsNNW1eyxRlqFEtI93QVk7+YK3WSsAtBYqxdxHmOHFz9Fr/k5lV01/p3
vf2W6S409pkR6wwRXFnKayQcprDSpSrnbASvCq4xmzKfhEWTR0SEcFUOKBWhBsjNwkvr5DultlFQ
sQhfYZcQ5RbVqEtEJeUvFcSGdaW4gpNnDYobuQ9p/elifqXa7vQEVWM73tGRxN0tXBwvxUYhjkd5
cvKSEpx6mYn5O+xmuBm69eEAwPD3OrFCkThz8InSTl4WJ/kliEIuxfKWHbr83OpJ8/v4t8AaJPxp
fVX1BU8sxVWWsMvr3cRrsXiVPMSizT1+p4Y9nRVbl6wcG8NqJ86u6BoOpqm1Xhaj2TDHI3EluJ5a
X3Svas5Kw7N8RMCuosW8wWiG8jbp2WrEXXBgZtZwXO23CZmc//rQZ/K1uEXqip1zZ+qseF1lMbTL
Sd28nAeKNsCm9SfGC5jvVxxIAXlNPhQhLH/lGtrFTRZWeTsNUShg7lGcuT3nuGDwrE1qCUb3a6W8
OsaOKLSVk/bGbBR8d3dF6Ubi4o9GZpN2OF6O5NawmxPFOkq+0uxqGOcPGaSGKOlp0vVNjls/G0Hc
DytpSPIjFU5yLpD+8wTzhY+05ON5hf4grkrmT0+ll7Ic+YYwfnh8FzT8JF8xpKX1BTbGatV1WaON
3RfDMglODjelrcQFJug6RTS8kHM4xxDjJW7e3ZrKBOiVraOpD0P0F25uq9rXaAWiCymvdDbmNJh2
VPUeNauGhnXcIgUO5avd7YGaeV5C4v+RYkswsOdb6gJzNbZ03Q/uX4/t7uwuFlZp2/QVRL8zK5sv
zOIS9QfXs9lSvdGJSG/X5kA2zg1axm6S8AbD/7Nq2uet81aITgzrM30keOJIeOdJH8al6ADIEnYQ
y/dlTJIoS0Rz0jlpikZE6ou6EN0mj2I41SJhq9+9LoldtFPlnSn1dF4gpY2Xt6mjrsS7SXgjK5K+
7ROfXcsixwMPAh4yF9BhfwEUjRUaCKLJtLEPNnsZrY4IZJOrnIEIEq7/K+XICmu9UvZWFAJj7Zip
Gkr5a+26XqgQSmUBj6jJke6KpWt4g4fwtbOIvNeWkND8wSh+i84A3bw8qAFkHm5O0yo84gLjYyFo
OD+ykVkbplIC+U/zXV8OvzsDwsEcA+n8VFrPlN4PXT5UPdWCagSQ6APBoVql5wMKJCF8uKB5C8dt
O5DLsIBmaTfPDKNgTvROwSIyLONRfhjUXTtsSip2hLu97ATnKGUwEaGnWs/ESJ+JxvhdHm1tuvwF
Re77g/gvO/bbphfMpW88JKPDuC42gG9NAb7E19v0yhmd3q5vgU3Z0nrk+OTV96MbaaTM9RfmUfDH
xGUO9UHD4KqxJwvUsW7e1eVPL2q78CaG/4tRm1VIfK0pkteXlERohUHFpSpa6yeKGS8WND6TEev3
GUWQSM2/Us/mxm7Sa0PUwrPLSdYHtmfprBF4okltZolbtzka4JpYa3krcX/32E0aya5cbWiGG6Od
UfgCcJFjR0kymI1NAWS7DuajTffT1/HDeHp9xGfGO39mzpSqST//x7rz7PrddUuC4mA5FlKc+iOu
BQUOG+fsbBM6syc3OHqH678mRQCyMMbxCRmkaxHmrifTnrggwxbdeEHpZadFEIJgzPSTs3skO/Zw
ix6sNQMfiBvDqnBAQw9m0hh+Tz6pLrJhdL9PYI+0yn4YRfcFOVWdFmqEmtTj9uG4y+/RXPgLQRU/
Enqg1qq6WUCNer75I3zzzS6X9t/bNB2GMu5paY+4Ak9k1Bm6Z6aM3b5j4AOl1+128muctidb9vKE
w25tuf6qxHbQepPUCFCiL/gptYmwmjOpWRaqHgtcjF23KTaHTpRd+c2tqFL3UnhFIFbJZ2sk1oX9
5o9toMWWPTuYLg1F4VrsVjw4cGRawqs+fGsXQ2ZUG2smc/LrPh5NqYRub01cadT8qe2zOZWN3ADf
S0VVX5HhNfrNdLj2+vDxqpNSFxmQ+wxWWrcyvenZRa8wERCpi7n7txfW2E6Dcy777vXyFvSq0z4z
gX4pVvzvlSgD2K0FuLqKh7oBZ0WyOqb3ehGe0SdqNtnyrq021LmjyjBlhA/CYRW7ymdxiE0DdpKy
MkQUGhcMZIm7K3k0sYx6WiBQRQpwpAr/e9xoswWzsDOeMeajX2jrfAK2upqoHUXyG7kxRYeQ9E+F
Tj7dhU8ikFQGtNxUDO+P8b2nFgDzdhwrF1JpCK689MgUcC8gExNLQqEn0Gc2sZZjzGfATIFHsdFB
7Da+9nHO+K2hNPBaUgn6hxVUEXfak24xkqxe11DMQyqK8+I3Pp0qQ94HEpZquxSqsSAm0WJGekCe
tTlVrw2D7Qp5N2VpLTKjtEse34Hglg3K8yQcSfGdrB+Ae6vxwBI4VU7vuD34VZGEEA6VFnvsV600
1V0LcxP1J6cMU1VhlLbmX7No9UKDiE4VLAZilo+jazY+I9ePdrUKd87ufTqWD+ByBWALmX9VaCgp
hgL6StRtUEWZNWa6T3jO7TBH61YzuM+S9gckZEBPhTf+awE5PnZAgPsiOYMgRlKkwtpLGI3kZ5kl
QlJacz+hrolSUnRl7etewsNTrwZwa1U90N2Gpdletgbu3YkgUXhg1zfJjVkL4SRDUdpVnVfP58ch
a8A0vc7XYzDqZtmPX2dedn40I/xPdZWn2fCq3DHs9zUkCmzKQWenUkUzCNIXHc940CT+ifhVj50C
E6NVwo3IY/i0HYacckiEfe+VrzqeNdMkLswqmT+bdQQx7o0DDbi8pEVtcTNOnsRAVuZxireTaaxp
5yxPCZR2F4sawJyRQsleysPot5F9ydCgpDAGHFJ2DgBr94XeQMzz/kq0mpwRoGRs3+kSfJsr0zU8
aGbGYzekObu8QFlrB6DFGlf5W7U9HrtcMyASQhesqzFQn7QTw2TnVqnSJB6Ii5r/7e41wyYajlc+
ZryTU0TkyM0v4xLciJmSTgLnB2mLpZYKar1vuFUQ3+gqELqs730f7xbV3WGv8Pu+Ru6tUtpTWxL4
cKoZNnA7ZQuzVJSSNmZbtvyJWa5JiP+xkE2//WSS93hozwKkmjBYlltyb+0fO2JqPKLr7tcODfgm
qP04fbet/U7ZiM4BOyDfunBLvNKol5gPapl/4TtLbqw1im1V5laUmdWtEVq3Mntyg7AtateZOFLs
TuX3xvCcRSrps0UcIxtuq1BFJFLziDjCJy7Nx1DVRbu6LUmtmHzuLr66RsidAb6NQjhLM0NIJNVV
9zq7deOpyO7ElIuifkbQkzbWLalMxmTKNWSohir5/+aym9nFkpTnrVR+JsbFL7ZKwuNYLMk2b9d3
oNGmGQqJ7CjO6GEwbeurNuifvjMl5vKc7xYxf+E/Gkqb/n/qlWbMlURUSyBwElnyVnIBIsKH32af
s/U7ZJwy3BDCK6D3Sro+8mmyy2kYypIuBu6QMKSWzJGgDXmY2zwt/JxhpUCPTOu/iakgqY8lsJDa
iI+M3I3+lqv5RwwMDbzNo/PsORotq8tX813tRGMQP7SkVVWR51aQRg27Zf2aefnI84ZzQpmO/EyJ
LQW6t4QGFbkTBr3gqjsIXL3mGulwosG0vwuEUF+MIvvzzvrJZhNRgvpvcKhScyjAuNAIsbUSnyLc
BlDrkdmqNqqs1mEtwYnMhAxGiUNLJRRvGFbsbTRC5j1tyRzlwQBuWGDg0pQsiMSqt/HscHBrokKn
JSyr9kFaeBPVlnWzrQ750CSv60lY7jv2P3SkIZ69f5jV8cCYvbMND7B4lX2kjuuURiBf2rzB+r8t
wz5mEjpn40HWThK4SF6qiPSQv+uByuCMydnOsTKdR1hHj05eYrjFYukCCx4ixzLb72C6VyH170qv
mMIWYU+wZV2i1E1F5L2LkhUST/9is2c1AbqGiwg63LbN3yjKuBKsIc1kH8P3cfvaGkEVEH88r78o
UeM3fxka7Xjt4MZB1sKArT8EPyxuP019XxT0ndteLlaiWh6N/7Nfxm2taVdCd67lV7oWYfa3ACWv
GPgjynUe1od3XUYF3cNBOJZlAFSbM/cxtZXbTk7sC19R3s/U6ejvS+G/9QXf8XI3DFdFtFnNrUKd
EblUEqPdZxzLKu1m0DvY3pIkpWVTyZLljY3XN13wqvKbsJm4IVlWmdTfuqmdREPnHE8My1w/4S65
XbFV1z94M9SXX12lafbxZBPlRja0sQtYoxzcMpcGVgYDLaympw4DqZcmIhQVq3OPrCg5973boHbs
S3BgtNoDMIysr9TcDcPImlGE+bSeg83QCMsCybEoSgT+2XRkHQoAXggQomndQqz7xSKDLgnorKGY
mCbnSZpweF2Vjtm6hZmvqLrKS6XbwjFfTH7pOyWmTg3vhNxotUjq6oR85KhZKOcoL33T4XsONxAV
Jmb6Tva1TNbyuA8FV0Zng6VcxdjLMKDvrPqUmWxrAlBElOSGNx7MbNQxFtTDpkXLlZgJ3WPJTwaT
em75ugZnxFaUmbDLu4KiN1V32dRaXpfxCUu3cz+3zTcyUArJCE5LW/+yovH68wEb9Afk3HJliil1
eIzNYj8vTx6c/51rW7S8JpHif+juQNO66TLE3vQ3U6ypTNYpY2sGnGxPqro4qrM3WUjuV3xD/l/P
tXuz1D0y8jsDdTPDhMfn/TVXsMEpiYKf8cabdyoktQ5bso4V4tQboo4c5EV2Pb2QsRQhz8N2K+4i
xsMFnQKjvo2iIdUP2Sfd5mCxPLuDpIeqYB+LAIENLy3bZRpT6ekAKp/cfYbrz+TqmRvvWBFl8+LC
yOlo6PI52jtCg/drkAfKnVRnsVq1w611JajRyS74yVhiFwVU/3spsw8+YQym08vIRUW6kv5sn5jE
rIT24pXOVckV3n1yu4PxV7qV6LRcdMeoaxEasbW1aZG6z0UD4NMnuKWzUHs7jZRZts1QTlQ3Gl26
HI3rIuxRe8SjTgKXq2GmAsnz7C9QMIv438N+z/ZLSnu6GVGn1J8e0VQ5dAXLiCHOU3J8fO3yuN3y
1RRRYkNXFEij21vgaDjDP1LOmqLhUP/7y88Cy/4nvPkvsPVruS4Ms3GIziphuTtX5yYpsA+LaSnd
rvMuwxVbsBTosRbJsya27f0g77wzq4fRFWZcrQPyfXPAAb6FmJOytrNAZjfd+tjSy8HDii1JM6+p
bRYTdTPiRbUx3CArm+mpltOAsaUFxZeg62CANKaDs4SWNUi4MD4Q3jIQoQBPtuekb3ka3vDHSQIe
/yed4Yd7KrIyT6W/8Dbmad7uP2qiSHZJoQsCiQqRgDIv9QalOk5R8BbvhZWjc9xUu+8gP1HQOpoP
827P3oNMpT+NsPhisF9ayDGchwcMw/UfIe5meOYdddSRQixtI6YNYBfZNWyST1TEe345RGUzGVR7
XWYqHggaUQzAV5lsMIAZMe1q2DNq9NCVQwlYw7F/4GqTUDlWL96gMX3/qMCH0ydFWLyryF67VVON
swR7AqPv9U0LPy45l7ugUmxkrecenxiGgZXuIWohZ1f4FO9uR8GYOslJ3NtFaOSGJeL3YLbSPAsc
oHAiEo4xs+VGcF1NxW98WEW3CHOAhGH4JUnysxyzG7qb7CIu78M0UYfMxBSaZinGNEAuIQ5FLdYc
K43ohG0qVlURC3eJHX78FeZ5CrDwVnDD63Uv9AkeraceXjwajpQz92mYBFkMC/38oslEBRGxc257
xv87yx9D7lV8EiErB3fSNdaHDrhNOlezfFrbStD5khgJ67X+O+6mr9Wdb/1jtBZ/es6QWm1i+uxv
ONqoL32p1O6g8IS3Tpn3uQrRjdlEno2SIE314ZToyqI31FYf7+uLawHnVS3PfIAZZVOVOPmjKnGe
adpKcMpjmuCtW958a6sJHj5ebsnvNIRXHzsyd2GhPMiKOEq2peYEG5jwRD188+0nN9HzFSIdcoLF
Mwze/2TpDSCTsaErWNfa+UlDifyFsLXNNClTbFQVsIrG8iESuOFJ/VOzdAIkPgyw6NvvdAY+YiYV
utAJVuhH8h44xdXYDilgj2GTwHEkWhdPm1SmEG+ETxOp6WD3kFbmla/u2jKnGwpQFK9kgpUR3y6o
8wtDyInnLj/LPuJgrLYbfkzc6UqPoKu93xlJ50mQVJddosW6OOR+SAG6cNRiFIQX9vXdAvwAmcFa
gOzlla4eCGPnu3XXAKCs4LvxTYHuhLm98fR2jRRiVMpf99XPOToerBgXQgQYBG+kkYoC5fCa2eUx
XX6hqW1NXJ0z/fQilIu7H/1TJnL0r4JkXJo/1HDfYek2kTAnw8bTgvuwoJxy+Bc04CyG6WztoPtr
WrpNFY1uVeziqAxFVJBFs3tJ+GCmmtMROUKVQMFPQY4Bt9387wE5xjN5CaiOgBUkU1kX2RjXyM1z
eHDNbgSulfuABk+Wk8N1Ed90UXHnIba8oDrAE3grsdeI/srkJtV46x0stXTwTqmS2b31I/65qLe8
SLcouKYP6Zl48KmJ1/5HHsFx6BsrTsXVeBLRvIpeEiLovyycUfbKd0UDOI5YJ+h7v9eD1yJj0wI3
F7OfFvYepQXr4lUTaW/BAPAjOfB3vwLBrbOmI1GaLEdXwJ5EXo4jFrOTsbv9fvhpE5WRaMuindHJ
DZBX36CvuDbsfM0Tz/8W1ickSWmmBCVYbL8PMh6+Cs7FazwXthOraQtARe9hL0dAIa1xUuxjr4IY
beEE60YDKomPUtpcQ8Go2xZDgOPn9cv4lQMGppxBsPYECdCHA4//3PQvGpO/s9K5aR29YO9QTQNf
INVcWwiWo8ggjbdojUQYeO1BAa/UOimPF5I2se3fcANBfeLYo/4qEnST97v2IPvAQQxL9psviZip
QPh5BWAQLGYpZS3h6W+2iVlzpniN06Ah51Q1xN9M5rXuuW4hIp2b/UbkPPWKzMp4X/1wExvQRcYl
aN/jrAMJ0MkG6+J2TXGnkUco3/enAxCk2lLxgvgp7vyx8ussYxBzNTaEtBqJYKU2NK0cZSXD5S4n
f3unDxwa3E3a+YWp3+Sc4p2tGAxygvjD4Rd0Sv33vgn+088TTrnGRwTOW9XLu4AnvkEOXpxoz2P7
FHRSpLSK5mqikDECZg19tT7PUCWPXKb8Blcom6zsEIrEPHwK93w3WCVPpSk8UcwEd0p54CBNCpdr
MYp90msfRZ60G056Of751yR6C7kyOKAkvP7CacjYhp9Fbnc69sgopUIOCZXeq8kh463l4PlmW8A2
WluHHKABGRKqBGfPghDae98yNhpGoIRPc6vsHEcqPv+0As9xlmrqfapCGSykGTzo2q6vdgaWN6J5
g1p1sAi51klRmUP5qp55WornaIsIUeLOBMY4E97albfWkc1WZYOliejjgMevtYMXrolRAr2wgQu0
/7S1WRiDmKZm+923AhO4zFbZ5PHQHpnucN+CCC8vRYbRCgcLjmyTBPkj86WFUkY+3HzeISf3ijRF
5JZzFEWuO/FHVFI1hF7eC9QtLrMXFQfMsaSaGiGgF5FRodKwzA0VwmKfTRzlG30TVYx1pVDNpnR3
5uG065RhwdmqnlcPVyfiLWjue4b2vY3qL/M+oaKOH4CQ12arD8flrVV1jv7vycM+Rm4i0blLIpcz
zTWtdBSg4M163ZmTH5/Nxs4hkar/YRI5FXei7pcCM2IUCCPo57JgLTVl3/JymDR029dKChmhiYPE
u8pItKMSpel2I7+pvtSE8ovpHfgk71y8nVEkByw809/920+CHzhtyIu4CX5R8dRBA3STDbZCtcSh
9esERFSTiB4l5uMEso8Iel7WWggVn0YrhOW2Lc+DYPfhZZ7TWIYv6MjrlJdK26yK44eU1tzp6Aze
AMMGsRnyRpuaCqDrtDL42qvca4QCmKkZRfYFjjMJZYRC6dCvbAzSK3QfqL+EEVw0nfXMcAlhVLSJ
Y9f8rU3dIa6BlQ9wCpDX2Nimy/sdKlnshX6lQyBctVmnzyrVb1yzDrg1tHqn/a/D1WYeYqO/i2iT
Y5WGnYp8xZz9/fQNXY7G2zK5F4w8yUNowyCO2fpgJM9IxHri3X3KdTGWr5h9cvHwUMCbYLg4lWWQ
bMKlwbVxpXY1VJUq+rbSmN1vbfzEk0SJuaV6khcqKmMbOciRdu5UsVZ24+Ek38gcq6dKdGCzQdf0
mEveZ+KMiHE7LfVBQY/KmWRUaGnASQx67jcyOQlukQVg5yeLydqPg92ouL/MHpIi4Tz33arxbJQ5
QeK8sPPtTKuRPXTp2CVQ8wNllgAb8Ym0r8ngLmraaXBbnU7QGCLjY1zCfZrZmbBlmQwXOeXN1utY
+ZdJLJYBgCAEAIwznL7uN+RJpYEh+6kuyWebdIsdSOZ0WqqRUrpqExVWKJ6wG5NwyLRlzqRtgjTy
xv+zGVvut1oHT93yGpUJyq6ZsDjy1xAGHNhNK25qOdq/uFT556PhURZX8XlUmCe9L2gCRRzmQ/Eq
OK8PzTJk38OUy4KEK6A87J61mK0RDA1vASp9ywD++y/3yWygA3I19FRxYHHk+Ie5Kw48RtfzLlfi
PwR7W50UQTz8kcVBun6VWnFBS3ExvDbpt3IdDBFotTqhlpPX1YElFbMmoE/QkS1qjI0NvENTAhKg
F+GoukbU5xQHXwYe+7uZ0rIfLlo7jf2Sj7IjtD4fUTqb0s9EUec3QMa53UAKAwmn3FmDTJqo2GiL
j9WgpNUJM/644lzH48fOCgfSv7yBnDRkVO8ekDtxxcViuDnrty9YtZG8MCdeCz9KFr4IDbvkD2Kd
BAJwPcj/cWLmDW35d5Rbf176/nrDv6wJF4B1z8cTS7KsZMAwrXhWvr5KlLuRHzlsrxC3HQ7dDLXF
ky2JZ34L4YOC53JPFmR0NoACJuryPlwrDeGwc/O05pU0XzpFP3TUB8OVMy6zikgwpGQuUycmSGmH
8y9N7x0hfy/TB4VRmpDvmDQaroLPbmGEJ32gZn0z4h4ax4fFapN8oopolakdfyExwTYIYbHicQWu
Y7BBLy5k6/H00afcQurqcvbsRhD1gYEBaVB/wA/FFQEPOvBY5FcC2FSq9Yjls885WMfkNdCtbtwk
ipmRXOsfEqiJmmdLbuzAiUrwyM8ZnxpYJqcGqrVpPHmNFhCgWdar9sA8AIeGelbdx9rbZVjJal4F
GK494pHDJPvp5ubrrhVHWHXx3wUbst7lij+OgU055ARcuTGN7Fcj01CQ1dadYmArb8GcKiqAFL2X
Irno0skm4hGdM3dH232i6MwVA8w/+lYNPfeH29AY6aStARLc3qkWVsQiHPyNH4hGU0/EETv1jlcg
6WTozxU0YOU1fFy9nC2YryZQscFB22TFA5yQ+MeewLKguRhTQAJXFd7RmB7nzJvmqWF5ZllJD6ti
505uQUunWI/rlTBaBu8Uiwc2Rueg7N8Xa86WHJrFls7frka92tPWl/+DzahNHZWwncvTP62EX2yj
rBbGwCRjo000o1p91Wm1/X3AvspI6QJGnp7n4dr1YrLiWslGKeN5u3kCqd1Xzi0CFQnNCwq9Y9x9
BOmmVNMBDt+Cdw+DKcHJmngqhghMPSRJUgxBEArzm+ilh/iey4q4lBnBOZosncXBZbgZbhC1BlnQ
5P8bTzaC7Nq6tDN1PTZeyVEPD8waNwnVCPNvE2jNwfbcUDdzDBryvhNrxY7A3QBF7cAOV2tEYyDi
32lvQ7PbYKasNuTq7NVDEDDBWyRyLaI8li/zs3+sYVE5bDQMCXTfBkcVmHaeBQmaaYlGu/9pKDe+
Cg8px2XP+26uYv0KG0D/G51zcoVzc3C8UZUSIhF5lEuatdUa4ZgSR52eOHzzGLjfCDxEhL0UYd1V
N2QzBjjVnI3hcL8cIQNvfh3POQgcUplHnLYSjWbbozzmpSUBzrcyGW3YGPW17NR6gKtU7RS4BKOA
2M5ZrGNaW5vXJwiML+FV52m4ruRStllNKiaNqMGO2RFHKvvFq2ggrARu3ZHvQpxmeZyB5l34UeEu
tDUgd8fa43Zlz+aZ7TLqfLFCFXa6ndp56hQts/yIxBa6EMWG23sLHF58yBI6g72Z/G/uS6ycLCy5
5q3Lyvwju2Cw2vTDaQuF/Do2tape/cpwPSixKCvUsqoTKkcYuTQroiXlGT6ZXhTy1Si4n2jQypxi
T7yirn1nt51WS6ki5zrx3fhvyp6CYHUxICXu084s6e/AlEPpI9AFT8aQ6MJWbWl4y76OMGDXRZ1i
8rppWvLRcSWSVHR1PhpSPU1JSJPmVB7Oy5YM65oy41jJj6G/B+uD6etIOoH40cOdAB1uM97zNcO1
d5TSny1Vsthf5y3/TbJfYR6ZnTvfo4Xei/m8J0gw0Xd+hZaxxAubZmmZxVyuaqu3wwY2LZFRtq/B
q7gHdICbLOGr/F7K9SHTR+vA7QXaBFPfCyok5y9e3j+1XFWvP3rGCrHcXpzhZJDWCyihg4NgEtsK
RhZyShbVpa6Fxci5rP0GuZPGyPYRKDm5AN1Zzdn3iZ9+uDoNJJapWbtKeh4mVY5eopx7ibHLG0Yq
GQMHV+iV/cfL26MCP/gJaZIfUNKDaN9U9w+vv0xUVshxD7qYOHMOkFiCJVQTABfjohDSj0y4hLqX
WZbOfCCggIhDUhTuLiwcEr9KRAsQtvpaBnChcvZ1RP1//cASBcOxgMm7hIvwU3UWqZWR9wVIjZJO
Kza0hlPJjZHUpGdzPhw/Zqq21QJKxSwBjk34RWOO7lRfGA3+cflbrJYPDlJl/XWyEL4zpqfzyiLD
fPEkVUPXrBFUVxSiDIJETNd0zCxU4IpNkKqCK34nUXm4t+ts8YG8cWjUccpgKdkw6TSdej3YBj4E
IPF7gyXlV4OOsylaBxnIQUhePXlZlq4TqTy5eQqrZ3ea9SGn2wW3ThOoY4tjHkZPjA7I+9wTlE9g
agjELu8lcZudVadrR58WmRMsfvfOqjn5I6pASa0hkGz0iJ/dpF/p9tDg/wy8O6ARCxhQdqsZxsqX
P8a8gIVYGXGQ/Bo9n7tdZ9h9y97agUSSn8OKZsz4wGIUwWlcl3Z+iVAOokomWOt/4MZnA8ssLneM
uYF4viv3hsFsV0dn0TUUAu+1WIGs8f1zZ1PF5nBS/ItnxoXckFgzm4c/kbtzmWzLh+ItmVis/pg2
5Ge83Z026BRlgGqcebunA/ZqZnGPw8PYJX5NWUYMaxwT/BQGGkksw4OaNDJf4YyZQe7tJj8i/H4d
aALImNZZBM8pEcOKPKZ8OCdNIZqeFHvQydHzZJKoMsuKCWFF1Mx6Nl6Rhv7jT1hY24hGrpu+aQyy
27mbXegey7dOndvoWbvECtwXJoDxMKeTdzm4Meha5Vuxb3PqjGf4FSaWGKZaSgSpQuOsEyahMHr6
jFzRJaAjjJBbRHwyyitYIyVfJ+rCCBsKl9eLI9m9OpiUQvprQpfTQpXxjfRb5MiM6/WvcF+aJDtA
7lH8dTPynE58ZdFl5C7kRbBdPVauGGkRiWbGQoAuPzcf4zXtyftDan9CD6T2TNcns6U061uyBL4I
FONKf5Dih3mjWDsz3MMObUeXDYFDXUJ6ZO52Cq4Ja+wJr9irGR4w4d3F72S288XCyluBxzMdr9qt
/SQocNZx2WAkJBjIh+aEnZquOiHisYEnYWhO5MGN4dyrNkWURWn6IL1W8rrNz6mTsWab/D6Bce4x
nnwHd6Gak5P5WHRqMypL3qZzTU+A6BogwO/TjzVN00YmZrnXXAbRw7uQxt38t1NsuOnsldyfDDnQ
EKGfn5gXuXNB9yLSin8n4J4/mOKXSJ5Iuac9VW0BSkByk7nOtz5lMWmK+QtpFtIJbbARqtiUFDKK
6DdAGd6I42v7ei0okdNkzrHlvU8mpg/+qCEPAgETIrRAXBRvZzFN3KOaPInCS49qBnatJ2CKtMdZ
8taLCgvJdSoV1gDiJM1dgn75Y8bODdYK7fklJIfY7tRwvnkJRY2RpI2WsTlsrxFWkP8VQmbfDDzS
9s8izJEWCcq/WnY8JWsOtmAJrydco+l66HPlGmCrenI7PD6FVCsNEHySsQBEj8T4+tkFxhMaTzjM
AihrOxzBDmNG1a0iT/TItXNpuqhmUYy1BjccgE/ftQRJ0B8qcISjDlHxkhNhsOEMP0J6K3PL/xPw
bzZimdd+zOl/OUk/omtch9QUzpWk1GVTrkJZiZzb0aj9jlJ6KxIB2ROM2wN32eulS5+xv6SfapG0
MLaquhZWpcUmdc7iAs+KHE/tFNuW5UkYFK6JeAyBGCj2/NTcu3eqZ6U6iSyzhEiTFM4akm2os2Jw
qd7iKdi078llemfkaBXJupECi2RWTx7Lrz0+dSegKyz9bLRGdtLwmsPuu7m6PTQ1+1qPgpwqaZEm
dRjjDGAr3122xKTXf9utI838kOvijFwjmWMBiijM7kvI6Gotk62cS25ldY8KOmA8TnqFGRDsQ6Bp
mjx9qk9gQQkYQCVjt47AXR65JVluU7Bu3w8V3H9vkUheBVQ4W0KZKj0eYmVmdO8TUg0Y12307RVM
vstOn86NCmdrPshufvNwlu43xEdSVRFMqu00hymwfBbrdRQuKdwt5ABqgCVhLv0Bj5ezRdEQVFWr
ZQ5p94o6UKmlDNoTB+16QZIDqJ0n+t7ZuqPv5SFo1al8099nfEzn+lh7ujlLhhfBMoZGE8DrsT8E
xrluPGw1Vm/R08D21y6ou+laudbWy21soenD6xVh7FcRBWu52euwz0gHPLpHlV/L4IqK+s9VOZxb
smAq4TAGOmYGoaQwgM7VmJ2cOucIpow6WNtlhRk6whGNRwuf5innXHBX/L4rrbio2587sD76oUiK
Oy4ff24vgmTzr/aEquiWPxTrJJfrY/HTEXMJFyt5kr/KJPAq2dQ4Huu7fpk1mILY0zge05z1RC57
8usUafpIPYFYXn5ahyvFOm7LhW/AELJ5Sm19M/qBmOrUyN1CXrvieXpZ+5tVwH5MXCOSlQIGvrqm
7x/430sYUKHGIIFy2b8C0MR8ijrln+3nDQba96jgtGmKdlxJsVea3ilByAvPMeg6Wu4uVsP8kLQN
PnpMMYwvuESD1y/7GFTkQNCDgJXa8GCkSKFsEjhMyCRobuDLHnYm3sr2eR5cglbNJs1K/QuaKEhP
Snlv5TITpxZY1/O7SPTDubrU10cB/hUNToCnU9Hy9KYUCjacN/aYmauUJlYAuzitC/XXWmjbJqUp
oA/sFNKGErQ2rP6kVmYFNR25cBC8fZ00Ak3kinoe9kfrxJBsgt+dwMMU2RauKYItvxzDggoyvjgB
HaKc6qB1i/0sZo6eKwAuFors8WH5H+6ZZT2C5yDUKEYyCNRfRVG09Z/BW8wez5nhuQsbdnqLrwio
EYtK3PTv3Zk5/03H9lcioN4yuhFXNpYct8MsGx1Ea6IeOmndnfM0LstjsfH48/kkgIH64etzeUzu
+I8WX30qOGW09+OPEe16gidfDshFaFQ5a5gChDe1ug7+4Ubpzvp1b3A0McISroly92uBpm5Rh78C
LKyGdQLZ5+eLARyZVgd+Bm5+KKeKKI2DRRkJU7mDU8CcaDLTYFAIMTPMt32GUBA6agdJxjynknEH
hVhIQL8rK/lHU06ohq0XOqpuknOMMyIs1fkOXdJWzhUbmfvBbsFTld6lPvQNMMpAYDXc5tDhoMeq
SGppses3zHHjb/uFOVocMSPAQLMlIo/MbdnJSa3gTviJQ1pNmP18BEhHj7an4rQhFosRYX9F9wBW
wigp4ZxVcapqyujDzIBu9MV6dVoZ+KwMnGPpBTxDkLQIykA9jVdKTzkWUcGdB+4pv+9rP10crrXj
SMwGJE0We+V+OCB4hezOAsQ7tpkwRAjYPUmbRiuXDa4X8GwofAzC/CBIqKqbq/NnfULPmMfDw8pQ
eKC+xPe0b/jqAFB0ywHJdzoD+0Lmb0V2MKp48YOpnF0fFYHp0IW8BcrpU1eINDr9BZeLeA/OJtrQ
mq8S47jec/5v9N02dZc9ssFStoHXdDcvmQGwTrs1DnZ8ajW6M6uIrwWB12EPWJIYPZJXYGhQ7FtE
EC0KU8WeVZ3FjCo4rvAx9Qu+Lui6Xnm0opMTpEpceZC8okHSgIyDZX4s1Z1bnoyfq/hkyQ+3hl7U
6pQdDzez6Boh/j/+oVfb4eBsYAcbNZcdfWkVwKqKACw/B15XxPVKIgYd1sGqTLPYOCh0FvDEDR/e
9z/F3pef2LV3DgAg/wl1CcXQ+RVN5BQAB7uzS5OAKgXMhkQdNqzS81UN/WwqSy3JFpnrcx+q5KKi
Suz/Y06m7xj/ZVZ1d83sCcdDeDY19Cr7ARzfEJ7VEppucYh+zs9wVJAFUX0Xo0JhW7bGf00TAaNV
Qj0iPy8h0lOxdDwL6mwxwaKTDmph5hqEsDF7vd9bhHvPYzGBscJr/MSvhNTb8s0WJmPJ5q7+8GeQ
8/qS9VU+0iVKLeHHMBSebm4VHuGjYuA8WxRC/JBKev//M3VhvWjjYJCSU2i0NXEoBPu94FVwze5i
PBPi7vuO7PfytqqppGRq8nSGKrv32B04jBWqJCUnY9VDfoQb+1C6Jb3P2utGJY/zgffRXrvavmT8
61kFbCwWzz00lYv49qECe9Chf5z00NjyZ7Mh6fvDURs/T9ifsYWOtlCroDw22QvmaLMfCQ/hJ88C
eLV9CI90PxveAf3Ob7p35By6/1Xas7Pq1DtKSrfFIxG0I5Cr0EqYhKQYvYq143YwMM5pIOSC9Q5V
0r2ZONttv6yluGjIW2k7KqVmVi/yTEQCROn0NpETC7wW98/xHLtMvwqi0gyoWu12EOUx7Rr6i/9h
+0HkMyvcanclpukrj60K1Qf47ALG6jfRORrziDz7R6foCSKGdW9vzZvtxemCJd1u9CO9vLo5dcHY
K4QB2QKex60SJl1YDcmgIecKeTtjC4XLAHSIu91POlP4qTlKEB+2KtzgL8j91zV14gJstf5JiF1t
2HNk/Y7+3PFLZmNs7sqIZnNSYB8CP7OqOsvqnSmAcfP8LfBh6//4RllQ58cpKH+ZL3YL3f8I6vww
yxvG08Mnc92H8i/t6Egy7o9V7F8UjY7DOSyv4oPSUXBmriccDrjAtD8GjYGPu3oUsU3R9ODsutAA
I38571hIiw3nulumFfIk/XLrID/GHcK1J15E9DXVLPHi2C4r5Nvw3uHq0unPVhxANpzEW4LtmhFf
ZNIHnc4rtqJGPQ5hHN+bsCf8S9b6H6afFrcVALZ712B5soeZ+PHknQM/ahed5uJl7Onn3u4ksQEa
r7pGcscGutqm6KS1YNz+1TBkT/CzbKQrmTYOcx6RgcrmxZq0p1jAuatRucZet/wpUxjwg+0tljBQ
IX4D7E7Ojj3U6tCakRoD6AD8Zt2JI9umxkjcIPaPSe6jSuG1YbwZnCnaPWsxWH6VEvakOtmoOyNr
qv16gJClznN3FX/qufp6YLkK5X9TNUpUcoGwsOxb01oapqqoHzuqs9UhBCKHETqHm0UhBHn/3i3Z
XI6LIaoi4daT+0jBWJQUFiAQhXsd/I2Udr96ywuhG35HVwOtEKTQbEVD0aSkUBu2zfxKvBqYdcw+
hfYsL2T/18eZKZ4LwUYTyoIh/0LlZLIH3EqzT3BaQuyK3Qa183tfidA3Kzkl7sJeKuODelqrX/k7
cfPNi7TkjIZKP6+dOPUoxfqIH1XtNcu8XASpB8ux5Njx7cP9Zh+6/FrQqbx9gqpIqYVKUubH/8HJ
0ncj7TlsiPOwzeZAYKYy8T6KzscytVuU5dK9DHBT/xTHr2qkiLahi+lriT3bRoiKFSk9Faz+/BrQ
dOrEFFDTIHWn56JeFKbpQTKRB2TEJEIP48vzuYvGIoe9qN5uGSZQGHiDpxRKT4sqaZVe9mxberRs
wEsT9r5FNptSnlytZfsLqAW3vq5YLhQN949mPRdc4XdWeX0DEFhI+UQfy8e6SUf4YULObPApSXEi
hD3nd3+m6z6aqjH8zCDc51M7fxVcMdsEdG3Avb/rrT6B+KKJSPxRLek/LaW8fuzWzPf4ZNVHkOb6
3gJOHdzfyyfH8HULtH4Q08yd7qD0iWybxbfhiLZcEqgj9+khDHvHazYoYapAqomQEGelfl0IAxc1
tw40YjKNxMJ2UT2qjzNs5B+3ljbT7IoCHlB0t1Q8/MxazyO7iCxBs9kbx5jp22QxdxK8RPJS1eeq
6JgsNEavuz2Mwi/0mrHQHyr64yLDE2Grfri7URr5f5MO/meVWvxZF48ja9kfRBE4J1z7r8s9mdEm
hWFay0hBEOJ/5eFAyR+GIqWw3SGWsmGGk8mT560427DMiwheBePFs1i+Bh1OI/cW/8rEwjI6Nnfj
lUKl2+QtD9RDt8evksTvvnD9HegCaQ7qmstY/8YmYxRgS7CwijEjP8vdRIblcbnhsbyM4gd3RvCm
qhfxvJyXZ8jDpFu8wPJmep6YVaZKhkmI4F2QYqFcp/YrpHAeQR625IE0iaJETRycqRZV6egD+DqG
3FRbgL0ptpExkfKAYSUYbEz5iOLW+AG8IBsVSGB2nF/3Z0+f/L827JEd+DcO1OOxysJNvdp6LLpT
1JciD2Wfq0Ubkv6Ozsw4iIWwA70iks1prh6PLRNxMuuLJvDvTrlFu7fCz/icWq2D76LIOJDn0rTL
SeE8mTt+/FRXSQzF/jMclmq0nzG3xLCO6ydyFNkFkzOUv998r4qBQ1rbFtQoM49VVx/DaoFLhU/8
rTZgnX7dKT77JvS5mxeQloKdztSezfG58GoYXzcxVMAE6NnDt3TNeWDv/hdW8cx+45UjgvGP+eKU
4Fv7cYOTHsQPqayFwl2kk7Wqzg+boB26ckdDPFGgYYMjYwsdQMpTI7ClQsYxEOv3EDRp4oQszVWo
7vVzYDHvRqrOubehYpm53CjEldUvCYdA1b60u2rbRAgwASgmPTetcI5LF9doNDjwWtC80Vrd8qDA
c0HMgHvxEE3SyFf99fsDUZXf84Tuf6fPvideqycnpZ46hBaKmYQrvoHj7jmvfMLgxxBQakvf55LL
l0hD14A7z5ATzvgWsDQ9dfmbMiGUuTHfaWfSL/AfOy+mrRL7OPcq3IyDd9syVlYxWlOMZRW9qVuJ
T0O0iqaCKb/fMZ1LK4JT8Z/1slNc7EXpqvJlZIVaJtdCpB/XvtvEs9IyMHgUuTnErMFSuP/qZGmS
VSUtiBJGLvsqsUO2Y4oRXZpkH5+DgizS4F2s3rcR0W46KwbHUj/fRL0267wCwVLNqLoNU+GSIPIs
IHfy2GfGpy3YGrQ9DpD43O+XhSgFZRLqtVyEvqyOrYLbd7Ow42eTf3vaafSrDLu5lvCcC+pYKT23
f4/+/NZ1IQJWFsQSXnFS4t3iP87zOLOtxLGMBld0j0G+qYFNvTQZl62izCyW+Xgt4bracSLexj1i
n/o88wAzNhd4vn+wZCbzY4bK+gOFEcqWmChzb/Lnedsh17w43BzRHcbQDmseIugHuPnbbbobOmh9
Glf2kc/teNOPBxvvI01lunql3mIulOgFam+vIxfhKxozBc9lIOQzSDcnJiVQPlevVNsFzi/bFAFj
/r4VmWqnXwRNMLNqKig/NRe/lfZsfNm4+/n+K0Ak2Zu3/gGyj9jpVuFxEyGlahY3StRKHQJPnqhV
gKPH+4cdjaiDCGl9hHy+dRHRBKXEOqXOHeuoCwCvzVcDvWJvu41r6XEEeBY2iz8HUspY/dB4+524
pHdyNV92YhinviwKCVeaKrXmdnWBKVBPmpoamK8w6KRxU1Jc2kqJNcucpktKtIKCMelc58PhXBLW
Mp/GmurMEtjYNr6Yn6tdz9GvxEVeA5y2IADk43xOa1H42UMr9zD47YFB6J71iompHFOgkreOhYlj
oabkZTJJcSlq/EFcokXB5F4HpcqtGcuzzlaDZTM60RewczxJBkz0Jt5DuFpFEoKGESxz+apxa/QF
9gNcIc0Kl2XgsdJz4YUFZbALoAU3G8Xv+tyGAuf25wLUCfYAGuu41lf3RKQhDpbCJlefYK+YSIiX
A+pvQjrZrv4tl+nynj1Ntzgp/43kXCq1dJE3aBf3dBiQJ3TkMJWAE8+wI+DPUIZeTfZLtvrXd6ck
CsUpFVXKkalUjks1J7GKvQ/wZAbpdXv4w3fl0sHsUiFT5clucrEaVR9ZjTFMQOuRcGp0ef22SolX
6+q3OPNrPCXM2lkFExv7aImwe2no+9T/ilqgGK8A1mZNYobk4wk+g7Lbhc1tCszbrKVO6/7++iZa
4NFMH2IlHvVtS+uHFBBDGEHSK5TJv2iiDfK8858x+2NzwE/ujiOYMm7UCEbeiyRcCw9KHsJF3zZ9
VNZOazWQSZ/Ex78Ld6uhUkB2Fwt4Y62s2mpxt5UGnzIoWltGZajmW6IyfI/nhXDjjtUOCgmy0GX4
/zNsxyfPWkeJj09g0A5UEhF4Z8kja5rAzF28I4ymtcJF21+Egqe85Ylx0DbYwDWJKnnrNOQKksit
tGYOj+mqUlmx+EhfUYWorhLF6EgJd+D/WutChsUnPYVrZasZ8a7bpL/tj3+818iJBicPdOAydPWA
KBOgENhqAVbm3A2O9ihlR9YaETQN7joImcFHqi6dahrNKStsZoMP2vEQAfgi/UXwXcETEcMQ1q3D
wqEuy5WuKW18arjVpLS9GAXs2EkrzKGgMqYMyzn8nw3CvAHx5dOK6Hlcy/D9HoFnLZhIIc9vNnAV
4ZxhnG54SpZUsoIfg7FfpNZCIrQsVv/T8PDq3fnXH+XL7LoMC1WjvsOu1QiGHxWio2CuLIkHJRfh
cjRyPJewvEFQz7KUZyP4I1C4JYC7RzvEtS83vRxTgAOjXK6rXKP40HkxpPMm5rRYZxEb3dGRkkhe
wGgWR26IjU6eVlKjRAg3A2XDm5+ES0D9m0EkBeofveNG8k70DcSUo8qmSNnIdh+xgwOPbYS6B95x
F3f+/otYYtkm/hoxRiPFNs54kJ6usnHG8brJ9XuIIjMRzh+OZ75j1sRKGcaPxpyJbLkgQCmiMvZa
qu1HmwkSKvwEpM0jJM94+qqwm2juEBjNwF+QrIO/wIWONym3NBR2V67qYl/DhtoOw0ADWeA70HxY
3PRFt9X+z0R/wv8qbzaHe8cHbJiHhTkW3WsFBC2d1r2q1yKShAfWTfBoTw21S0re8HBW+9OeD9ki
wEa7Tfg7XwUSwr+D043Gzokw63et3o1HsNxgU9gAeRFHrOgD47F4sCrXO2AhbgRNtdD62iFDwU8m
uDVgBiub0xVFgzxwRzHatKfw5Mw5yPACAtt/eGcQgySA3Lnggb9lu7in1qSCSFyfdCE6+rmZevu1
z1r8h28o6aj1wVwrscCl34vemqNJr83JVdAgzE3gzzq9uyuQl4rmb/PrQE1X21Ig3Cpftq7JEIM5
U+g62Tqy8ev9toBueUXqXCX76Q4QIljGmtoDvdmdiUZKGeQxaFJUnk6xWnNxa8QetptQOIu1LdRc
gvPaZLdzl0fS3IzaiG/loptXz3lIO5OXku6GYlewyzOc7SodS5r0AdaASuRc4dZlG2rDMzwGOxSI
1Htb3QoFUMTOoi6+/dntr8Sg29S4jvnroAAktMsoUNj10FzaxtEL9J0GVXH//mieyuP9vXtWYT24
WzWyaauKHQcc+RGVFMsuu7qHyjKdSAQdLXf0N6tGhE1kyDczLphfcWzkaSRrF2KRZj9svk2q+7+i
yVOUZYuUdpyL5rZY0pmkceDovsnNWcnmZHBdRCajMbBByyhDgBrtaRngfpNDaEG5RJ4NT+8wNr9F
3tUgPoA+3n5Nv9qGsvL9byEWOwYJ8iKehv5h5igqN9FA39Rod+FQSV4/gac2ynejg1b1OwU+kYuM
NIjNcsFTdRlzq+vKGByp+bsl5CoqbkkqGluBhWm4mXyVjx3tAKZyN5OogWrg1G4K+sdV8JV1I7gK
y/SJgoy0cgYwJEV7/GV28+8KXOQBm2miC0RJCG5eV6i6mtbsJf5S3w4koklx/l/VrjWvxPAgnXpM
PjoT0YKExh7GHd3ZlGE5IjWm+sd95YG8XVAPKRscAOec7LPRGCsSdCE6xj91GkM5GqZ5m9ud9D2V
7hgYrVDuH1qcIKihXIlY98ksCq2Ic/FKtvPLI1876ujCyTsO2rU5uuNddUxdMF/us1wL0E5JEdi6
KKZFPHtkB+Y5r1NIxhSUgACtzo9jELr0lZqDtcuVGpmUZ8EvQYCj5wecP9iG1DUaFSe9AO5B6Lhl
XJwXT9gCQ3ZDU+/mUxC4ytK6ZJ5apgIuL1MTfcJMIRkZa2oyE9Qaabsb5/+qEqz5TySzdFhqpq8L
6IgwY1wh/rP4Qxh7HGIFyEp31o8VRVqikZ8fADHqxgfoBbqIdwaclTsbA++VnNfgpOh+7dQg9883
EYGNEBB8I4I6mcBypLFqtB+YL0s7RNept1er6EAuKfRyxTJUjplXydMGF9/JQUTdrvht9HSOftj4
dfQRYUAkIo2oUXsoFGIL3pn1WJbJ9vkmTt8y5rJx+r0nzHWm7XbDSUay3s9ohfgD77RYMsCdNBT3
TsXrrTss67ur1hc+AmpWQ+cOq7L+d6J8E0dMmtuBjTl0sIhndJCXpptf4apdA3Sf0M/8kBNx3WR9
ctjbTXLAbQ0fodYVNlqJsZOXWq5Djk+VuCDex+/KsTJ6HZCprrjeB3AJyf2XAT6O05/5oUuEulvY
1o3cfDV0dg6li+CQFGpeUxn6go+aMYMLYhaErzRzsT//yzJ38DNDWK1OHkm4qhxVSFalP/geGU6w
cNNG4TpDNe0gfd58f93jO7naBGG9xId4n42WmqhdjjyIoROE07bfMSV4MGNardWgG3KxnM2ltumF
20PiKEn50rAns+fSyrXrLJNlqhW7HpeHPh4R2dzkpymbFuA3IIz9y2eJMcsSrqGkmkfdbRld0JNY
J6BEYGp2pjsFDibxLq+xx/4AANWfnAuYr+q/NA361wodaYa77Ar4h81Gz32H4pgIDdAH3vWj+IpC
vAmKcEy0mtTNeUU6qAnz5pUDdWx6BVrpC1JQws7ZOWmKxA71OHQp9UlkxqB5wdrHOW7TV3b1444m
G2TB5k1QXO05IpRfARAqdBi5TjeeYYlD+4MXoM8rlJTJ2rUUUjhqOJVlL6N1ahMm7rvlH5WGkKZt
l45/0XmP57nQrzWWIzeybT5jAOjKCXEHC5lMMcXdUVUag1ucVRkpzhC4Mbmlq1uvd9Cba6TTCZdX
FYRgW/BX9sJsBDwkFqiaO9hSjTOxUtXpp0PjKwE8ehBROWO75rPPzjG9arKGU0E9oy45onJqLRnh
JZ9dVevrTJxBmLQRvsw/Ed11EmRI+NaF/o44yDjWSR/xEBECfVJzpc/psRcaRD8HSga/RYAPbztF
foFDed2xrURwD/s27ySplGrI9e1OZZUyhzVvfnVIZPj5P/2zCBvWXMpzXj2wljed3pIuecmfbPtw
I8xxrTUG7jPyXC2lCwH8CzV1phvH/EDk4o3mDzVgkZsjALuhIMM+NkMl3MDd+MuEijR/dniPmlcm
7YFgnfNr8jtNTzt9TlT0wDvfKRnd0vfotyEXoToPkGYEHcdViYefQHuKCLnd9DoyaSXDJki8aI1S
qNS4ocmGeyKpwfqbg5FgpYPAoB7YIryOXsUxaJEmP/oeErqx1V8lwUDI9o1tbJesf4i1n3DZr9MN
zfVoKyKOTwflc1WRWp5G8T8BlvPmMbB5HV6RxI37RPVUkwlNbi9hmiHFz7mfLM9PkLNfYMFY0HWr
ECS2V7Ecp7gbupytISRGu8JMe9YVzKt9UypM0pZni/P7WICtN81sGU2tSlRRJ2+BMT4qnBbj2rFJ
pggrqFMAEzUYDUWecULzmuWSiXmwbrUryrhFDa1ov05WGXqNhrX39VDCsjSQotCAkf0P6jhsWXwN
2fTz7zvDk7W+Z8f+S8k+WvlBg+R8MH1/1SknTtAr/m/ZsdWC4TKR0th0NCzrJrOxgk5bakw4Q2JG
L0WnKWQZh0774MO5/uxxRvmXWu0VhsvIaHx7JBRwYRHr7wS/jAJinbX3SSOuorddm7GjVezegtEN
IgMcE5TqgjHP7PXXeSazybE+HiWFp/tUdlBaa+H8GxXwlbnwQW6UHhsXVPwm35EVq7d0PGrkW9v+
28KFxkqqw9FfTXcP7BagShag4SFHi2SkJurU00iP5xo7LVAWIz5wkNqfmZdhPCYIEsMrYgIrCqwT
dgoA+CD1471hlpIhh2Z53FAnkc9XaqsngnrCPy7Yh+HiKjxcOU6zhiGgo6D3yO3xYnSoOCbj+58g
+e0/MkR00BZhCVlLrHu7fDHEwOvw4rYQBmwkwMGasxXfA+daslP24Xr0UMcoyjwPQaWrX8Td1Bsq
X/JL6K4jdtME6SeqzAhAsJSzEU2HfYoJnLyhY0GdczyG9SWS8+GaoqGIXzJhcdf+Euy9VhMvRsYS
oLOU/CE3v8bxLcKJaeCalEV6v3Tum3QaTG64Pk7l0JhqGLOvyFenDfMqzsTc1Fg1EMCs6/Uorcw9
Iw/F1g/7/v2YL1T7xo3lDpniTAKg2uTbwTXvmMRURG7dhxHmn7LpMRUHDqzh3OaeffQCdC7wqwN/
F5xuorR7lrRr9MhCLV1ojDowKM7/UgBNSIvJtLxVyMrU3gjRw0C2oa2YjEzQ//f4RgwSEfKkIagk
rTWFike8QkTKaa3A4uzlhiiS2ZIY7JwymUdQUfOGii/Www28F1bWpsMq6pUw5BGbGlYAD4bEkngk
PAHbfjT41KxztvTX9q5qT2UEbjOCkrG6kfmc0byG+tq/zG7KgHqt8ucPz+ATiBFv++dR8AC+wQVu
s5BE0cLTTU6qPNx9xxMMWt7wG2qqy1OM+2VQ1G/d2WgRD83VxNSGQZj3w/hd36yYPLDSMG7NRO7O
jTIkwv2OaEYQij7kBgay1XtyD6i64GGJ9yZtf+OCUGRPYOdKmJcmoW6Bz3cFZwyJ3+HBexqv0FrA
LcN7YJyi7mkQ11unCvStzM15SuqUSu+QQAloHOYwM1LyqEfI/Bj4VQH5wUkY6cwfGrxw5MIrSIHi
gxijjYldfpdP/G+dk2uWhyAucjq4ThfOPtFqY33wXt0kEs6B1kBRa4ILeL2Sq44FiQA1sDKjeCp1
vGmuNknGNhmPZVkrivCQdqFJxgnu5GtkSHIJcy4ASrfZgrAEoXgmF1MJBjczL8NX+EaorzYRwF4x
h5rNQz/5+P4+pGXQJtkGWPhVLIZPPMGypxZgDa2Sn4dZ7PuZDUQIJC1/CWNJCQPO8YarDTksGmip
NOJK58KlcO7w7rRzFkGkVqLLm4lnzmF7jYnglAUtR06U/eMZHaWrPA4NpUCqKj+9ZU/NDSXiBRRP
368sG6vgq8yga0ZOXeWxJX3Ov/NjFQcquYmduc6Jydjk/RzFQW+0B47BFZ6+tp13h2c+X5xbg/iS
mcURMFPhNjSJY2aYaHjKwdirFgn6TZkEEM4NTDcg5PaMu7tRMNTpI3zfvEtmRiB9H+DJtRgOXT4T
XOXiVE14VAHv1tw3FsoiusL+YFda/hDCNK5cMIMSGW5ceSJR3AMJVS40XJXQsV0Uws6HlWmhSXOO
JSVF0CaStDE7XhW+PIZ+c2kKoQc1Hitm6/gdxy5uAsbgp9A0pqS845ZIgsFKbHBVvD9Yr06mT19W
VJhs/CKVDeF8j50lSO0Wde8wR8i7eKQ/t72xp4y7sWQty6On31swI8eNkFAtXW9Ez9N8i1VO4A8Q
i961RiuBDYlROf6nAXXN2auLOP7oNj8OhhddTCB/lzO+yOSEPio+UHq+wDkz66tLuHhbaf8WNoc6
nVvoLdoHQSj5yWxezM02UvtvciE65T5FzbB9ncZudZc0sdFSyr0al5tm0Uk5H8VFkaJHLjgxZ15P
ooXffSkDCNkX4suid/egOjPlhqaDiYQUPF1XGoyQduBckNus0YgTsT9iKB9tFulwdQrHUdUzXKbw
xKJXvGVe0kYx/6a9gmd0daJiUnTYURrw1M291ChfWdlaeH76d/qlW2MrjADKvFS5oGprxTtKrMn2
j+Sf98AhJ/+Xka+vIRsrHsMNkeM9Y83y71M/ZsThqaAsrUPIkBwmr05wtHnzfjfyeVynsvLy+RtD
A0m2bCV0g4QeNLIt/zObxKPr6GuOxaZ0FpRUhGLYKRlEdCh6NKLNkL35C/73X1RvGv7Xi1DCv33G
bjMfFloQFcGFbtDABXZqoW+HQ+teZe7iRTc6Q3f+aTmsZCTT3CmDUF9ovXRZnzr/HheMAjcYx78q
FL8XoRCSqLgBVCd9lTne4ALFDPs8lGCFms7xpYu0K4IVRBCroGiFMMrV1qI4xqPlhmgweLXX2UwJ
xkn9TvQ2vZQNsuDQcLJRQWoRk/EWS7G0jzJ9IseOLLlZrsZEtwGl3SyDj9I9GQFN40XtupKdxP7s
BIXe/aiWT4+Bsfb7mqVLRviw1j/TF4arTHNMHTZ1Qhd2hr8tfOy4EvHMeQZ9lhptNBmzoV/u3Sc0
e4Hmeg5es+0cZmUmji4orMVlG+oEYK32I1rUf67Lf+LcEYJrITRrW4nD2TYIoSlRc0ClttpzN6Mr
ZmOPdXfgCebixzwdYHkafMpxtBRaVOShVsmL5De0UKW4yF+BQLEt2yIm98uGjmWDSISIeAhGZZhL
kCeY3Mw8sriviTV4BNRrYP9gFDLWU1on0xwEtRap2ufOo1L1aKrfnyqKnazqf0YgLdnFhk1jpvmT
GWE0Mccy/f+OkZWsofq8IPsjzoiS8E9RPAbt0g7wvxuBwS7U5gaDiONewWJDtWzB0ppCaVZxq7tR
rIsFDfzByZ+IP3HRGv+71Q+qM3sLnbfAqPwncZPHuWgAxJ+257sSjkVkAjdDPIATqB9MirTtcMeJ
4nU6bJeVda09ee1du/vJirUAgSOGZo6scy3lm1yCODxOIhFleJnoTRSkndEyIDFVnKEJb3n3YQeI
pBrkksfSf+BwBcV9C4Ge3QYT+1HEWUkBalOU/XoiVhdriUMpo0jZgOGYYJVaaW/7pKSOir5QD9Rk
xaRUWwD20xIqtzkXLk7tSX6aSIoePHyv7rM3vKGT5jgULrNYukbubzYs71t0m6vdqzdAvaxsnWuQ
JG2rSbZvxV8XoCG2gS4AC7uNMe7YdxXcF6xkarVAmCHxyMRn903NOyN9nWRJ7vPrfY0HXUojHjsZ
ryuCcOl8g67ipkQ59wZnIzH5eb4ps/8cMFcjmS2E71RhHShH6rd873VokL6uQ5iawztN8I18kphp
w5Jq0GKt8z6gxP7Mw8TZpQuzTBOXXhd57r2Wg2Qv1Rct0Xa1QzgzR+m5YRu3FkUIY31TyonMu2ot
iCpKmgXou9l2daZhqzmsrS4YjyX4drarBLVuSfxi8F+x2EpoRrg0ifkWKNcVbi5Kmb9EHb+1eEN2
hawdDEJAIffZ/oJlvFjdbZ7ouU9BlKFuECcfscl6kDvduN7rSErF4EzpDQBvsRUXc5c+Ycq7CoF+
WxnmWuYLO9p9Lq/q3ge/1JjQNQtmN0Z6azNsUZpu8TMuM7VKLg8r77ZFM48tetQipK6VQgMzGEYo
g+2ZwJ3lOxa0tbp0nC+yjvWXp38goJTu8zHDLZVw3byeG79mCpCp5Uai1caQegiRxjxqzF0lATwN
ZwYIQtX0lXfD3krbs4ASDogoWk9+bIdLZr0DRyLJSl52gCwySvfgt5Hl0xO8TXedwo24Jv5OGuoK
KAXAFLs2SVaDBeuRMYezpnfHTKIQTet9n+93p9XQRw8igXRcOLt/oF2S4LEIsg5basam2CXXgA9H
+VtfNiSxA0FhhZ3OuzDmp2qYHsHrRq9w8wgST89HMWIZigJFr9uhMQTpAGiD7ZiPNWvy+Bh7FS5h
peQjEyn5m9KzkMZ5nO4qFIqU2GnzgyusoqCBEXntflm57v2AQBgOSG3CmSGxytwsUpsLqRsDIqj3
T+16v7ZBCpC3AwSe5uR4a3s/YQXsm0FVzdJ+P0283ChsilKgodbFEC7B389VZ3iMCX0NtJfBdfJP
ZUIaP3v0TWSrDlKob44CK9VJ2CHVkTdQlWLKLvAKOQAFdfFh6SbqLbsO+5l9YgZzVM1qKXJ8fpLg
zPyD452RBUrUVIAUxVGuwm0+OfmiYMG/KOxFsqcAkXFOzQFGW6x0vdilLVtc4MYkPwwN5XKktn+I
LGATVGPntFx+9qx5nUXlSjfU4O40Sh//QfJBEYAgcFrCIq74IZ1qiY7yC7elyj3CyLVWM6tT+/oD
WjnjpByl/DlcOAkMptURgf7yd1ynmrwm4pN5iaphaqVoQuhbjiF6lMXTD3R0v7JprvnfMTi0BdJA
K94VH/20ELBVubTcnjRQ/yb3f2x17EHrYyDIqleTxwTR2Bx89QoUVOrFZU4cyAA09A1O2RIC25rV
huYOqMik8iMtdgraakmVYzlChDFGhib4vvHf3DHLrFs6OoqhEwmlh/FNUe3d6XC7NcMB3shFB9He
9bFQY4PBKGvnYQnswOxd1DEcnbgqaRIaVT/qP0rfgch0q9PubphZhzCjQB/BqZ8zGI5duke1JWfu
+xhvKUDKugCt0guRv1JopjlUSpXVewGJ1WKdlpR+jQXjoY2TQUBBPDYRuN2eObfAGLuRJ/rW5Vjw
0czA2aK8odh/PJ85GOqzK0GD9cRXOj8GLEASUcB+KUKG3fSn8/bPQYlenLVsTg309rQYWr+LrJx9
iOo5P0CjARuCNy4nO/Br3VIukgJG0wt2WGaPmTd3KVUYRjbG59Eyh7Y5x/XpiT4hZvvD7N8+Kcz7
xlZclov3NbnA/Tx2hkoeqMGwT3tx86dky/f7tSLdNXUrCpgmLn4ILwTk8SRx9CmCT/xNREZ0+Lde
WoGu8EqHSZFYutC/y+s+jfoL49ULDBDOYoAqw3Y61q55PHE7c+e75xU3mv8errtoBfooji7Wuhay
KNqlpFK9kqaBHJ8ljt05gNzfSEOrSWNTp82AFQx58URm3s07sgXGFSs+UVxdrNF3fMPGxiVOu1ir
aECyNvxR2ixRdgGE3wiXV0k5daPewZbnPhKh6Q8XIsns2sDdlI51qMEuexCW5HL0HAWjO0HwvgOR
frX78ApCKd5K8uusE8hKIMD7ywmbqQ5azYshkPLQ8S/hfr+DizXwmPTVV+lTtX4FLnNj0NHtDKZ4
MQOLCVdHt9J+RXQFZwFN6UwC9Kma8G+S1jd6W7nI5BRpi5E0GNcSoRNBmOr1uOSIhw6mAU4aFvL0
VsrNtWA+ku9drQy39qbRFEJqc1G3ZSNJNeoXdAki2Cc4unjghbokRudFeqdR0+5r9BJuEyal5WgD
WBKahU15uj1dQwT+hlxbZ8GRladG8jXy+EUC9hu0On/sHKetFj5WmCs0QWqZzgKJr0SYh1d+WoxL
HhfINvaRUp+jeL8m9DVPrSRLnrsh3Rs6VjRwgYe1/FjVTHJUk+VExUR9u6OX9SjI4qZ66mBb9xVL
o6Wuzz530RZpYYzr2NBXnXyVuoy48nEPaZ5a7D906vEZhF00IMsxNToSo1tihpwQcUiAru+zJddN
qA3rzRm87d45z0S8W3wK7YGG/6aB9jd+Tp/ybn3CAXNzDz36OLhuBD/dPjfh1abHGpJQ8gupkwsN
cmxUhHeCbXCs//Cc3cJSwEn5Og0FnPsOZSRkDea3xDRnOcXC7hnaeMlyH7MyiETjocPGVlaeFcC6
tN7X3IQy7xFc05HmNDkocM/U8npAAsdU8V2ZncNTOGESiZ02oGPw84v4WLTrs3LT8VDpKrNdGod5
9UmVly+HMj2XKRTkuO9mMU9Nus/o4ArxGsrrnyR3+8UwP/zy6yfSFL+lIjWpahCoLkhzXtYrksEc
LmsZXMBycUk0DNu6N3Sx/Thet0msS4JYgF5ZDqQkY0ZlpFgrjtPqhjmSIWvBuKcHYf9T6AvrpCG9
WFTIpUcc23rE3p4WSRil60Z5Z3t5TeWhkqWD923VtCvsv56Wn/ihTAZPy3ZANAJxdcBRXIl86+Yt
vhQKr7k2BFHsRUBK7gM1DlF529/1SAivU2ZLTnXExVX/rZ+qlIRhPwcn1xkAx5WC7YRYfF1A+VOE
aZ0NPgf9IekPwm211UbSW5FE82+OYcF0HO3OrDzGECpKIpR+LHN2LdT5A7k3QYN3KxiiuchuzmKx
fw2EgMzJI/GSey1cPGGt2ZMa8A7faAIp36NLHuGvSz17eNyakok/UtJt/nAjZS42CBEi7BHDZB7O
yh5ioD+rCYyjycPZCUASTv/r7+Ucc4IB0ioSaVF7yTPhJdfby2a2CJKPSN558s2I9GK+oHJiT8rK
3GrC36v5K8cZwVLvSvlpNEpQDsDfQYhxVni6UIgt5SBjnOUgOLsFYjUXKl1srmHmiXUJNuezN7qF
qDNAjsm6JzirluIgKNgtsuGttaEknnZ0yeCKcwgNarJ1u+vAmprGafEbXjKdp+zZby5licq6MYVt
0rNMQI9zIox4z25wrlRgFYg5KKTV81Q2erHZK3bvWafu5niwsZsYyifjRwVC7ObuAfkDdWHh/OPI
u5T15NDz1ECZ6uNXJWPqvanz6pUrwVLZbsf6LDhnWJBPt5AkqPnx7n/9ebIMuuGD7jGWZyDRPMg9
nnu+ypswJ10OVMG2OmgHuj8meb5Uv3xv4QIrEdUoI//kCFve4K+emSZdEJTzR0UB17iw9oVeVaMk
PZQAPqqgrS7s0NEmP6Am/dJ/EP/ncUlSXjZpn/VyGjKJ5+VSVm6wI+Yu3iFU6lS7DOyYDPHZmSrp
lqw3Yv9MMHYLw/wXZSrA5UjL8yTG5XyaNei8I9UPf4Tl75ycLo4HX3IgJVJPQFeoMi0Hw0p5dkZL
EiArPGuQejkC2SwPVcHi5BqDURiA6wKWAgn7p7JyUq+NUrfS2hFKZxjpTY6HpYLt+Ll4i28jYbvO
BrDFA3QbO2vVXngvGg+JfJX2i1dKJp1vBcgS0tHyZ+/d27yFIg+QuVHWbCJeo81WhFXPsg4YyvC2
UM5PxVwH9AAYp+ba+wWNOcMiEKBuGOMPod9TAUr6X97+71MffkVOkhD+msTae22TYoJgKRBjHjfz
rSbBT/rukPyCAlD7iRSYJq4/F8rL2S4utkB3n7tDXixY/XziPYju2wSeHZ5dGrDPxT81KK0Dt0/K
1r5g9ORekMDAEucfvMpU4Mq5YJX3lvoSDDrEfpfu3HVcce7NmgK/kWXtPl45puTwKx3RPOwqdjrY
zSlTd7gEb47hBSXmGj7yM62gKPpO5kbqENazhth1q9XDzTiANTVqNlafygkymStyO89GWfNiaYLh
s09N6fFg2UA8rnjx+scrgLx9xGdqIpDpW4I5aijSpgqGORL4MHh/FPvUUtQXdw9/lIjg3dr5Qenu
bWSHdZ2zbbc7zclnHuSRutWe/cGiP1FO6u8x116bH2ptRi0QJG+TfGqzd8q6/6cTgpHav72TasN8
tvelL9I3qGRkOJaZYx8rJkcZHWD05C93VWBfuXNwlWgv0HUgJVbeNONG+WfVGGZ8xVlWu/6Ug0Gg
GNY+SROjcZE87BSvkfBLeyn+CkwZVs310dLPUr4An1cbfW10nQocZ+VhP/j90GiRHFbuyQ0P4rjn
OQRhVexUgNbOmVpUtJB5xw8bt3ObxCMXco+Be/ZWQILh2W4RdEDaKsG0zehibHNyhfrW019krIcl
LN2kSC1t7unGmcwVfJItmm+kPSgR0ljoKt5HaREh2wuS+IO18yt9WXJD9aFsxo3DnLJnSZCwgpcX
23zz1QBMrvQGXWIURqPqrCsoGPF9zfrkT+5SOfWGm1K4YT8+4sDRViZnD4f7dEfjCsedLGQXlzj2
TkiTRHoTLA7/O2ausPIzGVIYb5+k/Y59dHNSy/F/tcyJTJYS51Y9WnFGptrPCkSFJDFRyxnQgeqd
DuT0Gqq+b59pwVDmSSBeS7Coc2xTHax78hZGIcM+Qnj1hAGS0+Ve58DvVlRCPd+fBW1f7lQFbq2Z
guHRWRfIBGSg2qz46nDBQf/fEQbws47kis4j3XYmO/gO0qc9d5+URTbxi5qi9GdUh4gZcIDC43OE
LrNb65BJUt0lUkN1b5iPeTB8urUQYpjY73a5EicjnWjBmrz5N3nrDaAYZ3GLkPHH0dvC33g9halv
LrpRd6mdkB1TBx4zrx455f7WcSyyMRX71AFVSk5NgjCnXj4TrEjn1aQMzMmNUGROG9lqAEqPa4PP
5K3CehY/3fwKxFrBk6hI1eAu4Irk+PcwLMt3/qHGrqbH7icS+P+1CTTgw8Pr7NhcZPe5MDKXOvbm
SIfcjw5+/ogAOkZeuyzWag7bfucNVZZt1DBV+0x9kFWdF+qKW3daaY1cFbXKNYwpBJZCWSJyhLr5
mt4RbIm+wgHdm3vBB5bdfzhjjFb9LhJGnA/FpjnBjF/bMXkw5b3qlrUT+xGtKZ4CnXoY8ISxZDkX
nMhfMEgPKzgbr6hYWMR2/Z4k01S89JhcIjGaSZVP6QA3tRdTDQdAECohaT8/QAz0a0el2OBh8rbx
PFiIQZ4pnSaig1ZH4OO4+BttllRtLla2M+SIQ7nQ7vCYpeQiVHbtRRxMA85KqPZaYQj5jYnrNsh8
6bn72OUIjN35Fu1A35/Bijj91ypOk2LNE9lodLr3ry2p4VmcdvkAoaQpIv9l6AjjTXegDXkpkgtv
1UAs3Z8k1Gcgj2fWEPswN6v1okAi+ranZ5F9YUpFZ6uLu0N9hxFthfTm1B9yoQ77VrVHrGd1oBzp
N1e/NUNU8n8EhKeDWggFHvKA6b04EwgksNkmH/X+tDDvvKPnEUF21letMZrsGv28uEQAfbnIFsuJ
Hqbkq05m10hG4ToFV8l0t287y2SmFEHmLIo1ns8LDEi+uIiPri82Kt0P9vRebTzrUT1VaIv6URLB
mgDi/KwnHYrd0BlYRxCMamJPk965Cz0qkQ+AvPFxzjDZ+U8eEjOH56lT3Du6Q6zuopeA+6WxrtHh
1DeS42hJZ7vYF/GeTXf/DcO3CY5NFd/UNLe10QoppujxNqIK+88izxIPQhYbqMSXrffMJe56JHsP
8UH/QFRH0xAwkUUs25DQsejeh1i4JDLcFG9o+mh13+k4bZPzvWvDXZYMM+kN3pdShTxwKpgv6dCM
A3cJDVPmKoq4YrsZ1IoEmWVb5utl54Sof6DpJEfx5GOZwDn29G7IyxVKYRs6GcqOorGWekyB+czC
X8VC8fIi/BJE3WbjXUlmlFgvWyE1nRoM8yMmNH/wjr2kHAxHnfM2FNtSD3HmKhaLeAxlIN/UAb0/
T11cKeyhOaytf8CbzDfnacpTA9Kepa8H/GuaGSs/pCTLOA7t3o14ckUpVZ2WA1tk6Do9EYNXc6Fk
tjTBt0cF0ePu8ffNxKMk7XVYuehNZpPIdztLfRMsPLpCMXnwa64pS5gA73l+UoV10FHM7gvZiPka
mIFCReqxlS+mqaVuZbdbPxX9dzcZX+W3OEQ3bHNb3VUnrXc0td+LZ2yXCU9YT69Hff2bVerZIxmE
cg9JkJSg/lYLViaX2nGK06qVs0+QLG+C6gsNHKEmAdrBD01sbDuvU5YxLevfSh2BPohMEbzdt2yW
uJ/dukbP+LuZ1a+ov/AIs0o5jOzIyHturCx2dKNlWbJfvxSNV4B1jEMiiHBKoJxQmbBNvBQv1mSc
nCymS51jeq6TJuEvPoKf/6r9NmlTDd9jHgyaNUahaO0bMlZg3FwUvr85en8ZW+FiAfnnZD5UIDNs
bXsDvrZxYR4otBE5RtWOPu99oTwSlRkbzl0JlxMWLqESuZvQ24rP2FoaRJgXf46XDCwEAK40kSer
ejNJKqtBvzxQjXNyuNB+hx5i+ZhJy23crEYsUyYKG7Bm1gQYghZ94YaeLDFBjTPeKyCqeLgLaYnC
YHg4OpYYZxK+kGFRZ1k3fmaBTOESfZMkiHSUrA2+5loJEMQL+w0OcbWFbTsCAd4jaW59yOzOvtih
AQXw3Xi6b/zcmutGqYfU++Auz0eGxz0FAPZeNid/ZnOyPFQufPxBblr6t+fnEAYIApgnAveiLzE5
dndbfnGt6Mzl/v20VchukcEwqLv1pYRncB00K5aXz7av6l7mhgEqG2ELUjtLo8YNjrao30n+9hG7
TPoC5JM1jXUmCpDkVaSpYxI+vGAYjeQIgikEYcIxc4AbQXal5JYfiiFy1pu0tMDURvmpkCNhe1Ci
SOehXUddYq5Uo5qNngkGCvAi6PKBPI56R8xybiMw4n33V0psadszB6dINv27Garxw6DhVlk7J4cI
hj6vvTS9wDgrKWdbLV1khu2jcu6ht86fWr8nfurCLxL1PDGQz60efaffxqO7i3uMSk0lMS99eCVa
LGck74xliYSwz0DjbG3j84TAtJO4Z7CvP5y55Xi91m6KSq8rCPvsUT/IEXSsObBs2Xa0FhuAqhOM
2lSPFF01u7SPKG5YzCUUCxOdclpk6sbsPzPLwhhxhUDfs2b3D5cPs5eetcp+ay7/fDZK8Jyo7BmZ
wliXGqJa9WO2dz7jdP5xB7LcIyXeyrfv9SGKk+4RpEkAeXdk0mDzK5md6E0G/gNtb7XuoNsM3oOm
rBQ2USiIsS2GkIPZIKQZuP8DfJ719dk44QGS+e27bSzHIcRabtD/E/HLH5uZtsTkbQEwUk0NDYM2
3v7gHnBkejnXeJiuka74EBLnozN4dnvI4Ur1lB1bO5a3+86mdhX57iR0wQEnVznTcqviCvbyvAML
YDWjXNceuublLcPGDWI2W2W5HKD+D10jxz8t2A9mILfWJ53EX4tVWbKxVeDOWaiUySOI81fVdqMq
CW9bWssAa0nyw7aUn3RsQ0sD7miwUSUWmENAwxY2UCBE2AmwEjG4oCic4hXu+rBrsPos+URoT87q
U/R+OKI70tzX9WpNWlzuP72J7GGX4T07aiqRhZdAzlZvT4ZEsXgj0W1YDiCNXYssbHDvnWuHGEpL
toYmV+auOu6OASlS0QkT83dSz5xVLfrzLNoSUAucn0Nr6m/Y5+2nlgp063qltQ5XjVz08tnGhuLx
jMZRCTOZHV+o+kRwVcRxTm5iCynqAgxjwUgNYe8q4S5ufhk2fHlB4ZoaTYhC9bWG1pTI4pzeMuqk
l+R/dLpqFIYhXP9G4LfPb9Ri7v98xCBiihwQQJhCl48RAKICFa5wDrGJVfrm1Ra/9i1QELw4/55k
M8Ixbe0h5QsgXrZWC4BGTawYPkCVRkHJXflLR9nWlg2nViubXRcYNXy7GuWFrgdZXI47AiYq8YI9
sRhEH1iY2xT7wjtNJD6YlN5kxvhf76ZFqAjUwsiLLf1bAldeD3/SIClmOTYcYx/o3DsE5jC97AUw
TxBNyXZpcrfozk+oAMjpklPCHUJ5ZpeYgDqmC4zv9yZiXSA1wnQF9LZUD/jLVQyo67mS+hVda7cm
JLhul8oFNr7uv5dHcr+EJKdX68zhLdqa4Psru6NHTbFl0ARI9FZRkLm9Qs3RfP0rc6kdvxQgKGoa
lDHa96W5Oiq6Uh/qP/NuP6WwppW1jtyS0eJ7Sl7Lgoeg6GUyAU0plvHEagjikMw0bGCuWEKb8pAG
8HvUVewsczqUyeFAn55ib1RvFxO7ukN30/ccOCi+bPGd+GX87FN+xHU+cejZCsGK/VuRwI1oF3r+
DpyfTl3RzwFj6f4gf0yv/xPcxvziTrQz+AYOTDKyMs++nLbbqzDJhEn3Rh3G4iFRYlg0Rln2gzr0
I7V+16Wko0rq16EVvCFEDBT1b6ogsJ+zLMhEqY3nFDILqIrWXu4bn7bYDr7gPXvuCI1hX5VRQfTf
lBpAf179LKz2Kp+enWxn6VI4N7Jw4opjS3xC4+/mDSJNPiKEuO/TqSzBBYtUxxngniKKG9QKC804
AFjldDyIHrAEOoDxIV2UDwrIZUP3Ny9hB4rF4pT2VawV4gFWtRplVZO4Sl6WF+svg9J7LxqyczPk
06FTzy09Y/b3/c/TDOJFNnbaqDr0aybOfEH367VyrlxaOli7f7Pre3nB7v6YgsiehxQFEadVLXkQ
kIRe2teF1MAyr/MWPHNM/oWpQrVZpcMl+ZAnvQUkdjaevv7eT13+CH73OjrkllEj5tRW8supkV1f
5loqec5LjwdnM8XczPq6/eTrW6m5wd+aGlsF9Kbewysdd/LbC5nsB7+fqLmi7MHhhPVLiwmpRDxk
UE0McnXWZC6Hz4l5dMrIeE1XCpOfoZL9ax77b1QJ5waVuVEm9tN33/4Eo/XoBQ3YoYHH998xw7RF
/aokPsWVrPpfouCVXbb+Gf6DH6gGCRf4ntg8i1tW5vVPK5Vc/RgO1M0BLQBOcpU2GskmRP7z+9wr
b8qulhiIpKcWg9eYBNZeb8Di5hvkGg7pMxhUo3UtwVu6Xc+zZRhBe8UuXmNe6IOtkP05DH9UND5D
2m6Sqdcl0wHVKeQqUXF2DxM/KALGeD43M97yQjuBAz+fe2Aafez/JnlnPqaWtpPoVIv16+4DPKer
RJXHUxofyAa4gVISvOUzsAnOqLl+fpQzraU9LIYyggNcVqVDK3z0mW1pW6gQncmENrTfBcj5SbkN
L8q3RkWfvbR646eYuz+i5jY6rAHF8Z7bXV5io4GQnsTAygTomeGe8LlIBeuMQc/Y/G6y0O0eOcZQ
KJOC9WPIK4AUYJHeNfnrBbXUHVLEcJyuCeP6Jb4GHQYF/QgaaQyc891xdaoNOLbK2ppD0CNGmTTS
tM1pzvhEwHMx+67fzXTch1ucWCGSlDpfuUXsWTTavbh71b/rzpKNL86vvZPvx7wTNpHBfUMut+0P
Rqe68TWw8pYkoBsOCoQ1D8v3trs3ehasM3NrKCHO3a1HwWhLS3j+UTkGU7QyuqDE5uutfUUhh8Dq
fLCm68PuqQ2dV9kZnUSrzyP3N5ceez1So5I/cF4Mrjk8NnfviBBMXWpVK+j4TMwP0T5xRvg33RMQ
4m1nQ4FmR/ezDWtb3wIdtUNUUzpKBXVPLGIk6Q4hsv1i/fSABP5J0a9RNrd6jnaiRXO6g9Nk/nOz
Al5ft4wi0woNakR1zcUSoy4Vv7YGcYijSK+5cjWm9zlkv2JSH5PA6Bvv+mCvyL7L7oVJ9rwIxHT0
dWOJWu64G51HdNb9AreBkFWl7rzmhIbUTVcR5KZXmORDFS/KOK4CAlOOl/QYdZWtfww4k4B7CCGb
Kxi7xxjFIt/jDBdzTVSTvxhfTEvZJvVFnMWavKWad5eJqtcZiIrZVFTTpC71cv+LhKY+AY209/OS
utj0GF/FceD8jfToO7RtezHoT86DY64hwmpAoHhBbDosRbD3UDLYiaVYJ5rIYDUZvBjsUnqn+4qG
vpXWrnlnSl4r2znlRd4OFJ5jin4//CKD5PINXoz9SL16lQxRC9o5xV9k5L9D02bfOZeerwkZhfS0
xVH9rdBWKZ402BIdJJP4S0LtIXxpSS2zUyA4jNshCh5nftHnJhZpv5Vee5xrt5d4IivcCQBKB3ON
DPTJ+oitohEOhRYYArIhsawjwCS6bL9uaYskEi7ELNI+wl0sQTjthPGOp84jJwZOghzwKUHsg76c
LxbAs5f2TdNDEiIm7bvVwoecvD2irNLZvZYbiF0qUNy3MtUVJ56Ch4sXszLv/8HwTt0nDXCRd2Eq
tRAfznBCePjQg8MwtN4jSeNUQ1y+2JDTVp6EWEoN68AvlpwSP8fAPwMvjh5+/UGFSValTRraPrpW
jx5jySVphovcDS86UbXkC65MHjbnRD1CMp2vR9Y7p3oF25/SLdtAWuK8O1IoKLnwejzFpcq594kq
hjmCYx38Q54+fl1rixU6uDz/vPbWLSYvh2nToGB2bdyUE6bvcDCvJAvQ7FRqPrcZZdwI0mv9eXtv
A0AzKJN38ptuuCYgIPwqz9eD1dSC7Y7sJeYXG7rAYtCTWerBVat0DOxSZOmxehQFtuAkUIWD51yQ
sIbzUwuJ0FxrOtZDYaD+BNHU4Jj+rBe9qIBLruFo2UaWVOfV7ePjmNSuQBRXRaTUaVbfq38dV9eA
L4OgNM5PJ0aYeD846iZ7Jl06CsEbUaEpmQm+yF+jH4b9gLz51sqW+YXBWyahIKdPh6UREgJm+V5l
pkgFRpHkYJ+2uscaxnhC+z1s+vXT9ASpCKw4cx6PEUPQSJ3h7kKK1tBwfIE7sy/CWi2Gz4+UCtxH
fuvDkrgueGV2KM2OnXqx4Mp0ri02WhGIlfKCWIojxHzYJGI1wV7fnaYX+jdIhZbV/MU4cGUpBe6O
4cGq/arEm+uZjA6We4rDeObLaqDeZVJcHLvR8E/bgBQCYYRMbXzn9+kc6QUl+DBUTJMklfo3kxL4
Kv2Z8+htsg6kVYEUH0VLlVyhOHZWQtl7i7ppAD4taqeyCEXsU6S/Fh30JZjAUcd+8VAZbIfxc7Jm
gmO70hxCmTkpyzYTIEtDq7U484FRlD+YqKeCa9AQ6mgvhNF1d6zyksmtUYnvBAOSjvw5R3ia2dkN
eyaqADb2pb3zOHcuAQHJbqaiDdLlRxXJgXzXDMeyStOCugPxTdT8nT8yd9d8dgFfIPL6HsqORFOR
/To3U3dYyDOe/NtE53Pl6Zrs2N3jhgrTKOi5aTwAiI3/64BdJe8KxlebMcPfy+RFHrjYFLykafF3
0oPO2QLPQKYlxS+RlfvZyE89+yU0uPQGHWjZdhGyCHAHyyT52DUG20ht334bLyb2LWENjjsqA8Ek
iObrjuN77o6JRQJIHP7e3Vv9XYBbjTX3U6Xt2M/OPAAwPtKxqDJe7XqIaDaoWIpr+TlWmyaVp+Qb
M953witswegBDmWnJBg8Saa/qI4tx2QwVUdqe3zxX6ub2JPwaf4afMR1BloXWzDNr7e1xLXK8zxD
EWqxwmw+vtSBMTXsrOqAVfacupw/NtlE+Rk9ZeSqskaXvxBNnKpngTul6k8B0kSemHk/FQia5Rh8
u/F2hv1KDSJe1oY25YJx86v1IV0KFpCt3L3J8ZYTmXQg0+oSz15BDQq2HX/faI5BpCkA8jGuZoTv
TjlrFuK33p9W2h77STovfiRC0SJ75Ez1twI4qLnzi94g11Ya7c5w5LRaJnAbDaIHzPOQygHj4zrw
kNqFCzqt64016OM1RdqjY3ZG0aWOnFqTIslK6TCqOoGztLcyPmDEWJCyi4DkJVzl8Yt5AdO1JEhd
Tfpm1ZKGhBhzxG5+1XMvDFCJaz/80xT2PUqxHoMWN6dCQwv0xjV65YA8qUtJHPgjTU+DhVrC7qJN
xoXGvWOjFaBuAXPs6hxqKNCGGE9Lc8HI29GeeMYDNs8z4XdmgMfH/DOMn/VZ3FRxc/JPF8pqISMj
VXz8yBTJE0Onzr9amuRV+03ilOJERDVl6ixMtr/9HlXW8NFLm7wS8W6qs8wmF9ptshTWTav/uyPH
a/Vv6EZXKLPkkcfQcdG7oXgt6PQUMPTu5lsXmw3O3QOeEElMONExW5cV7VEyTnmj9aq27aHDng6M
/0d1/4fhe5XqjHRT2hSMqMjqrXk82GbcSKD/Tq6eGvhhoZOwrwMGfNlK920ZUMWht6rD+a6OBR3T
i/LSGBfJXZZJoouGZoFZCWPE5bZbUzfrx+4marj7IYPSKeYciDrJFFlNtLe6dJpBsne7XxZ6v70E
zkUVm7+Snr78xe+cugLdegKGJVr1IXYEafZkRhpNP+Jh2QxeXSQvNoaWeHrTfELdCFHr2x0NB/7v
kyJoe/IkBeKLiNh0ACjRjMNtt9lZXn5d4f4bPcy9MjDpN5zTMGcZFzmoP9LncWwMxjBdgb50+Sw1
wWAJIQmUowWgIxL2CW9g2urmBUlcMdzPqcakhRUqpdAMrwq/tM6l6bqZiGhZLQFSzeRPwVk/sAVn
m7cEQj/6HrFXtluLmfJlaePGl1ImQdcMP2I7zrw/kUDxL9AeTpYaZ9s049wAAnbLgHgjCADYcbbg
5sBIcCZwV/Ib4UO5P2QRcLaTnqA6lYBimXqI7NwmnCnyoLA1YraYyZzFomTkJVlUbLuOBgRV1Mh+
ULf3PNAonbZ6OUKNSdaMN50SQLpF+LaKCmWwRM98VBeOtMi8srISwe1UkhEqm1qkVn7I8NtuDYSh
ClTRgRRZgkYjQjMDWS++SIkvuiR/PD3R3PZEbeJEbiSFosF1r4mYpurpwAAd/7CF1kwkgagnm6u0
0IqH/Xm4CNCgTW4hJ/K8eICf8rPkxlFkJyAVnh2sAT5qFZE0vtzi9woPaNvZVx+Pm0f+F0Y21iIJ
QjPYjt+wEDIJrxF2SFYxg9z1KdyPk20HfanPunQXyQkhlkDwzqiytmI/peKa2xD41z9NBO0eH0rR
vcG+d4/VEA9tzSg5n7C8f84lFMLQUFNF+jYeGF5YwFjY9pgliRzeGN/++kp4gPtQu2nJ4JbRDiDA
dBp75k7Nu59q+ieLnr/wwbjjSvly94Yg6HYlPC3zoHU2Nbsaxa/aPDwuGvFAd7feXWUJTp2ezZV/
CPBpL+f0oy2B50KTmSsr5k8ucxE7Uecm3zfva44To7eLz8BOT98TgOUl/4wOXVKC5sWWX+Xl55b8
FH5VlUni2pEH1z8zgxcWR7BwLYwYrdUVj5GMB+U9Kuyt4ruitYOLWu4Z48VD/duQzYflM9FqQ3+o
G8a2QKQ+hH1/zx0jSi+IgBUiVOGauPLFTFx196pHNxWcywXaYiNP5bpc0v2axGwnY/pXBkp1r/KV
fuionR+CYCE7RXRMoF1OfQnB9tkrWteWM9floPwcHxTBH3PkbOnu2slAnIH7RfN6veRDKk9d4TGJ
iEvo+d+a9K13QYAoFmz9vCvMsIlYICumLGAE8gCgrQDk5CCpvH8w9fd4iglYWVfkkz+WGflo0O6/
lEKlSP/AJtNhV9h0MWBYYRPdhiFYdrQgSXqIYXPG6wiafXKBPihN5g4KIPeju/HxAnkgt6RnRq0e
H+EBj2aWD0ekalOoBsYz0bQmxCO7zYYt2/UyKSF5mPgNwM6glJNl+zZQ8uV4/skegaqZGn77AzxV
/InEbOGYw5r8YZghkzn0TziMUCpbHR2s0RHokQvpFhrnGHuGmgiKX6f4iu6xRAm2fvs8tBLqo8vA
jM8UzOzZb87V0ZrImAJ1nH9QbozEB03qDtWR677ctpRw12waLMLFdT3jy8MK9nEjaC4PGFcLPh7M
UTLKQI3HMibDJZgRASObMUGnbgXy3S/WmTP+RpylcQzl1q70mI/3etIAYJR7cp6ZVvRY74q5oQkT
8xQGas6tIdMi94CoLGrFvCWB8CFxt9OMeMg4rwuxarJJ5IMZeN1JC3yjt9Ltv9+uvZ2IEq3cW/Um
Z2sWJO7Qgr+gjSR2CX5JLnWfvF+9U4ER44sTV0WuOjstMdN7SLSmJyQc2jK/IlFUpM4YwfKvj57c
yvnIeMzO5X3PiCOXzAvzioCIthys9+BfsarefDFk7YWTd1BVSqlZ0c16BOH9WdGAPk8jzZZx/tua
M0teO4nDFfVwgEy2tHVYKsCHgZ/Ot/Bzs2UvE8r5WaL0aakK0QuDrQUXIzce+wamfYgmcgBWhWUG
l8Z+6mqSk5koDOij9rJlb9OznX/FCutZ8NUeZ5YlsxO2gxgP7yGkYSfsoB00PcyqR/sjZ9GYe86c
t6QXlsZg1zm5oLUUDWCVibztqOjE8IWHU0+exJyEB90TX6WPZxQ4/Kdw7PagNemQZ/597wwQJOP1
Wc5Jp0o36OFPrx1/IWt22LZFgcGTKbUgn7pyfiUTMvB0lVo04xNzRBeIxnvjcNCcKRij4Dxe1qfN
V8syLljvCX2kYxcAiJrfZA+Vyq0Pi7ywIZVrwE8xpSfE07PaGhO0AIJsVPAc7rGmqMfgD2CW47P6
erhtVktA9Bhf5KQMSKVeT5gSR+Kr60IghsGsQ7nEQbGVib2Y0kqv4fBwOmWB3Xw1hTRPKoReF6Ir
zLd5DCYZxNGcbeLujX+T6cDjf1kryOw7vjfNhjEaeHwfa3OlWZ3sIALkB6BH9wyqLOhV+MurpiGK
BDl0+b9/T42Gk54WWRXoXGgfBcr7f80GP3jr9rUIqiH2dVgtDwUgfl8MbqR5ERVX7e6wKNBLCR+e
pr6XzlpvGko/5EN3o/7WeT8XuiLAkGe9RLqk1fLdCDBnyB1TXyCf5duH352ep+XMwytoIjVBqC27
1vMwmbDlwFKsK59l/Ifu2E2ZAoj9TZklPh78jlAeRSjVJKfSwThAUVu282cg9FnDc7wi709RpFi6
dUOZpHz/nc+mHYIpvU4OQMa5Hk4vxTMvmGnf+VaoR9QZA89VSRfVGIKugi7G72Kp2oPk9uPT7ioV
65CbYDTMWMLiq4etvqGishGWtEpCen9EVOjDvnMlUO4K3uKcL+gp4Iwhy0yjQR7zAu1KowJM08fJ
cgBVriyzytd4rALKrA5/c/4zTs4Umt413+pi2z8E6Qu1WOfCkEbF3P8j6CdBJHxtmp/IZFi+1/QP
2vujCa4CdR3uu/92m7Gvgm3oP+XxAQEGVGTXHqwuL0dMqLkBi551AFf5jQFe/8wirnMXh3YgDPTj
bkaEOVp4h/CY1v731Ay0YUVm44YrZu/O1/a/4rESu91f5nhUrhjQmINKTK5i6jiy4apzlF2lh5Sy
Tg8XcjNd6XkE+AqN9cr7zXwPBnv/ckOMzR+xf8lrKYtfxWzZ2yUR6NdD1Sj3SqoUFUm2SgHDyqpU
wD3XSE0h5MEy1MjaCyabWXsMIo7WZnVzZpslbcQ5zlTjuKQJO8wQaRniF96n6xh9rl9BNGC0aSUy
HvzSuX5lvIiH4WzRDFE4dna5EhyngXGYH1pBCwrbZZ1ZyLBAah1O3IslkN70zZ+Cv3E1VPqiMQvK
fpTglySlbQKSs+y0cBIFmOzsKWYtsE17+12FVtB+M3Bz68BF5vLjklz9oQQJ9xbrHaAQ4r3b9hrU
gKLYTc+FI/WSkLNUcQ3f0wiLr3rRhWiWvX+XmgS7nVLvhNg74O1oI0jJtWZe/DJemL+AMz2rmZwJ
c+z1O5GhmPmbXU2n8pg0K7r0xGr+sfI9ieWl8++wzrgCssNylqBT2P2T77zff3316AoqRMUgagvy
GfRx/QzxUhGgitXpmMUMJTPwF3IkbqTaw7fixSpqtfvSj4A5Ku2rt7W3nOII9drPg+k7LtjhVvRd
Ms1NoJFz+rgjE50I0GOyw+ijK9wsJAaR/IpSAolUa4Mu9Wyo/SrOXEhYOUzXOqMsU4LL9ZPhPza3
AuT73OOszZtVL85ji8kawDbvjt77v+KllFiZcbz7RMqMxyybcPFcbmO1hfsKF86bls2t3TMWq3w2
0DLtr5UzDbmBAmmU6K2xqBv3JinFtEU5e0rYjjEpA0GmbhaflqABd5fD0Op1MacxiELXFBaGTioI
fscX11rq1XZvrXJZLIA4K87HeAQVonMXZoe/LJWuyuXwdMa4QGnkNYbrETMJfnH+xaSkGnDSfa3k
/lq9/GMjrvGJm5xIGWiBdL5pEugipALH7EG6pr4TrREhB3RI0VCJSbnUa9+tj2jEDHalLUdx9nZh
+Sn4QmVNukpFMfYFymfuprCfEa0jdAJdi33bnboZGb0a5nge21o3eBrnnFYm9CR1Yjxup0DB2aEC
+/O+NhHR3gDCC/TawjsiflBR1ie1GNuhThouYg1Jb77Yna7cohLCc6LgSPWa+LDpAO5PrV6SeiT7
qBmP5MRCz+YfW+AxRjRD70unzGmwPAnhsZmy1ws2ZWDh2oPa/hoaBvLo7XTN/IKUhYhzNb1mnEcJ
UTOCPtMtfA2KlrGtXTTZhcmO+b/leq+nxljsxtpn0LFOOYg1T/EIA76W2HN7YPazPUdYXq6zn9Yx
2xC+FkpRiq+vSdrO/itG5uyDV6hndw8QfxeZ5wJeM0yBKfk4DgmRhc+p3pIh5iUJFN4gqMQd2E8u
mF1NlhVLLOAt9Gn953jWrrGtttQJF2PVbPzXwp9dLdcVcRN5HXMtZKdE3KamXEsH/k3/mn0hQ/iC
bxvhZsThxrjKi1kBzJctYP1k9Su91r2ZAh8u8JT4xgjxVp9Ye6xgM5r23VC020VEbScjS5WSmxkm
PkWDkcuvd1QOAxn40FCn8ZMS8nitVKVm8n4MoQOY4ZAp5KcrEWNToQ/tpTcI8DCSrhXBsV9PozjZ
S2EwFKGfXdc7eWOwdFcp/UtA5sWhWpWJ3qWWa2WHQpfhm9gQR2Oai6HRdQt4JHxrZL5rgQev0MqT
ZT20JpWMriJn3wNreHB0aqvYvqhJJZl/9evfWIVn0r1ASqK46bnr0o85OLsAaVRKY2gmxpaWJDXR
/NmZPbf1/r4LVoR8c+4xP7nunFnZ7zsSleNBUoUFEiXy5CUUEwVt2r0Bsj8I4kbyjkWLS4tf8e9l
R7WadsNzdbLQwBsfm86vba0aQ5cKW4a4TpBeyDHBEk4rpiJPD/nDlqaq8uf5xRpbLc11gg8pkZux
J+REMvw7dVfjPWZhYzv0fIh5nfnsI7k7b17fjwzxRtWh3+23LO6py9Si3wO0ND+GclxLV+Fl7MHs
Uk4dkZ7sDrBAXDA/Dz2g1fFxhKrhCti8KiDx2o4BGvsMhIbp+csiRzqY0hD5VHOvvMNidr+rZSvL
Edym0A6/gHyVRTB05U658kjVyy1qcVzpUgh3SIDQu5hlkdScJecJ42SFl55zwMPHHiyYAMWW/jJK
kaomjK6e8ax3cLdpLy7wwJ98HqYBviD7A7Mwk5N0TO8uZlVwa/KcAtjOCo5MkIwj4nG9jQ/Zyp7O
ntnSVySIueWINhScv1r6SSrCXw0cW86gb+44FnnnnBUUeGNwBe/FYSpW5AO8gOqWjAp+mnGBFgo0
F+lHruQPbCTxCESaOmEB2D9Ep0hri18st8iCf95+aiahGfkk9OHbfmFJQXCJjqIw+u3fK+cc3mSZ
stjFaZ7/hNUNqtW2lvQi58RxtXyoFPMUYj16LBmG7v8Uk0kXeg/0XBCyCplxHE1DxGkxWqAJmAzj
/Byv2YcDserZePnW8rFBCfSXFEyOHcLklq7x7/aNzUJoC0TzRKHV8ZymSV8VIFEcHf6lsJWvg9SB
dkC/i0AUPdNPoiM/DGAnxBnoDIiPp+FqwUkRrjaDUypvbX1j/KmebvEjInjNeCRU4Qw7AMaT8tv4
bZpzGUA3niophmDiBqE/VZCFn3dvNDo+kZFyMTHfyhzCvP8K6vhTJNWxF+K+nhkXxXGhjR8rqyQR
dG3rUE/14aJBKfWbQ5ylGT+eQ1atlmJIAq590/JcNgLA6+veIEcy8Be3VBEzwpWGSZtzYflNWHRj
ecct7BYyjaEB3BQ6Ch3ZJ1IYUSXIXCY6ytSKGNCnn2bkeYo8iDUshLJst5H/lFBBQF6mEGLzi4zw
9y1ZVWvEgUJ7bCau3WZUlsdYN4+Hjfrp3edxbvrdXbeCQ86FSnK3+EZYyp5HKq9b6U/XcJGC4S+r
9n29FpQHLxlE2glGtvt9S74ro8S7IDGj6s6h7xk2GTvX5RhadafnLMOIFMbMWbedGS405xb1lz5d
3BY2NA2bd9/NmTva2Ru9cSHZDRpqCil33oe1WJd/FuOVEzcsuJyps0F/RTjit/PTsUMzg8es7Sp4
kjxowKPzqOpwpGPUK1hl0EqdWTPaQ9X17osiS7nJAQTSZ4qsINhn27dSv9A2x2yalTHJ7oyjkQ/b
Cx92rLwmS4Gny0GJ6AtpKG0nFCqLklTH1CvnsHCRFhPblgRYyI/ozXrztBsyBamYMDXqM+X8OdQD
JbJcolMQZ+mrsH7ulLsa5WCp0mV2MEbawC5EZdp4lbkFdRibFbR6quQtaYdloWdEMjTL29iPUBJg
cih/D1QD26yocXTuVSpGY4yVQ2cjh0GQe4DMozyGdDwa0YohaKiXkL9b4BW3fn1A/lE50oSSiZxj
Fj/GaQ3gWL3ZU88Scj/5FYjg2CVC+28vds2Iaif/bssEEG5LqJWQVRt7VVHRN/2hrfwcyOjBW63G
GYZiabZ9agWx8DlpDADcJisQFYFEblWbQw6ZRTALQpF1LzDzs45RF0HklLfB01ITRdQgW4ujZJmq
e/8AKolIgoEy9e1XnjtSqw2/jwps9VuVhfCTRFVf0dEyqgy4DP4arphWiNpjtHpRg7qpUklXzR5Y
UPYKAmINlVHKmPpLDkBO8Ddi7/pWcYALv3dTcrZxFdaU6NCsAY0kS/GnJnezMpvMTwUo8vB2HQlt
TAjUAomIU5YOSnQOCqxDg2Ys/paLOQ1meQ6lyoa7Z9hl/A+13sIfuo/c7l/zRDI7wOmrrF6iDA8e
CVa8DSfrAMtWJbCq/n8ikzgEQsePt4X+tMMdzTqDUPR2/tXgtGyN+ipgTaZmk1lp6ts76yDLMnQy
Y8TIjvYGTI7kloOE4KrG21as4RCeaOi/+PTnsZXhgcdfj2YB2BNkH8zKNCpfvneLdgrrUtzOtggU
mtVc2VPnRHR3OWTwHPdbDtI2ys28eO3NeXBpCkJ9S0jAtWONTAG1b+6wXjENwdheLuvMmcYkObo+
4J2TkaZjS19zYHFAuq9rTzohffqixDvZ5szJnICq+h/WrVEGV423Ewx8ZE0iWeQJxBsbrdl4fCVU
YN3TzTaCIkiu8O9ECNYJcfNv255J3ptWxmF8feD0ZHHtf+Lb2uLSLc/nn6tQWpAYs504JLWNiRXz
KsETh1WdZ7xAGZ8p7OIaCeMmQQuBSAD9FpSCSiVn1cncNNW1ErTXOz6m/KzttrerxDbg7zKc/1R4
DujlBltlbN7v5cbknTsFe+ci0qJ72BWDTWq7Hl1T6sAtJpxtdbsMLJ7BWuyHD43Jt1qt1k9XWhPr
oRnWpcBXuEIIid/w7lW+vuP/IxJ9gX8UBHnkXny8BRqh7VS/a+Wes1DsceoeSezITIS7OWbwo06v
nSKnQzVT1KznO5oZt9Ks0nyfyVSO2J0e29hORoJuyG+AN32hYKwArixM6StkRfLy3w31c04bDC6j
DjrqhGmFgZp/S9WELevu3Ptwbq8EZStraheU1r6d3JYP7kdDfbpcEMrYNuzG6DFBBtC7v2Jenl5u
ONv7thW0gvEhL9OxznTrcIrCvsFWY2TjJ/cuezX0/MGWKki/4NM5+xnIGGqiuSU2sXYjUL/oWRmW
9SR+TdoU++rXszYZDIYpVbdmcxFGRwSzpvL7zNbfW1mO12gjaAruOjIewr56L2dpVu1ZE/0cLqn/
M0HzhkTVI9I05zfutKttcOHhhVuicJF3x75FA2XOf7UOXy/vcrk32xihdJlQLEFShR2H7/e+dgB3
iiqvUBmzoV9zw1I53E5LbcD5lfzM5jujgnGCDWjSD96DTgtSs6jAwA7fsBNDfZS8mPPeLsqwRug9
0RR/4+ADugcUn9ISTWkOVyCJHMeRfPo1j/LXKVpnPRBtNRIGExs0fDZgOBNUSx3v/NhR0pGQdnXH
Vj3agrAiBhm125rc6Rp4hI5c2Yceg7CJCNEKlh5xl2y57zUCg42hzuvqyBL7LrG8tKCZvbQdKv9f
fLYaUrXP7nFu8jLF5Er7atCqBu4NOJ2/bjGyzhW01dBhgba2UrtnDqK4wFHBbd6LZSF7KDBMyrQQ
+nYZlcsiSCp7BJ3ojWYgYPKk257roPmLy5PtGo7Ad1PlqoXU6ieRVRvxIzuB0Nqa2C72KikDVg8j
rUub43L5bG9r00/DMP+n8kJPdz6MOYbviGaNO+RMjpVFwKtQDlNCNUgcuZ5gm82U9NSjaiM/zReJ
L29mg/qb2fRbKFVchjVBsA8qKnsNd+LgQS1ojKJ5p9nyjkglHG6BUGGf3aqloxXVeSG3RYhumtwu
NT3PrtSfhRTBe9kOWjYjAp38/oyNzwx/dUrBOXZEeyZXXiIQCeMnzGZxghjsYQjF5SGQqegXrSZW
75iO2mZABOh4X7U08EQy1JOFNoqLSjDbNtJaeFUSjunebC4hx6GAN+T4fChQX1qfvuc+IPf8+GDh
OVQP1Cd1JPztk2oWrzsIJpsqhZqr5YMMAQSEJDxwMpxvL0i2Hl3q2BaKRE9v76LseyGI2ikKJkRA
2FrHVA2SbOZuSFCw4k3cwQ8iJMFu09q5Gi2YBaICFlIAu7tA2f4N7xQhGm3j3P9rKB1YxEGxZuSP
4f3rWzCafU1n4OjC7UqM9/zPJA1FF01FFXnALWc2FPIkZJ/714SxCEKQX5lrdLi5em8Cl9MIMK7E
OtT9Wvx7pVA6E/WH5K6Vj61ZYcj2OGKBmkPDisb6Yshhn/UA83OAgD2UwMuY7LYxpq2vJFun62c4
lFs+xR7VEZ0/AKnFfFJup+UPcS7eMXFeH0og4Lk26rVzvJ5gB7WB+/EcyABPesyazK0mH5p6ZUWE
yNDeCK8/zEKakUQeeMcfCl7YPGG9RYiCgygigfJ+NYwq1ArivGup5j+3pkgX+cbBnYPtNepOrX0M
gMbu3lbM1VEvJ5Fh09Z7iLJPXuVxUwwQaBoOi274Fg53JEYrPt9WR7dz5BnxdWxcT/dh6pLV0JzS
Ah1+5OzwgzGCCejESkqiFmK9+RTFvpUAnvm0mwOs6ivQ3Umx3D9qj/h+QRgB1pqDqZ+tQPTn4ggQ
kjQFsBwX5kl29pu7fC7ooVFNxQqeuo8YT8xuF3/ssJz3KdkTQo99eqj2RCmm6z74A2N0upWf0fLB
wP4Y+i9GS4qGiBfXlaZqGWjrs1ydi8wrnlM+JBXo3qizgEwLnkbnqewJFopgx76qUg/zNOoXwKtm
Ym3e6kS0JzpoQL6vMw2fTeh967GtNG/E1C73WJA2BmRfo1TT+iNfjvFYUqfC6v9/UpieWzi77TRm
qASvsOOJGkMK7zciSq72fPIxh1KRfL30uZtINBvOdeyTFoGbTAwqnNRXrfsJPNSlNi/Eul8UH3Yw
xEeDu4uwcJacUW1cp0nSqgPnc3vbzEH0760KT0dkuaIxheooca1jGlLSdijCEd+uR6Mxm+iObQcw
k7SKW6xkU+DgrLElaKBVu1vdY3d8UrSLRKQBXdcOxYbnUmX1mC/Xx3mCrZykNndODLLTrNskmb+1
p7kEf8KGbkD03f9GGX32orSNbfBgyhGqdDF1DSuvnQqZf3xk29VwlGHqBMY56lQ8zu0Yq0NkB4w/
pXWdkHxmtDlxeorMnQjuar1Crl9dG+lnLArBsbRvjSj4SATQvyG5CjM6jqaxqK04PxBz2xL0ga+e
aRCuPL8hCb4z24gxr06iNHXkseCYP9R8ixbZaic3MqZg1sVf2wrv1Yg5mDPTnhsxyWl7L6v6rIIc
xjjOxK6fEejiZN7LPbJl0UUP+b8rmQha6nRWexWvnE3jq8YnjJ3m9zuTjqQbExcsTTKRh5yfsb08
FOQCiOimvnAmqneYNEYdQKItKbtLvI1KkZGFwpSBa1DXQfhiHvrAOS/C8lDtzHPNU1ZXsZ3SbqKi
DrY8XiHS2l4UkoFniYAwnGpEFtS0agEl1PArOLCHPvV1xwV0zhspreqTB9he36JlLP0wv9zSD5Bk
r2hHO3BMi8l7R85ncg4oLetLR3P/575eh7G0gbVAzL5paQng6FZbLwcP+7KJxGWZF+0BVmCqOJIQ
szSW+DskBFxMNC6BwsEH2DRJm2IAEpWg/4nae9UIxzxsx24KoyYjvAYfjouRf8WSw0oscupi5fyv
oDTaeTZZ5szs5fF/0scbf/qvgD2E5aqc3zb/8npXb42piLAI8GS1KD/mUPrfNx5DSZCUgzf57fkh
SKFszHi//qwCk347l0zUIiIgQ4PHWvNOfObxhD+AII6wwOmjV9ywudbkwPGBGSYmHC+IKUh35YQl
b2oygwFF3g9Cw1izy+HFNlDB3+Iw3+LcQGUhBzwX5Lpm+Ob9LT9+QnK85SrWyuB/Qo/3DGf6fveR
/dGSpOFLw4lwLKXKqbLshtnHmrJlcQdXK4CyjPjpbz8EQwawo+HGPF98lG9uM8H3qPQurcF73FLM
atVgGokbM8afRFpXMCEHPs+1/lHoHP/10qqCglBZcxFh3v6Dt3r9eXagwihBsPgAFSvSoYzycFQs
ky2D6kTQ2VuCzcqYUXGHcpF9Kg1VZzbzADqiSg8FgZN185SVy/MZpFaL8t3AAzmJzb57NwnIIvbs
sTnwiI41nSDTm1VJUrgwsj3g7HoI3WaT0cqxZJ/ouaez/CaaUVBlWluGo3STBojqnCGUBCSEUBy0
oqT8c9bQwkzMcnPuO8U4b9ImcOGU3YVFUOfcKMO5XYlzr4lDQWBVk7aKN2L6fm+TORLnOuVWRsQQ
4o987mpppBqNbnMVvbr/xGAE1uOspmnshuOp2q/7wERuXQ/8sBGTtieLtLaHP/zA5BWvAaaHQ+U0
PcaLcpXtS+mr/uRvt0Hs4AL0MGaFDXLFScsLSjSEVEWbIpRGeAqH5jgri9Rw6XiObRDkzVz84c3u
O+a14TlnSLKuZiTwDeTLgaugs+81eqM5RvHH04aMT5uXMdMIdAlhWk9wSli2Q2KcH4P1k4zYaUKO
encMamQYl37kkBy3zBDd/u5w51MBpJ3DJFKioHxE+qFjOpQhadTazhv9SGI18qqHxNAKqwBERDWV
XNPbzAwSbBcACjiBZnAFhnkQp4gvCzMOBD0BwRPtWaEcSRoDQZtsPfTuLjINjQOcU0aIwbrvbtWe
lwNJgJyjgNMfUqtGy8vQZS2czLH4H+6FK2DfqnSV22V9R+3iqHXeyP2kzinAMjeQcRInI5SHNWWV
WlBfPYYk3qSo4ZPRjybQNtnOpHXXLPWetuKyLlGrZaFyimWhezX0TlGFA730r+WiLBEWB7Rz4X2n
9NznmPtmVnMaFlOgeiS/vpDehElCS+GSXKTs4M5UoDUB0RO4R6ZjkR5lPWeklvb2/HVWcZL9E3S1
52mOqrnMyWsXqCDnz4peTFxVIoQCAOF8mGvyqnnU1N8t3nz9jZ2/z8SVUSf4M4vQ5Bcp2xZpqC5g
MXrNct+Tx4F97P6uMMtY0GulC9bpxbH9jqtYhi6qXf6rk+mGA9BtsXsn+ERCJFDeGXepVqJkzHdg
A7qTwHtapLCMgioQLMp5hNBrU9F2zxPXvc5S95+jiXtU0KODZ1W6Xh6zvFjICwhJPE+NCmRhBbAi
kp8TCg9PGz6RlKxASsEB6tgF70ZyWGIza3pjEyLJUDsp7rpxVWUu4ZZj+j9szB7kGrW8/nHE3rnH
VJ35mXpa8pmS/lQoDgbRUL/yIfE4+lr+DlGLfvSXJxPlZmWth5wrHCddIcvUat1BtnMhskwTSLP5
xxfURMBxY+Ozd+PhRjHH/A47RFcQDoBw8zrqkHyW5Qa9lNo5EaR2izNNJqG6iKxgipAVVDfvHGPe
jSjhpTJBiLlupzAx4BvhymOIw2bJUuUO5LtDeFTE1O6YQJglwjc+TULRMpZT+Y06YNYNa0HjLbCR
40QxYdvnUW/CTn10jOE98WIMQ/w9WKIMwgUhX/b8YSN+2Im7irELv2kEUqZdtwyHbYTdWIDY9p0G
NBLYgqJib14dEOPTbz2vE+X3AvuOwttYmPTeZQWTtQLnH3gSWaYhwAL4JYSjDGZI69RkXJaGCPmy
apMe80ThXPlPhGx9Vo2cX3CR23jGzGUo5cxrcqj/Ftj2o0E1U1o04FxtsJXBZbDY7HBfcI9hQDTX
WzpPUHH8GEYPHkO0dxCKMjBgL6qUuhScLuvLJD74X+zZsov5w/NuBkZJj08+qAPb2l61/x9IPEwx
V1CEYjnR05I+CkGnA11uzkx1ZG7CNN98xI3snMOqbVR0nmbClKW25dQcgJ7H6pGGa7u5doy2G7bL
HKBREROAlmbEkq6+n61JSpE+wg/KWHJ2hLp0n5WRzIqMBqPa9fEUXk0vY2LU77Eg3CuQu08+Z//L
PZSRKmCKsoVw3g1aUyoc9y63nUtqqMwFmjEmCN80eb1K7kBSMdoaWrYrzuXLdV2BmKOFAntJnYD4
JHT4AhGbbE3iBCtGdFGT3hhh+2UMBaG7hwbKdjnwyiNu8+nzZGaGPNYA8PzBpXCNZPSPa/GiX/QK
pCQI3CrXRsXFPGREReLp1qSUtFXJYXd/H1M7oEPYGBF4J20ufmN6cLHYxtLBTNYKVZk7ImCkB/wY
wszjXek65x1mwP3RetFsrU5EIxIMll7bVlVmsbV1hsLDOkvhIGbMlIfjFTs8ToTnzTigQUjXgEyf
s4rHMaNmGNt+m39qhChsE6zs3wDMhV1L0S3WYV664XcPTYe6OamtOfeuqtt0K/ugdm7/6oFg7eKK
5vO9uTu2VjCAY6kBz5YbS/8Ck0TXU+DFpNsemyzV2Q6SZJvcgyAcD893HrbODbPPgxGTGTPpC8FJ
3/uH9HLE4ZNeWSnXgcsjQLx9xvbuuNzynw3FqbCKdRrA0AeAYZ7EmzoJB3oHRHY+I4aFYtDn8UuG
62VEls1kRMkXLNYbU+9WUVxZAj3MflpMbIjk6BiIiuCBiqMThHQRTBXcx5zpc+rQ3tRltQe2qfA4
UbmWETcVLL65N9U+2PIiuZR+oCriZRvZin9BDLTjJ1cRmQMxZz53/Z0M7ndLDW24afryaVTItJx+
T5v0E3b7TBYXuMFO0cyFHSZNdqg+BDZwuZRtRPSixqGFSpC4hws6aQJy2f9e+MaL6aGQX7HYlIA+
0vNABSmpN82IUW4YI2mQGHsz99vT+hgCzlAo1Fg8lGnPk2xjkLkyBxaK3FyzwEz7Vei+st56uC+k
4Gmu5pq38pA7zYuthCgPQztq7QBVhRvPDmK919BaYHfPPqv3zdYcmEm8YZyuFfURG0Qs4rrhCoGK
WkMtwMZnl+bKStOseH5k386XNySmqA6Zo6cNejp9gxLAoyOZh+wCdEXZh2dnR6/KYTJ1+mSv8XiF
xZTpBirGNB0ORIFOnjoq4ncN7WFCcN3E2SbabHMq44BQ79CEv2UqZGYeJOQzFIiDmpOuYWEHTg45
ueCbn1MEz/OlpdEzUyazY4d52Vn9MmremVSlUhG20dNf2cBADsX/L9HLb8jV/symSO1qyLBcVtJ3
Ot6tsJMSSiHzU7qeaHiplqTacLy9rLUnDEl8b7W3LI1wKHYfdHozImJBVPzEAt6oAHCt29t9HJcm
7/Ag6mtzApcsrcYO4DBa0f78QDIRqtuMeNY68nlR7Gge/+ogEjgSsOg7pUPiUsg60DXWUuB7K5Zc
Voy5mkpiLO5oJygrKLJdBcB0zIKtrE8T5vn2+VqEMDwyJwsJ/k0U0N6d3QGxLApipiVUTf/DNvQv
AayXAL2WdCfoVNOElXbzNBmajMrMU8ZpNhS57KJhJIQIe1IDGyUKedsAD3+UOLMeub8GzVW9saXt
7iy6XcElneNvdRmJUCpyyoPreNwPXoXFiVpSai0ZoLNkBTFTzZBazmcJO+QpaL1m3M6/nofyBlWj
4Xz7ZIhb3L0cc85ce64b8hZEOqnXTBTR+bP53qM1ONV5tAHPV+IpjHoJANFFsDvdU3VXQEtEUuU9
2HrmSbUTJsA7ebsZk2FbAVSeWy1tmes15VwV1RpB079Z8qY/41RRNI4DCPrH3GA1jy/kXEG0XHbv
HgT9059OGpB0LruZpUjj2d8MVhs/1xjfKb8m55OMHqo82COUj6jXp9eghMD70idglnmK+k+f4Oh4
/VkNiul8+AH6MagD7RbFSqewBvuAvRGmhrjEaZG9oiyPxPkJ73ri6GLIMJS0CoFWJ+9jtSGBCLaR
DE0wvYhjjDUPAOSNC55jHNCmKuxENZv9nbnFZRADhG5wnrzolIexuJwp7m5bYol6vPCfc2pPubFy
hFzMWYC0WhKRYdn4u9QFe4weVKSM5T5J/swZYz0mbKtC5cZq+tu2IAZ6NnF8tnPBrDw9uW3OvWNU
JPEltjqeRa5xQ3IvlhVsKUgTl0j9sNJG6MtvWRHA4OR0XjIDNvL52/jGmx8nyA739QVz0FVRyWim
Rei3ACoXfV4LbEDt+ZSzVMdhTg9N17OiEYbNkzOfkqUVuAxlNzlW4luVl5nYXyH0lD4pIYq8BEQD
qhLK+1r0TH7bZX+8pHpCdlbdPs9qgEe98QSGCQioP3H9VPFV6OFjjmE32MCsmwpJiSzQZ3BOrWDs
eN6MPYpNsY3FXSkgXnStL7kJIIRJEoQd7vSBnTCU0xBZkT/rJLr15c+y2KCF9Lx3ETXg6cFVcjdb
x1SUwQ1/puv5JNIyszaOBAYdh6C3JuiNXYKKDh+tTZbBRb5KgiF5H2J6xnel2TrDWZEfYjFh+6/x
ph87ZUlHp4gYopVxNGIciAgICOqdvGCgvv3X/hjbpdpFsbbqg0k0XfQU/zssEQTLXztxR2pcLhCc
HSI3EaWBxE+JUQOllLDnNWFNu6QpfW18nkt8ZnNxTCvoLnF5qzgMcg6mp832D8T+eo+0P/Zmq0Wl
/EoZCzpk8SbZ7SdMy/zp4cSTntIgPGMsd13elNySOodBekwSFKYy2MdBIFH29W8OGg8cvCqUissm
p4+cFwVmn6PmXVV4baXcZxSjCvaCEidtnqwYVlikbBuzHdqGOOsCUoOtU8Z7AWNPRlWzrK3aNwMq
zo3tXEQU4mxrogljlpW/PvbsaA0xEe/60ivOpc07me7kl0G+4pz1wF6kFD8jwldlTK4TzMgaJhfk
TJsRlyliqQdVeoGYosjOHLnnFoG5oaefQ/BsIMQYWol2aGSN23lrLSEkO7DDOKwYnDC779jiQQIq
rtm/NMyN2b+RiXa/szHuz4uyCZ7hta76vinn7EAJcR+IJFJ++bN6LolLToW7gF3IIeD62E7gBipW
6g6WiJloVPg5XrXv8feWpTCDUhvjQZF7t3PfcJ+p6pOxLB5BLqFdlSPStL+65bvPgqygzhoWG1Iq
lRjPrBNcPO3sAMFrscTXdk7meQSO6LGZDje4UKD45hoTCtzxAqHk9ZKUZS/53wMf6NuRNegKYcGt
yoCrQ2+s6PDJUNLS5kbG4DIAsW8mHmuaaM5uNUgecwOPXKjMyo/Hsz6WUejgNaI9wpZgDa6WR0Re
KSDJBgNkbbKqTpPt9M3uhHclooAwTsrRxYrCBLyDRNb9XqGutfmjSYrpwHf9gbG5mJdCoxjGGdiG
90qh6N24jLnLv9c/4xZjkDlpxNXbaLHilJaA4EpfhJuZOQVmjwJq2h7cXPmROto5wtXW9NNUEXVi
ndftsFe9+upHhCBegviQ0SCQgvEwnL/IreHNxJD4t23ST0EMZj8xOcYmsdOHZ6YRP+D5u4dUt9hP
HpU3jaA39VeyHQ2PR4ynPuf3MNY+RcgfXMtawFKdNpu3+1guy5GaaI7giP5dAymM2CcC/i4/TBNU
z5UGZdsfPVMiFj+DmL6XF2Av/0clYyrEFMCquxnkfHdJpURb0i3idKYgg981OeF/rHbMFEBhqdyi
Xa0JaENYdv4k7gZvriHA3kvicTrdbmBrNYcin9xcd0Vm72VLM4oAjXDPglReGmeFD9iMGmlxz9UG
9hPx6EPHdHZE2TIuorxvTJv5eVOdCHRfQ4CW+KofMVpFNt1wKR+9rDaZwgt45+cydeKMol+brGbE
sPLTyzAoySyB5wE2y7FfEQXq9EYWP4JDA6oVJIeAhjl4k8UNxW1WsFHm5vxr+8LlmchWSrqdxtSB
2ruWuza1CO2SiS5mFViAQ79/LENzqwBsk5Etj6YfcgfQ4ae3pc0qhS+Rq08CIjGCRgbvlQLuUX/X
58xkuukIKEsy7kURqXWoE40TAnIF9t7/ZPKSW/W5RB3APlrp0qyRNyOUJYPe72e9Rl/4yb6iOcVb
KXsUSj2fXHFsZKMmEorPa8YF7FR7CYDNdoWFZjyBZnOHWKicE6HX6R5pCKMSC7B1iPgvuNPwr63g
mYwBXIFQhk4n5lrbHkO++hLUKjB5/NYlCwPwPieJMGsOJdQiq27KpD2w+rq0sfC77pEMOGu5x0eS
8qtXx/yNzfd+GvvdvOwnVndmb/JcdSRTsL7xsKIOUEJENRSzFq45A1ieSSQKOaojlljaOkRrMVym
JY6lSHahbumcWyv7Hf2uxRaioLtD7jsfhBkaqxaXcpo9zPYEX1f9JvIB6k7Lb7ZkObLJW7HlvFNq
nF+WSDAGuzsLHLbJ1dXMte/j0KLBxhVOkg4TRnrfV5lWZQdL0Cz+phOzzfuRiwCnSbLB/2qjmgqd
sQ3aAQTeiclSXKKzHFPVqHGNF7q6OQYAE94VEHcqwJtUiOaT6F2B++Af3+9iEpyY3CqIjyaEHHFn
D6QLv9FuvsCBgzHQSNaLc+quKyxduNzpLdMToDMO7KpzldwA+cGaRUq6AFdPxwbX1ly9UkuNGdl1
xqCkJ/21zYwc/swAVtVmnI/hcjjgkrY4BbPp+03eCI7yzFZIwtujxhx57CMWKSnvxOd6aNogrJkb
MIPtFHeVev4lhlUZ/yiCVa00eNYv9yYngtj7CORcT5tSRH5YC3JDelETzcvWeu1CFEHp11Cuc/R4
0eyuG4EObhhHODrAUcy7XJ8TVysch2wnNqhoSQmD5vAKjxrJt9NjqC7gdHqPnq5MNoo818BMWl5r
mnbLQDYjh6kKxtF7nG+L4/YnG9kwPDLK1tsfO8Q4GqSW9SsALgHMNB2bnJ6accbtkUT29uLFVObL
Rrm2jZ1qw5ALjRzlhjlZOhBxOq7CyemeC5RDL8VMeaMxUXvlUhNumByUKcz2hlYNgcf3h0jkWZhP
TA4XeJZXd+hwWUqPpyCCq2fDvXdufkjw38PIxzMidwSZEfE/ozOiT+RblL7/lW6QPICc0jaqQTN9
aK/aepZM5vCHEVzUAo9RBDlYXmXBT9Y1w6h4ZwjhfFamBxzAlBasiL/hwYmukM/Eu4DozwDv+wX0
jZBQ9hjidmo0zPgmd0Hfm/UjC2HdxWaypLRU+ijOlys6iDxpN9NoM1gvLwI9e6PLrVYWMHz9+CFp
k5TLS6sagrc2/UQOJRlgV0sNuaZJRsivLbtgZ+V9QxX2aySeq39wNtRyHBE2V4VgAVIzJbIH4Lze
qOmVYuUzB4Zaxp3xuCT4d7gSibBVPiCGye6Q7m98aLJKQ5Habf7+erfDbHWGecgWP38LOoVJK9nU
na7eD0ADEGt9nzTfmRdKUiDsY2qM6imy9pJsoLR1hRD8XfPlEJqNfIUjlMPLmimH4pfSJLbk5302
pv5e65aeBxC8I0B3mCCe+h7sBM36qXvBEaePU7Arjubnz00sG7cOC/PZdYxrXW9oyvEBDM6ZhHcj
W8T4DHNSNnywpz+g2a0iqk9e2H1m+F1b7YYK3NX6D1WaCw5mfmUd6Plx+cgq2tek+YRZUM2SD+Kl
/HqMH0aqobrjLA94ZabnBOHlzbr32owxQ2qmi4vCW5Jab9djBnbw3JHVzkGS4l7eO5KYfpF3P9Ge
PM19PcYeFFJ7EKaxLwdOGyOE6Rz/qfqXcMU68eSBsqy0mhU5TqMo4KSEBXR7JSTyXi9aK6Lc4BNn
SnNCYyroAtEjxBEBDAkAso+Z6a0UoE0Oh2s2bMTz1+jZHF/YkWFfZFXgHl7WCqR9TsKdpCDoPqEO
gm/exVSpFRq6X3nwXDojuKO7xmnWzqCtFmiXblGzS4nTqTb6CDIqK9twPki9NJ7/eopsLPpy/WE7
aVeh2WBMe6Dl+ZHIYFj+hYiPylzsDaVJiu2Qvhc0+yUnh45pRambK2eeYuz34Q3zgipSRdXDJHST
9OajNp+jeStYaRWTGdnrowUqmb8xto0mBGhSrW4rIQMeZg955vK68cONrwEnq7AHphJu4GS4db+x
ARDXEEwPo9pmqbuovPNb4gDHgkkuc2LVq7Pykts1M21PeOciG2c70O/tILY+WLRv/dSWfW0d0vnb
lGa8KndsoEP60kVvvXZWEHwekEc260ydllkXz3Two3S2HO9hnZFe1BHdiUHmSzGv47n+1OEArbXe
0bCdzm+Rg+tnEPH3nAIij5ZZEWQCPxcmn6J4Q9B0kyWMhS6s2GjmWVxtXen1SVbKAqKlv0HrJHOO
h6g9s2CW53MIh1T0r6ipDIxjWN9+bK2oajFXEa/ul6CSz6biddMGfLVGeAUiAjWASz6QzLPYsItZ
0pM0vuZRvcLFtydqLz9nNkjZG3RU2k8xtzuOcoWuSfpiQ2uilI0cNBwjinRRIy33bRY7D+tZXl2D
w7q+97Ovapb2BeHwWARBKinISTIkMabG5A/aDQZdeOLo+GUsUb6BdlgHLiyYoSx+NDKFqxUuEctF
L/k3O75iWxwMWpJgmBXAFyYoU6YLXXFi/+76rDlUVGJqBF4KB0oZcvjCL/SxQyTCQhzaNFkppH5T
W91hRk+ucVqDlAPuKnlrIsdHwHJb3/eF9gqbu+0m/xAVNhiPKU68H7RgMwhgQehgEotYxj8Do8ag
NvtasTuZLP+ocZFQtE8Qol8kfHTzmFJhuwt/HWr5L6iHn4vv3fmIqbs2d0KlMr77vHUaT+uiu2CF
ZqqZy3qciYBg8rqfewcA0ofbZaNEVAwWAi4eoyBISWCiZjxOf6VqnLfGJbx8Z+PSscP4lhj0axCc
mnBV5L8hVvkjbpPAQSQS7cU9N7AonmvEm3dJqknjfTaddPBFSK9XN42VC0P6Nnd0yRi2frY3Du28
HyGjZmlCaqx+tm0o6s+sP53BWBcZP23c5m2oqZC4E2PCZJ3iXxnAqanCi78kqrsDnSB/ZDpFTykR
gx7M3I/Mrkwo+dRdrFc4g7uBovYrPb1uPkry2P/aapQsm5tXW4CYGyYot2k1a6mS3Cb4uhmJ7jWa
ln4VttbHLgAmA+1ryTg1b/shpL6bzKPXv3cCj8+UWtF2JpRfI/Xn0/ulF/Eve3zvZ6kYR6/W3i14
34etqts5cWBBE7/ARUrGMsZ7DPK6BDq7cGGxARVOLgpxtq+8Ri3hz8LjDq/YcC9OU2jpdUkA9YMZ
3FLpV/dFPe/N0F5+fkbXRjQTNTqxDXV2Aqg9MLZyJW/WiyIPNsd1Eqziml9qecjEzgpitMhcs6TJ
6SDYRUFqId0jaYMVdBSgNJFRyrAvXbzWlvJVTrDOvFludVdE9cgTaySB9YL/7Z5ynMtCCnpN4pkW
IEsBk71nXK7S6Eft8Kqxq/MnfEd0q221aj5RcUaxtP1Vl73smFuMGD7rHKEFlj95VswoQJiZH8c1
iIzvSxXkh7xu8yHwlOo4XVmAAuXdncfW7M/JN6YC2taVRo6t0sJSu0tTdbHeNcgnWD877UUqlnZo
Y9ylsUsqXvelhKgprt/++Q/IjhbsBGAZefE4Oaa6hH4tECSNJGksSABBTGend/JlyuS+VBzjo/u6
ZNgVxx+PTK79CChlSwqxQAd955j+NY7Hc1QWKy0UJkWVdb8ZQMd+f/Ie9+HqgApChcuKpMZp4HRN
Gu4sbepOTR64VPWuZcpQl/h8H2+kZRA73b1YOJ0kUPxv94fbI5X0GNI2vR/Rj1yHvsqAtfU85UXp
/cI8lh/TJrJdt0WwxSZ44+kRCvlA2kP/l5BHHXihtX9r7p3j54EQvz0DcIUrTysQS0RFm7/VKVKf
CEALAorFiitbKb/CDCsIKgC4W1I2tRiP4pK71GJCfk39ZN707qV2F1Gcq6kN7pEWlrqyJM2xEBRD
aPkQscgBFkDk5s0y7sgTC0muJkrcq4948BNFhHFzUyl1GSxpZ85Vm0Qc0YgzCOa75L5FXX5G1DOc
yal1k3afOjJLyy8bLL5a1Bl/E244K5G/lb8oBuRl7os7miFwYvis5l1yBj5pvY1HAfYsdtfPGORn
l2Cf+T8Q4Mvh3Ld6DSfZwRZXXz9ikt4g+xKbcZLS3+w6yhcE4WD6T25QPOPNPWoWXx9nW7+GdtUC
NDJSpjU9sSfzJ29Fi3IskeevC27DG0hsvrWNiAxLEy/LAp5qmBEXa4c7gY/sqC0EXMCVJlPGA2S+
JH4FuWsUCRvXIPphGAiHaay6aSAuoJ18OwR2+1mK9WWOMA4GjiVxfILKzBlvc3FNx8vRr9M91Urn
on5Gc8LFY5t9oqKVPbLFdFFocjrSfZutk68pKa4FmwumKUVijTmpzv7eXRv9OeAv/TWPVkNNmu7X
lqaZMoqSNaZYyd1nwaVlwLSDCc+lSm94JPSKoIrxaPPtSeQUiXHRoUJ4/tcFNwNEBANvQ5FgPjlW
//1P5XqI7VRpqjfTtDs0pOJIGepnTEN+DHLxrRk2d32YuOq++P2QokKx5nmIwJeHOKJ3ZsRxh6dK
JnugdaMKjBKCziIwLCDJuuBl5K34KTZhjdo7igaCduVQhw5RSSe7ZYMWHlM4rJuPl0rHP2G827EK
vgu58qkUBurG/ppUdU8OsdNhN/U8OhXAA7HfqEePcsd6kbT9ZZ7FrL9TIKXQv3vwsjBShA4QrcVK
w1GtJHE+UmSTmCdrt9jH8HcFrtePzNhQTHhNsS2/MBA40zgJuWaABdDf7te2edYH+rTkUP/JezLk
3V7WTWffauW9oLEjdR76i7TYsSrZIT9JSfNm0VzeJEDyXkOBlFsGnBSuY9xfATUsVO66QJIhPemZ
gOWd2M9INATrW/ton6I5jUJb9HMTZf4sA5ainHJK6zLA3p6B3CmOn3V2fColZQArsNTpW90GJk2S
WBZ3Tya2fSF2NOU8a+YiJBUrxSCUtH5p17J3BSXPnx/QHFMLruL9wAU5ymcreli0gvL2Ck7FLNsH
NSyJkld2BlPEKJvJC+BtSNRvjJbkQfWN3D+8GZJEkF+gYQtknHe65x8XLHu8Bc2kv4+W6OXDU+iX
HNKkq4uyTT90s9yq6KiULVtHVF+KNxTL16xpN+Gnqt+l0b4XjQr7oyLaza1rCWzdy0ILUmxSKpnA
rftss4jbHIgMCEbs+CT/rnED5gkS1baO0R7u4RgaFNCHdgxSX6S/CLISnZtDe270KwKlqXuHSduD
qekTcczmNdb2fJw2CaF3pbgxNSGkHfGdtg2jzAUhEOZbJfqy1op0UPSzDte4pRZ6pS5rUXjCKJck
rdfzIXYyQqJMq82MOzMyhvxRBXqJagq/b1IeBOLMHkLSKlebAP1blRqeUzH8ODvLb+aVy5yg5Nt8
HsJVQf/vguBiwSfttjaCtwSc9LTbU/lstqq9oPIQg0TVnHLL0x50txKUBZR6NsIlJ5JWjsT+5j8U
2IoJcbcFzyW1XJRqGvYxcvKwfUtXy+3JMMVR/atgtRY1JD7nJGxJwmFDwp1BPkPwe80BunegAywt
cKaLin55V3qu6bVnS4hKDKgOZh7X9fx9RU+Ucu7dx1Agt2uUAhvrZIweVroJTDOfYoo2HOhfPlCy
fFAPnD33mbqqV93ppyBz7mIoSVATkpe99zzaTRmQEf1lZHN2Kglc8t+sBQaGLyfCsHDtDzyjP3fV
OmQN7MoAHc13WgzytsjlqcuXXiCnGiv9GDVduIqeth98A9JDhiQ73wb30PGmmTr+gBzmSr1av0Sv
9SxcONDMr3XddTU9JtQRI47W4fhjs82s4A/8KxjSu7AgeOubKgPEFhhWAMLM1U/iD+Snm7JeNjeK
4HThy5pY1TL2j0Vq4jlXs0jeCtiDsCHkvQk03Ve4jnnQZakeyEXnFbvoPc0rN3ncLkhFTiLO/Zqa
pS29SwcjiE+G6GMhNhe17KUOlubP/UxqHazaWZlgFkgKhrgyQ0eh6Z2z+2bsY978hFpFT8+UKitK
0BSGn7yXJd4X55GJKI0Y50IQIifm7jBhRNeEQnPruhIrJR0Zb14+fqtHinYTa6r+2l9V5WzajXhV
XDiikW397mBDhC+J9YpWVxa3VlVPoqqUOewobr6r5AdyBFXonE3fg5tQ7P9a926j7qAkMlC8Ft1p
BJeFRo+WOBIofABProKG45UIKal51DrczWCx37Y06q6oJuEIzSNjq5vtIDh4NA6prDQhx8lpG4va
8TUhGIgD2m/T9OXQdyoCuuoy0PGRqM1TRWomJl1pYtZqt1eM/hChcyHjCSCfG9+TzWPiatQr5XvF
sm1YzH1Vnk6TlPuEyRj4ERy4OKaWxMWgpB3J7CS+rif9luEyMxXN+Hql01NoRctiKctIf5xk6xen
WiwYwaQaxmGerv9uQ/ly/aykwJICJlGMWHHhLW8aDrcBSH+hkyYQbReRproK4wiyCKSb2Z2IEyJC
RZLqrLofQ5WB8g6/6nDWkeUYwmSrtRxkeQHPilZvT0ecZF48xfu2T6SJramfJc+ALbN3HENlyNS8
TZtzEADdNpZ4NLCFcGfq9WVVSvjqRZ/5EUj5fVIPCLYkrQt3GW+dEAs1b+hpA+jIXyiACu9p+7NS
55k0cy6VD87iMPTFoh0lp6DEhCH2pj6UU2oPkc/xAp4efvsm16Elk8AYDz4w58L4rcQLBiZyOeOV
ZlgIL2Eh9cZaAZXpSnfYCTUpcPQxbLvHRUU+U3ZkzI+NuF9DGFxoa73DL02dd7BFeL4D9DlPMHc6
M4eK1TyGjHvq0cTkEFpy4Vz2kicOhUTUSTFBeLCkXklFFZkg16yXpdYPgprTZX7Sf3G++oFx5x/H
zKFnV0UkYt1Nsp3Xe9XupcyUN5G8KVgWyMI1+u7nI1xQmbSXdJMCbtpavO6EZHbrgzMU8Vg5jRzh
CT1asFyJzvptk3l4StuishfEKm/OXsmVNQuo5d1TtjAPsCmaKAFXvH466za4SgL/ANYUWCCNj0Ww
SjeRhnl2zygkYF+kF0+BJakRJuSRwYmOG1wRKcGBghgc+6RggEh9PppYbWBxdiVCRVGbQAcvewyI
RdaMj2so2sSSQc/F4MZP/nOWJQL3/n51M0lT68mHAk8Hwwv3MXRGNJN68W1j9WFXVFuCzWwycm2Q
2CNg8eTlUuQqW9mXIDokCgwOomwRp2F+sfz6b8d7uBAsuQtbP+234oc4NjORyMGrITbvgdMmOwoG
6Dd601bJ2WqFYv4QMPCQj+aljIfJe8Ba5Q+W4S+cl59suo4TVfgOBtINKP3QUyYkdm+kDH4Y/LVw
q9N/rbjfQrkaMg2GHSvH93Ci7cvzr8w0UTqt7dbZk8wpWwAuwJQ4LAssUiNwbnEw/1aseMUm4ncd
tsjcZr6WZa7T8Ql7s65MoLe7PgpeIqrFd6iJ2TpuSc3sA9aJmWVxUOK7e2qveX+C+iZ743eumaRS
Zn8BV8ZgGT81TWa7sn+IlPW6wC6IYQXnlbGmztPYTtiyFNMiPBB1Sr5cR27GZSPbbqK48s+sE5nK
vpoqlATjKmc34B+le08IOJ44P6ckZCazklDQnDed2aHQmOaEdXLXNpZCvigb97NRM/NDRb+EeKSi
oafzkJ3VZophbEVLBsE8KdiZpirRizFgBWfsdnfr7zxz3FMkw3YuMubYDuet1FVpzix7LZbdaI5/
PPd8W2rhym7ezXeKOkyLmWqE6bx9iihEsSt1NRaveYbL27fqMiGuadLgqRH8lGb0+LPWJOmh3ywH
JA2Rk3fyN8s5WcsqgZ0zEWLY5wROZPOSt7whJO94DV+atQeemOKiAX1a/GJoH/P+n98PL9919U0I
ZB8q5oYsdJyKxABYmUcqG56Yk+DUtPBYsafGdfj85bflsiVhskPgRThWYu+0uHFMCWmSDiDEjHsW
YVtWIl0M3Tg+qcaknvpr1BpO17cDBD7UqJ97Zqn4KmQQBGk4g5+MvhscNGd+ZEqtY59WQUxrM/q9
GDC0MkRiTwQM4S2i/J1sHSY2YKIk4XdFPgvAA3AxKpdgfb6x80L6gKGR8IgTdD0jh8+MfxuCRc1r
5kc0loggOIqieaKJR+h0BeIL1HN9vF/U2FML/BUJmOZsIdJnNR9yHgDkZAmRlyGaMJbIr1KfnI6O
THAXd5Zgl6J2yRzCy/PaNijoYyewEW4ROmrbZZPvOrDHeM6/8RKA1yQqJ+uaNwrAeQAfc1NvH2Em
yn4BJYeMZyXALv0Xj931IFy+xtNISAD+iDq5pyeDA0HZf5OGl6zyo886Ce38e1crlOCqQEHC2nbH
8MUs3j2qf21Dl92o7MmSC260egtuhmkFpWd7Q0cDqJQqr6pDkTVDhrMIKJj/Lu1ORWCxEbP8sDAk
e8+brHyYVtOJe690FcXijlUUuXBEGJU82XYKQnY9yGOfSe/v6nbuWTDSQB4r+SXqOA/gbc9zMawp
ndlusR+1nJp6ZeCFW698UTtJ831PrPfnAKUVIt11YX0gGyHInm6M12CRyAZ1YUFceTlJOm7YGd1E
QSN2n8zmHVjXU18yS+lPZsvZnEZQU+DCgAhJQ5QpWv8JmVApK3WlztXtzisXrQpRDocwxYjh85eU
m2j7Su9CCrKFh7R90iiOXjkVnLj9PvemvjNzOAQKyLcvmS4pTAXbT9t1NKV/WW+gxRQsoYozKyC5
lMTopqPEsFCCUnYxLyOImBiix+EQL4JhTY3e7gYxQLh1pA1/fX8F+gqley6UdpQBMJ0d7iybVq20
6mOAvOw9ES0TJcb4Ijev6IU48Ep3bo1U/PI4f9QPHe78cqwPDUewaIFjovdoMjp90wjcmj2zulc7
v+i0ijQss3ZkCOfuuJrLKaiEgJu9tBvxe0XPKtuCJX4+DE8s7JWiS0E0V7q3KR3XLCFrqSsdia2B
esXxUlM4djQudXP0lM4gmQUpmn0U2Hrb5L+U4+sF9d8x36A1qcer7OhO/TUB1MGPW7OePw1orF0H
DLYHO7szinGIAO8Ax47VoaIwtB8NVzK8Lh4oeKU7ez/TYs3KcyEckK3DNawrUqgN10PyVwrVt8tr
0ojmkRzLsbCcvEapCcaVBiGbW2hKqysJuhZcDOZzmF478IXOo+5zlsv8Lr1xenXqO3V368hWFmEN
s60Kfku9QpCBfW2IYAhyspda9pVKw7LBjpn3ZkHm+lGg1ZZN750uaLOZ27mYYVkLqjuo2D89Ke2a
GsCPboWMs0P3WwlZRuQou9yUz5bzZaxKKQy6zwYvQmy6DBVFAynjw1qf1haH7w04s4LJumJKta0s
2xthyE6Z4k/NJiuCiV4yBLC7dX6uUn6m49nkGGvt8bW0JzYIxhC7sBx5xrb1XD2+92ptFCcD/5H1
1zJA9MnOF24H/iAjxtxQZPJKxSwbt9CvX317cAYRLWvCbpLjhoA/Ha93RaKkEhtYzll8rSW/Fmlb
GBFOE7qmOOMpcJPUPe7vZBaIAm60MKeGq4oruAmHtTY7y1F/4OtlC1kMM6juXQ+Av0uxuiiwm5eC
HP3uMBuo2onAiYB0lOrV+RE5r09jz3S94h4nPvpiwWIYW7d+K+VGg/UcDlb5/0ej+J0KgL2hyEh6
4Q0MtMdDEHPAqU4tuVKA+g/g2dJsVF8Vb68Hd3Ik9vUCj4U7OBBUy+PY+zRZT5vVunsbl4xj8eY0
mn7qOxYvy92BOTrLVvMBxUgJtuv7cztIvRdgavO3E/WinTMSdHgKIB2v+L91UwlQ1BMj6XQUlrws
4BMQo6Z0LTqSooX+Vzl8w/r1HLWI9S9n7wu0vw61m3zodasYeO3Cs5YR2W0MpNvmydKGvzGNedeL
g2G4kBeJIXYFC5xBzNun7UOyxE5EjQDMMJLyoAUZcWbopdI3lcH5hc6pCfndBSfvRv/SoGtk/N+7
N+aM0AZnlUfLWGFIxVpPK0+KOT2Js1J6NHNT9RlztWx4ilxp9ttGV2Dd67dYV+lwh7YfVobvMWhT
0T3TkwXcpHQARAZv1/PNZWBYsSa7owqzmecgU6Hi1RBEnNJqNmSVwMap4qkLU+REEhGujAaPYvBS
oII3puH3LEh23ziIsyL4M24aSMQ/PU/WTpDZt9wtpmKukgao7v/Zc9XYuBkJ1w55YGxPha9V8wSa
IZaV93hwx70wq75ZXXvLVBL1Zj0T0zOO7hWw5fx44Kivl4P6qiLBu2vXduKucR7rYQPqAlFQnOk7
/S2iVIiFrhPFcicdKbUYhHT9Swc6tLD/OanhPzSwC+2LisKOp3X8qttOI+7SuC6avDuEwXOUpcpg
NltdoB7/aLRMcn6J5oln6YrFHFj6BcHG4K2h8fb4LFRTUClb+3SnGoYhruYrNDI4du8fetod17Vm
wm9wk3Y1VYjruZdAeSuMFvHgfQFZjrvv6X4ZFJAyv2SJllT0lCHrekD/mJARmTSjGzl37VijmxsT
GbPTORZyT6lrfqFNj9hvarGFTkHb0S8raZC8wzbM0F+DJNTiywCuaS3d5tk5brmk5WTOE5FjAQUG
9HHMNxmA5XPjS0TCuuSV27ejf6M4M8dVjTCcUHWfQJqtNAmG/hPamsS72wxzRx1Y2yIXH3a+Bcbn
EKe8aE7+I1Ya3oneCWEQs9YEYMzbILvSF+/mrtCKnFRe1XUffddTUm3u1qOZIL44GtTHBj6WJcLz
6HeQWUThk45FbLqq8b0B8S6nyjl4l02tqi0Cop5fIrZhB9FO9DLpoenXYemjV117urqt3oL9ht1e
NZWZh9A8IESmYPvfSEQOnF0vOFQRLiLOx30m/Nb1VK7tX8N11UD7TPWorcEono02AT9ZewoSpt+Z
OdukQ0mkHaTqGFN3uDAbVChEdnFfRlmNZ0zRrOMmEyOKPg4+fFzB25Kx0xcYP7i5gIal8OfEmagN
8OMhO6/F71H2JASEoVIJhtdCG+DsSST4udBSSJllEnOKQduU9A36rxZHAeljHIUIP0mRagvCAtA4
FyPHN0EbJcjDh0GliiP2AC3YaL2RDMj6NXImdBok8UXbiwqDjzjqMrxSwhcDJnKK1LHHx9e/xy0+
LHnU3IfKloxlUAFnt0BYi+FCHmiXe+2A+e31kHkjtAqPmUOxJshLx96+6WOVaTkDpWecKsRuelHK
E9tkaTNy8xob2Fwbi+OwzA8yzIDj4eEqCxFAorF5SCSPX8XRMFdPKhPW+E98eGB4AFzQ4M8IDYTP
2fb75OP9acU0CoEbOkF5QlrS3ADfM72E+mU72HkY0X1vka4A1a8fh+akjy+l+hvGtcuMfn1Sz+iN
aeTpmZFoZtMIiAaEfvLHEAPxrXhznj7fKURVcL1R+ZySUoOhF2TqP2uo33m5wKa00puBbPwJaxGS
9SE73M3/JF5zLgp5011nHB+ri7nzojCpm6AF2Icxac5puZHLzsr0TSZHiWMsxQBNHvj6gSe1t2Xp
BtANVLJPB5bydpZldlaS/Z0o9TviVbkRIiehIgnPNagc/c+HgfT09HQYO4LJZJhLQ8rOpoHaLhu8
MlTZtuuq6DjcuXZb1UdsHZY4rzNUhLKLyYQ8184xMMb535mw3VFIkPq4uDoIJvboz++KTT1IjCSs
R8MIYNAb5HEu7ppo5vl+guCuoPlkTnyi2CB4JmPsjv1oEz+s57PFoke9WkT7qn2kU4nhQWOOAyGF
ZWgR1kiS05Zz7RgC7BdNkg7pQgCu52IIXi0pb6Qzxfnm4E4Pw/bMcCPy6m3O/MPE0GgBa3DQRa+S
weK+7HbCad4bLB9e/TQrsbkb89tVTYxcBaKKqdcO2aGp/yb6VeaCF/8XrQ8WbKFCM7bL9P91YaS3
XiJc2UfylD7x6+uBt1lUk8hPkqevGLj4/W2IbFf5lT83yt5niHyGO5t+LrIchNWqo7vqFzMdtlwP
cWm2+zLwxP9xZ/2S5cTj+j8XA1ISDD8EOJFD3gbDUesH8X92eUdhuS78kh96LUD9lz5uCto9tH0B
8ndZyHHheUvr6RClJgu5lNXlKwU9kQ7UeEy54LoMwXkd/KeE1uOjp+6WTSa/e1y+PKw/NDjFwvWr
ux3uozKvADkHBtjuWOLntXFN/YfIWk451y0rJbRBatlg+C+LFPFW6VIPvoKapjEqD9tGu+PxZN8w
h/ZSA74duDfOznCjz0CYQ1rtHh9jZyJwHUGj1wsT2GfHi2+POB0qHv0cJr6EysjJ6g/lcySyIDd9
IxS1Un2JDBMrLXjQZJYlLYxpU+Z03teVVEYjzDMQrKz7Hk4wqdTg3K1b822/XpVy2npqlneDSiTA
WYxBKjRzc+qvUyoLrNLMeeXSqrAKcxjDX0jHYGSohEHkdrB1vrBSQz2lXTMjUYHPSaOQK7Yh0N6V
b/eWvcBE7IbIcP0pO+ipZkZJGI/p2/z0W5RzZk1jUSM1avA8xz09z50VdwjWO9a6U+IQA702lEZf
+DeA+psCvk7owmxV6K2I/IQUqfMdpM1h9I9xop1A2DLOBOkY+KaSop14Fn8olDBAm3t4Xz2HPbY2
11vHjEUrhabxZbdp1pdO2eAfQMlLkeTEo2ynO/70h1R8C+4/Kc7808CAW61kJ8i28NjCeofiyNt7
EAieyq3JLeDyLOLBWRude6vSfKghyOpOYDKe8bJY/m6XweXyhcL5i7VuSwfaqg4w6sfqUQ7iaUyo
jj/YDPslBM5G5scExOcPIEmiZaGUXhT3PnVaMz+HLmSBqraJ5TNAF/Eo/5JvB2F49ysVRis6jZRo
hnlwQdrM71Pr/iWXOXGx9bnr+Qm+VCaOLU861Q1eh8fe3QETIXLhMWrQrfR5BVnJG952uYrMFgm5
I330J1kk01EG2cy87U2p5Q6HFlO73avet9iPLmOVddG7ZszgOWWRRmKbubz8QMVTnU4tfcbS5gHo
uT1gzALVV7uYW0J18qiSfIj+2eLuqe7p0nIq0tjmYr6+jFatEbTUvrxT+4N0kSyq/aa3g1uM7cxk
P9OXaigE0WF7hdG3RRyim2S5Ee39nYyIF3+y7B5xuuDDzjEluKmKuGa3pkNHMcd0oRjyUNYWhdcI
KJMWuGgXIdOD/ZgdXvKQLbTk1im0DtmesG37NZn5hC/RSo+ywmeJgRR4osow7KA7K7BrifQtTPwd
8bID6T5k9WgJsWDzm65JjESP0GTYFDLuIt73crN+co4I5qKc1WdHnNV7S5wS3HOWm9xJ3irypTXk
d5u4T7nE3jMRfiXFGuuJ0F2bUhJMb2GD/c1zcAyk+9QQXAuHAJID1Xl84A6/tPVN954dQalHN0Ug
V9OeS65rrHtTQEVnbNs2s0vF50MZgagToJtdZbQLVNi/o/kvl5M2U4H+w0USZoE0lN+Xr4eDYKPp
ccjtaEb+cNZVtlDVDqDbM7wqd0r7HAtq2SG2fP4l1YV0ZRMThBTxNmSGbCnRM5gPIgd1qza5OwWN
HpdBHmTkiaKFV/IkJfUHcJYuxy3oiAoFykVuNvFg6+sZBfe3g7Zr0oc0jQGpyhSKUldcausHj7Sz
bTE+wyw9EoJMf8fBcaIXDCC5GEcor9vFvEJtg6VbH4FBMesXPKs2VOgtsRNbcYzSUzI7NmJLjIfw
BKXSWE7JFQHktBvWfLhEeDg/cHOL4m/BMIQY8tEulBsPYZK9K9VBCN95plOoVFYKONuu0tTtGwBm
yUZC+4zbrYYvncs49unAOpcThj0kXYpKat80eHFVSFc3WRwRpCzw79KCLey9NnkFyENVPBdIWlYP
pUOkSFRtzt2wx74XAfotDM4oafwjFE+V1/8S6jrRLLTUQ027EEPBNo9a5VBNqt2tQ8s8WW+O/fXO
MDuEDCHmjyy8HkEar4eF3aj/qO0AQZR+zs/anzbRkdKObSn09OtaXNssyW+r7LbHSV/tY75mwAi2
HxfIpMo/wkrnB3ANFWamROGsjKmQwWf5Jt6iHmZ4kkToRLt5ABPKxUQSlfsaEixbyAhCaWTGFca5
FUhWDVNCUSz+DOHU0vksrZTtYQORaiLY1FYPniFS3VjusdfBQaBOuhjL5oZ2bFgQjULWvsL0STgz
9vzFCjKCOd7Mm9jSXR0V3siygjy/HbukMHYZ3VPno6pcTIr0nfHAHoxlKGhotgyqOqgRbam3+nhe
0zAd6CGLcdOaiYsaL5WmfDXKlWk0zF5lDy/nvmDlM71CTNvgKe6Olro+u5XpvSbpLetOcV0/YBsU
YyqDc5OSX98LbYFP3C21pCvyADGfhAplCaWTv39ZXWfTRq0Y2P8QY743FOZgvivsvo3xuIdLMeIS
ekqH1Zm1MZZk0l11wEB/EISIkT0gKYMiZov2pdUfW19z4v3klmYFxkXMKoSUgQLF2mH41SUpeYEh
o69pOwhoWoM+XLbEuRAuvTdz78P4c6O8GNn2Ss0Otozp0nPWceA3Jm1zlHPktzdlwxd9uJDy6uYW
N9l7LNtO3hoFWt+NOlD9Q12OOq8m+SAas3QqMs8EFI4geDhDzbfUHB8xHYAfA/vUBgpFByZT8tzZ
UyZiOXKCT3SHizt3g5JSxYrlmVLxJt3jubDvggmFyBznMm83gGq6xpUarmpKWJHqDWu03rwHkn4P
F5jNApoXtkbzepVsNR0O65d28uBQ7MphgaeV+SnotMu/UG0EpKtPl+KDxVtev2YMUhiq20zlc0Y9
I9zOeno4g19At4/Ez4gkGiC3XeBdPlRJMGk9LDQ5ISJ9XzHep/7KoMJ0wi9B5AGTsFQrO2x/Yo3r
exsxwGRAf3ZWSRvQA7blj/hWw5dqzLJrQhrFykMH635YVn5qL7QN211GsYo16Mwk4PWHydjxBMic
P1mqtELLBj/mZ52gDbzhlsRCiOTCfIKBsvjPM3bi0cjTpRKZEszp/mh4txJq6vYbttW3tkPpOhTe
RQDxpeIZEFryciLeSa7U2hCkEWlxPa7+M9e+WTfeZ+fvpZfuYqk7HA9BSxL4rzC1T0tM1L6h6IH/
y4hrCbjZMQAM025tOjwgeeiHugSDG5GIECRnz5NzJgtg9cqV59DjVGSrCsLElfdxeMPP+5ObbkMq
NagvPBweQ0bXl4IbfSnRhvTHbdfCdYy4HVTwx3Mkh1Up9SHswXI/bikMF6uDENauG7t7Wk8Gfp+r
V7HJkoOD2cJiBViMLUG/skfo5YTKgbRqj4xbI5gs5v/WXxwl90asospdzezf6G8FjPuNqBWnACoA
EjvP1cctrYIICGPnHdF1GbKXMxmLdaCswunM3yXoo+NHhFKLizQgY07ljqa5+hzeaXQcjjkudVWw
1UocXgVLKqa0Xr2b4c647b3JzwxazFQkiwwz/tT+P26w7hdkxW1Qs+R6Um6FInE4JNtvuG5/6qHE
OcagZNxOFw2twG92B4PgG3NUZiWjmHxf4HXlHHd6NZDQQ8rXS9qniA2CUh1AfnMo05aHl6bMzrQa
DqoO+xWTdMCW/Z4fV+rs3R4IO+dDHRYM/Rtprq//kZdYC4toZWmDWHjaX1c9gYwgEnPb7YewnrDX
u5Ecd2dvJHQ3tkdEtwcnydX3YI5BQgz8bDCs9gxEswJJqlYXYdGrrqUwYi/wjX0mHRRL1oUtsBx9
r8fzvyLr1hg5xqBAeDDNhcQ/V71LTq8tqx5PzFAbg7w+/rSlEG+n8E541EaKXT9MHY1q2MMaey3y
5QnXRO5brFIRBPi/IG94tWHtd74GaaJ/dWYeg8FlmW7k8NnSzAQn1Tg4k7DK0h0IOKzom9CDsz38
1nZrbEQ0KSJHSZ1urqcNKnY5z+OGtZmZ2VEkwzpSdEAm9GY4xOf6qooXxd0+V47YsKXl1zkNEbTR
XRGl0zCBm9bqFCdxwr13dpqPmzE1tC+CFxSOoLDCFJJUVqJovDbaFMYK0jckM4AnANDJftoh24mN
lCpmKnj/gxP1ULmcJDNn3/bHDw5reVjwMFo4Ji4UJGaLAyq3repwiPD4DTegLkROTlR93wUQZbxX
KCFyfa+PtgylIiDxcwhOvsKWf+I0nTu52W7AIYI3X29Q6HvdRmZv+fwV37ctvVUjzLo8byOcEHds
uc2w5kXmF6BqTD+UJufu+mRXCvF2usz1JnmgNPckc4UBhXoEMG/ycpQ7yBlRbTcaD+GrAGVftWUT
0VAVMeie3pjb4o3/wc+MDrARCZq6e+uAc9o4iU/DocCzQuDGPCmlFT2QGwRfZyUIKaI+ODdUMwtb
i7mpHDXBCqzpmTc/vVJsh+28DMAI1indKMmeQmnToCJTZEW2BuVfzUCKSnt16DqQxvOW+g8Z+ihS
dopEi5132WK8UX/RL0zjRnmF6BqYE48LHFuQyqcbRooFN5PubTXFh+4Bq8RCShsHWjtRPuN/XPh8
wOs/MqW1CTa7cBhRmopkjuFjqbHVgOe1Q3P+mfq3DVla9cKL3NklkZK1ANAEpj/dIptvhw0Z/hZk
Y9OpJCQO1NHrRih2xyiKJdZS9qWCpvOkC7kB/esbT2aDSeBJWsWASRLWKl5rbLsjsBaRB9jxS4va
3MZqkTm8X0oFP8gX2aWH7nbeEYK1RtknnmU6H7nKSiTTm6nPkpa2YADO1mGF4dwB2bO1zLEGTBOK
eBINQ90GHj+21Bdel5lzmFSG106vkUmmlJQ0hGqJqX2xBjDgK4osjibll2oDe+DJSle9l0RMQQmi
4EweicEVJkNGdEMada69nvh9ObRtxNx7GMyIpwulrjYqkIfK8dHSLox9VeEEj5md2+HH+Vah5xCD
l0A1/PspybJKvX7eoYvkVr1cGObkNB3f4VGHE9M04MKyD4YUv2iyOx0/mu0VPSGIdOw3synp+qVV
WP+rNtYGXIXZYwhZXJgSFI70zjCVjLtiwO1GoE6kbjhvYXOWyLM+B+REZwLMecSGd/FB3x6nf1Pq
Io6Eq+1rvXVr04Ml443P1kdXb03c+efPHnfkeQ5BobUssu860TyXalIQmL9vx25hQMbABKGkJzyN
CgdhhmflbZC93voR7cKwXRTgWHPnCdJBhGFk1mGa6+fgiKTMiBmJlRZAacVDZ7U55Ejj9h9pgtVY
W7xrvC0K11jse5OWDuOK0DaQGDt2op5nN/TpS4/fBLYWKD6+vNf6/zF/civxUreCmLQqT/fR5AcZ
trNQFlkzc8bhSMs+r9KMvQuHf3LOR7N7WhLOqra/k0H/sTIQLY4JUbax5RJZLjnNv5iHU3VTm9rZ
JS0ICTo0oBMN0FQ+AJIZjMsvIyuOBpZmrPsygbRy2d7XUbtjLb4osLSe71B4dKoTxj2xpZHV7RTr
y1HYnIyRXsygrH2Rx+M0bToNYT4Ag9g7a8HPIY9rCDDsY9YBtUN2ZIhcIglvFYENQGmBCctF5zWR
e6kstHx4tZH1cjTcnI4JPzFH8SwNefObXqlmZ5sPO4qwaYCHp0uxLbRTOvTxyB3g2udP8H/mJZYd
KJlB3CZk/1Bf5gGCssYeirWnCkYE9BGEEjYqbS/IrQPKgBOuPsN2zClyXJcCRLIhZAhuNItxN6q5
GBQDtS3rEVr0ZCi0cPcpPFOTzNLlGcGfhhgdSLAs7D/HawZNmXyjxLh0cG/f0eAMbcn9AeI6L0XX
dugfllHIG+WjmfkDoSboQfHo/ZZOZtH7T+lCIzTCa5pPeL6ljq4KRKi1ePmX9Hmax4mC2uxndSHO
BW45wKKIHKrce47b+W/a8m4C40iBnSc3ydYlUEh3fhwDIouIRnAnAIYCtZJ9VQbeiQ4VJXDPC0bd
aO5WFFE6LAO+e3VuXWgN9PBup0wyoapLJv3jPlwkVFyEEUupn4rfpWU6STTUoeU+PsBf6ZENOuhr
cKwTJfhDipS07q2A4KbDruYh/snx6gyvsJaw/mBqwiQwbflIVU8a0A7YY9PV0ZHtp0/7tGcXUK3+
evvt74W9b6Medj2EwMH/21/cVa/uN8svPJf7/fqHY1yEMgbZwWdzB/Xqz9cNbdHg3UwkJ2n9VJQ1
FsIw/PmHlcndbI9lT2t1JC552hoUktWN84+wQxh+54K3aMO4hzn3+XwMFN89y69DMSiCKOsCkCPc
6TBJUiJ8jNOvBY9UVetvWq/kW8+156Ixgc8A9PtilQug9i3+02GZPMoQ2NapDhWPdUJ/X9UC0A87
ARTSJ4hIWvKzbRVQJxOZL7IRrubNXmPOYS2NioozKb0TZea2p5SPmAh5ErgZNsRVuqs2vv3h6a8S
jKDhIHOTExO5pqf6tV0FHIwrcVi6SiKrn4BlP4oHTqV50dW1Quee6CQrZwxgMYY74lqG6egsSNMj
d/1+Oop5hR/fsO9wGDdJaooaABV1hbtPpP5x/VCgeBPZhiC1vDT9qZk1Vlhk32JcTFx2gwapCQUV
4AS3uPq84Aj/R8GZxNBjQuRUw3n3O8zqsGXndCgJWAr0SFdWbkqg6eGSYnmAJ9nW9gC1KihoByB+
taOFbJr4n/puADD013nWRGGhWNufOzvnTAHRf920EAB3PCmpm6CGtfcoSFRj6tsgiGNvuTLuaebc
Ys4pCnpA0bZ4e2Li7m3hSdrs33XqZ91ksYpik792prO0gldbv36H25x6NAbVlU0pQ458tInBTwfR
fFbyH1naCFrr9SuisrUcZHhfUKHtIaaCpLbEjv72hG9SOfwmmjOM/JUnsOcTzw/ore1ETfK7mBDa
7d7qLvrKeC0zlQFN92RcvCtRgf0yqUL3G/gwiMqTC3L3tRJ7ae5h1XGvIXcNr1CDyLMiVW1QHo+f
3SZuNjLpx6tqvNzALk0zzeG64+lEBP/XQtZCgNo/Cjvo7GwE2JgCWgTWh2MBJILTdmFKP4r/po6C
zIwjZ1CasjYci4OldjOAH/RjMYyZ2rGv2jJ2cw/+w+OJNml4QdzUw3ugY7iX1E2F3ACk/eu+GHr6
w9qCh3+Srmyh4PTzGSW6TupDBLNuRRh3Pw4Pu3aMtAb3hF0OIq2DTPcxC28Ogm31APdnbID2i6kU
3mVGomFHxEJklTBoHF+HWA9N3NMQkTF6/DmW05x/wIr1A2Sw9Ij/tRMo0n6hXNjUYEyfpLo/jES1
GPbrTxKk5c62bNrkWHyg979ryJxk/94XG0NirvdSn0xKvoV+Qyv9xigvNhRY6qAcplkyeNYa4DPL
4T5ShkAR0ukfz7qHWnmr1YvRijP6Q4H89+77WamcRPN7uGBKT2N13MkdCPRKsJXZDcUaLlUuglHd
TYSfRTLxQAFkNDAknoLdWrFegMSTOQT8P4oY7edX2f7YK2qVZgDo+jSn4Ooy4mdBLcb/qloK3Uz/
5Umf2IcTP04O5GpHPgbLgudMHW+jQaVMFKWki5twXixf47x3hdBq7UHlCYohAVQ7Uh1L14GML8wM
vNS1N6TOten0vVVS1ctsgCvUdsFaEWuWrqriHLlb+waDFMefEgJSvZkg00sz+dJ1v7CyRyGQCE1x
kiVzsdTdxNg2/duISKEewNhsGAydxtk/1GUuP0cy8p6jWSNqGwnvMnhlVVtfRV6PDcv7c/UGF48s
4uOPQYTTBwM5g9rYcPMP76Mq26X29U2re9X/993bJOY1hKb2BmDxraIMWtTDPd4J2iLz0LZn5nfZ
1hOd7IO79J+PIxZzFfg6ygbjkSYn/cPwvxQ+OAHgNMtR23tnyg0IkgeZQcUfx9Nh3gIaRW/By5fz
Hbf+dgCpsP5hmcvFu8uxeUyZyZpF1k90HPLTED50VHvJ63zDtWtdOAA/PMsN6BukeTTF96TgxfHI
J+Vah7NsEfbH4e6aWHkF0B1WUGwFdmkzbc3HnseADNNDV0OgPhJfHS+yyTNIZxylGW3fqq0rUHcg
RrHgSCGWq94WrqyQdPeZqWVtBH7a0bKHTCXoOWeTEDN3WYGvR0ZRHaeS7gfdDUTcgSK72GQU4oRS
TCRvw4NsfWWy2fRJoEPmj+M1xtgITMsxCIQ6fe1JfkqjLhFzZCrVizMDgC1xrUEVpgl6ynj1CiVE
ojDYdwPq0oIdAlfbW5QSYjoXkKySrnOien6VTKm9MRpB87e7ko8opdz1jajWXxAmjX6gme5Gh2W2
8lg9GGS74bMTEB8Dk5Szh7WcviTfmvmXH3A80iADb9ZSv+vSWKgc/aL9wMbKDIbCMv4pN0OTYLPo
ilCr9KlAlYAgdF1Kt+WnWAm8DDxSotD4gKKMj7+MmioYdHNLTomwH6r6R6dvf6cSfTRzG69zhmNC
Iy6pNTt5vQJEMFWUzV6Yl6MFaeOP2n2xr+b4tmvftDO99cfKaLrs077ibw/OYGyeR2aeACggiF26
F5RF5C44KjAiDPvQWFgVtQFx0MWsw1Nw9caXVuKvk7SOpVgUgrCY0/e2maWTdBD2q8SVEmYujwcm
g6A4P1Jw862kg7z18NI618crW2c/CMcT/2qoY1WQUB+Wkilfvv9xwiZj5vIojdx9AtvV6fkmQrSZ
EeyeLoOI1Thja8JKVQXzWDYDXOoJylKDDOR1J9Vo30bcsHYxL01KDjTPqQzsu/RV/O+EjYLWp/+1
5JF6aHzmluJ4vjDOediequDP5nx/98sVdj22a32mrq0oTRlbxX6YZN5fZfggeaEMSg+DlMbJ8rNm
DqkZ/XC7MJTormtQuw8CA8U7Z9WA1I5XfNqYEL4OYpcpu/8Md3eGC5xFUiVs6mSg6nckf9RfhrpH
PDgAP+V3v3o7UePcwQudJtPHrw1wySDJALR6jYpaSBopLKkiqZbI/IQ2eCBFh+w85N72ohbxZI84
ueVaYzmorbgZ1FMgKz5ktN1OQrouSvId9Bbs0MPthdJ0MOsXPVvJZsUzljlgyJqj9PJOWJd9FveV
F0wIPon2MGKq12EXAQmPe4GGg/89HOALwPsO16KqdAJsoMYbACJ70WPRG1pfCHJKc0fGz/DnvrrB
Agy6V+BCB1EoRe+ChGOfYNBRQEFt0tY82Z0543b/CKRceoJVAEnUfTmE8X/wPTAXGhsL9OYZICOz
RPpHDEkn8evgRxfknU6zs3mEY6iTlDPhrHUQ2uGsGNioEZ1vTan0dnQURA0BV0Mn29F/uMGqxyDy
KSXl6OcIdZ7yMQ2w0QwwgYRKqA1DuUhkR7DzbCTle772DGZtLqvclYQcBSbvvRRPmE3D4idjaOP0
6BqTScn9mt4bWHcOcgkC/m6juiqSeaUDPjVMQlNP2gaFZeMKejiZdNxOPVWtFIGD7vpjHWB1rzng
78pZwLs2iiTkI0WkIthnuDwNJlE+fSOgdf3cpayTkoMsZrP6uEkIDyfPASxj0Me2zSd+CoKrze8w
XvXyy0JXNxw0awsDbMYvwi5EqNcVjjHt3uvePNECfmNyALfDlEjCt2rlRRLZO/hlVYMHNCAojhH/
WXSGhBGH7XEtBAmMg3ihEYDSxcBa1L+IJ6MhSg8HhSo+6T9zxx3fj5S26EQ9RhjH6F7DKNsBZCD+
2F1qMwqkXhkzKGrWohsSm24kG0wEEJpiPoZich2MO0jAbtUu/zUM9+pzP5ZXfTkcUSN/9RPdibwF
xhkWrx7XC5dRAPkGouQZE+jZ32yLZE7LnsXgQg0rIu2jylUSTR0IPUvgBEEwk+eEiLA/CUMTmu+U
QE3NSrMAfWdpzDEoQCIYTrz/zU60zxrr92m6F/+kwJzWmNBTAnFIT3mfRG2aMClOJ/vwSPiDCcZD
dT8m0Brp5IChpsOK7RosNeKUM//I8aDzeCZw364cik67oq44urLl7g4TjKoIq0eNzbmKUkrlPvB+
WqIzgvuITz2w0QoCdg8ODrlDEyt6sBiP31DhSM6C3biVC5nxdH/worehqMvzyJsVx4qtYpsq3tQy
GTmrj6Sb0hhD2UEs+TbAkP1J7grpfYXcFL59VvA9K0ZfilUJpztpalMxKoGNTppNaUkJhkBx0iET
AOMwucD8oKJOjfUmMD4f8KMdVAHxE0zHWxgHxQdY8ke4w2EBwen3HpvkhUWqm+kbqFTR1GAeKOJi
25u05UxNj+IgVBqBPaUMeXA4YhDJPydowZgVCh3jKC0G650GF4vecXree7VXBmjgFq02hU2lDQCj
ACqG3f9KZ+mLY0vEjzUDG+uPW5oJS729pK4wvb8F8s2atthnDxxxE0nTLZgyBgB0vpXDluwN58uk
e5V9ndgGO0pZm/fnHFhuNjSAJgQoBSGUyQAMyfqEx5s4dReCZ/33TfIV9U9CFuVfPR3L8u/7BZk3
g1/LysoQ7M4vS1vOXhyCrCa5buvvChUthRX6vltugxdAcrbZm2rXquDKbpM49Iz+qfioPfj8X7Vv
5OfSRI0/PYH6vgKaAsA/fIKARyN0q6wKfqk/5cH6g3H/+eR+ySVEyRek9LnlbYe2oA2vkGCbBhZi
bZ/N4S8OQ+FSGbcR9Th65EMFBXFJIVRWs7HTs2Mk4J0Xd8JCihifgXMCToxKVTJ+apgDd48hQuya
TARh5j1I6TSr5wKuwbPpocfFX6wTHuWxL2URjVJwl85vLiNpfGreAtyYoFVYfrNNFy5DcG1F1ixc
eAQ0Lgac3qpDUzEqjuElYJFBwBwWkMtAUb4BCld93a0pDKYl7pSMWMhVd0tblqm6rk3t7rcU4ysG
nIYk65KQM2IS9XUHIfyf2fIqTb2JU53quAkjw8Z9pHZcknsVM8ldgz4ZpPDb4oX06M9HwoVbizuZ
h3ns9S7eIFsNQWvtBsj9lQ1hIixXCV6B2p4rSS6MeK8kmSf5AIuiq0f2ExJOeDXE04Ra7s3p7FMO
QSILxThW1gJ7BLtyBaNq37k+SM600kveFnNARU8nS00zmr5IiZsCR7wg74hrbZWkxds5LNX8BBRj
T1SrYCWOdRC5O71z75g39LlQ34CCVyR/vPg/rbENivLSg7iaOV0ZPO8ivj1MP4K9WUnWn71Y9voo
H7D56QZRCKFWEvPnwxY6nwf3BjuYNAbMmVpLQWW+rDK/xwa7B3tW0vKfS8AXuAEoUlWO7F6T4jIz
CN1doU7p8tz3qkb0uL4+jB9n1OlQUpWNsYf8EyZUse0M+0HLa3itR9KPsHvbAZXgEnJcEvF26XhB
NmnguCoe12BZm4fY7a5Ptfq6V5o/dQ1/5cKsPM6tzWNTeBwWe1QZHTKJqbLer9MmjnKFlfs34jma
Oh0Fc06MHXLmXAoijUjneg1ToYEPsaOQNman35B7frFfatLgRtTbN83pSr+SK7K+plXsmyRfLj1K
up/lYsMsq4lNZIPGQS3N5sMMvSGDQJbsFHtQf7wL4a6kwhf+dgjuT71a1yR0ONfxrgwUyXnGoWJt
N1nIWTFtYoag9ZpOF5A/7uFjt0yMoROKH38NRZLEftimoHHb9SO+pK8fJ7SxJ0uNcuKsBLe4SvNW
5DDcuq9uC3rKEZhSMD7HCbrpCWtqNmDgbcDGbAamXci257Zw7Vd1r1fZ0YZwoBJ7XGJ5Ac0rXs18
jiQTWVtwBJpxtQIkKLSMNnwuqt1+m10v6dIUJnZMZKM2htiUdad5TeoJA0JCw1z1MxmE5v6ObDmT
dg8Xzwmw2wyUgc83mZCR3BwDLau09/idoj93tVWgy4WEd84FQV2p5MnPCfznJAgaJD7EjhrZKCrl
LPDTlEteBgSbDYyNi6yUHXiTNh8Rh7lUwpDZRFGtARXcaxx+G1YGypbgFv+vMYMloQfDsvwKMOrI
Uu7YCDrc5PAyGBSW5kdcmm1uTNFViPonqL9TkA+6EK5REXjcWmZ1+YTicZMX6kEBTtCbyOBSzMr5
zay6ll8QzXLU79rWUrvbzCfUt084v7fIsTUSbLWqvhS6C/YRWdDRudsum59wAc5JZQsYv5l5ZCjy
1FaDzhj6zbe1obOQptF05E9Wuvke4cBpusiUkLtc5GEXsNzS76rkgMuCMno2EgT/rp7XegAIR7X/
HTC2CQkI0gAdim98OxrwGZfZmVphC7SLA9m4zRi35q3NoF0lvL+9yO1wF2QtiPqpXc/qdyQEY7qm
4H+rnjid7HHpyQexp2yhcwfbPMnUe2k70rcwpwj96RWz4DNar2H0L8tz0UO1VHFMXwqXi8HGStnn
lq7t2HjW1KbWIGyuzfwr8PiDZic9q0ygjYNW1E6+TZbyra3WoW5pKsnkV+qmCXi8z3DSjFqsLf4/
h2r/Qt6F45enAK//FTsSgLxV5whKN+/dMgTkOnAicHPes0pyuEC34GIKa+3QPYhOw4W3mKQZCz1B
20GHT0Da1KTEZ49guG/OByh4/GG1N3vtHzxGCfyhaFvggER9Aj9nGKxYPy6n1YdW6APaqmFQcvFd
Jp3VU/EI/84AoDcHoEi5j0sMUkGdRyRwqu9vkuxJ9WcoVcoW+H1dnTXFtcg9i4V7Dhe5X1O/AChJ
o2qlOHbCES2SkFopa8spS0EuRR3amGNJLJtR6+RqzuyET17qkZwRyM1VHpLK+ysH/q3yhOKAGlG1
tljgTKqzzwoAsER26une58tOB5Og6C+P3VDtRYs8jaNtn1iHCj4phHZI7ryX3MlNKGkpszZovFmR
fXKIqMXzmqxWUsveSyaPNCn3zWzpY5lHhOO3daKXsQaimuZ+F7iBGJPGXDChcxLIbmFi8h4YeEuF
EdlhTfStDBhe0u5EkH2yE7k8aNup1KXFhjhNmfOGPF65IwFhBhLPZhwIa4+CVhe62l2ulEnjjgJD
KDDpYRQ1ckgGgA7korzXUr7jQ0p4sTL4PrMOTqHjVkyasiZ3eM9UYfkQPdMDQXmmH+OdL9gIC8U7
NDmrqs2psHqh1sUjWeL5e/qXRRdfF6F/JJBQK6ZC1uPSVam5UllCndl7u5Ulz1pcMqDiVtzEi7js
mJ9U0GXYmEmNOgsxZAGSPaLxldSsNm0yjBjqNrutZdgQLTdzJdQ0KAt0pY3MZAHEmodPlfziSUTB
iBTPo5ZqGnQirGhg/0cnVnFs/ChvnjszQYuPwgMotGB7kyrLcg9pGHNfJYGCmSf17AKpP5Fuj/tR
h1IlGAm5z+UTlS2/CCRDZsX4Laug46I/hhVAZoCqtcSr80KvgtMzDQeUZy3aF0hu097+7S4Cuavz
isuToIBiZrC8iD9HSgElG+8kF00tZMevNsUF9k8AEE7SdBB/0kZpIQbR7T2A6wdKpEHxGmBqdETl
FSb6NXy9Vn9utvrPbb/x79pBHhpRWflA9S8UIrzgWT0oXM8PMCGTNTpbefXgZ5ue3rpOesP4za9E
c+YNzNocZLNeE2RZEhLA3R9ADrCasT5F+h0BawJz/jOh5hqtk4Jir/2wM51wg5ycfWSG3f7qyJ1G
Kunw4/ZRWRa17r+93+hdSaRso2FktqCeHUO5Z1Y/BSdDlDt4JE8I1QvlgrQOmNGGbgfzKEj+4yrN
6duGd99xWi+/ae9XkhdvXX46A0QiV2tzBImwQplJ7e2i3bUvnzwBw3oTtGCwk7qjlmuRGfEUZNwh
dEhbzoFcGcCja0lOh3/xcrXqW3+h9JRr5T8ys1jxZDp3Gkqeyqed46ua8k7Y3NFjFjWUIkugUng4
JRUwPv4UdJixgDs5arOGMmAkiX7zclJQonRBbLjtPPVNWMyc4B3xAA3g6ZAYhjfHyKc3vieZMKEi
qgGQgG2OspIa4xcYnKa82tdSlY7Gl20AVU3cyrPPVacQn3e+Fs7vcdaImGgG6QB9KP0qSMr21tQE
KNL5JShIrwFR9WXRP9OjFJs0iPVSm54nLt0sXyTqcxunrcwCILn2Tjkt82Z8lP+MK3H26U9Ndlyt
kXNtsCyPAfwNUs5p2c1/5FqXR+2t6c6T6wKu89Ve9DYHC4uQRwQCcpJXT0YAkCOjGUTycTrbgx1Y
9ayrxxEr+Zu+ul+UlgbUSyMmHL8ChP2xO9ZGGpLdH3tb9Lg2HRZNSERXqO9oR7VLjzTL4WNbaB+6
jSLtbshzpmjPPb5iJ//za0ms1oeyV6kCOfebhG0n4jZSWU794Ii34TK3sLVb/WC8yxaOwONroE+g
EXtqCZHDm8ZHPHrKwmNHxP4YMZWAA1cfErLAOCx3nyAyjvRMWnmjiYqfN02xrnno6wIl8+kQ4T9N
XAGV8jw+CX/gXlYP1jO0mT0wpMWzLotTetZaj5V3fKZEPbR+CEF7106JX0bf3Y+ppD0uPl/ubgNi
MRp2XYUNOyjRtH/fx4ErNEcKp5nkouvJqcsRXIdJeLLuCIFMr+lZPUYa+cl+V2GqCS5OC3aaI3F2
xcJf4YTNqnFY5AMTveS1FXghxeZN/YuC08x/S0aqaZAjIA16CAuWK+gmzIfPvApCl3vRQqw9qiVQ
CFMl7zaepjsf/ddA7Hp6F/wOfO/Hmtpbcaju94VrenbR2LUXAoN4EE5lislpdAV4ow5Nsq0ToH/R
FVJUkki8XJ7AV8bnNOo6py6U2cuKxhwUBKU5H4tyY0f15MfBTGwPF2hhcTFya4E4JbPyYJA9rPi0
oFP43ttejLcAQ6ICrNmm4vle9zV45ObumFjwU3hTXOLTPQ3sF1SGBV8ducrD6k8n/LlqNvJra3Qf
O+PMmOcpSYRevDXmMj6TF0lLSnyhDtJidFn0yAajPBeC6BbgcnGMAcblpCgsE7u/Vbm8PYzGP/Bu
34hZnBJEph+1lZh3VoIRN9UHIBO9gArhmS4IiLAP+C86dPNwF5y08Fl99yqCRT5/Xd+M4IGL1toZ
DXaH3vdQJtpHyvGhN9DXUOyiQr9KkOxofDmWlgZjwxymaUllqa2HnzsTcNq62gfyHUN/EvFtrxut
HaS4XP4+31bSmIO4pknhan17cHNlKEVjMww4+fiTGYA+w/lTHTQfD9UJ6cT4/fS5uxi1FT+Btegn
uoerFZdk+4J+y5DsslQQ0myUGVxVD/v8uwiAy7EPt8lsY67UcRqdngoLT1/An8XMfjalEjRwaWjt
MShy5Te5qVu+DNf2IfsYJLUd08YbaUaFuoQEPdIW+YUkX09XkOIpm8BwV5zYz3FqEsBHhtrOam9a
JQVfbg1ItR8u3bOK/KlzCK3YfoxYcfEMkuRtamYuBz1EDHTlykS5kIJE4M7lYH3lW7rLUXO/9mY7
IoQBqNI/P/vtIxA4Lh21kurTMFWtATMGH7tOWAa9jBVdm8P6Eu8ZDT2YjhBwU0pZW1+U4SKoXFXv
FcTC23SYmHwAvs45/YF2fWKOFJ1OCqAJlQrdh3fBSe6dNk6lrjP2YWwMdVTBexOe2Rdcb8ytbKcx
pFVu5uo/45ZF+FswykAZq/qfcEE3pO1z/T7JxUjs8pfKjq0IwQG/9cQShJOMbqUQXDwjlWkz57fX
WZzHlcf6BgUyITZtwLogXFlGefGfIAujjh2pbQV1iqMT+SU8T6dmjk9xTc3p0l999VjTdt8tvsnk
Ucm0LTDO24ZOJusnyOMZwxksQRs6zstrvN7ta/A37aeVqq3BXzMI7k7pJZUIfZNYS06vGd6Nryoc
57L/9GHXo6mrgoP5eYM01aAt9XtTwy3fHaThVSdrz3gUB8Cm9oCZQGfSgbgq+dHd6pXTVlemtETl
B+Gbuc1sBHrTrKZVmtNdE6V+2lT/j1YVypby2RqG6Wrd8w+LD8FclN4ouJJwd+jLv56LNBfBDTqR
FGGr7pIyG0N5PuZt04vj4Ie2zBYb3pjnmnufWGElM0QjJLWEna3GVq3FXgbGyvEaDgtVZWjRXf7h
Uw2AwkDGCX+ZUo7896EwRW2R3VLz7kE9rawiX3bIVFJnAKNsZ0jiHZuMP3fFXEO4qALzWShufDZ2
+90CDTV/LD5hhcvQKK2dz3zqmzSv8WyfHOzB+cfahqCENqEWavodEy7+vTWepCXArO0rM80fFspy
1rhsZbQI8RXMDHL8n2q7Lm/guTgTR8LkhzaLUWWycnS4/9J9o0X9aj4khViBnf6uP5RGv6/k7NW4
rBm9PJyEkwrpOjE2xU9UjSed7pDRh6QrJiJAJhpQv83qkXtoar93EIDKxiLhJ8tuPDt0ijdrhCeQ
qX5Se/Bm0ASlJ7C29n74xo4UJCvXvUDcIS2kPAzxu5Zs/ZGkEsmR/EwDctahzTewWBWPPDetl9Zo
geOrzrmaXFLqqLWUbd2eaapJCpA2Z0QhoDMQz6aQ3Tui8MVEqOl8htdb5RKQY8zteaUNofSfB3as
eYOjAuhdP6G9XYsWW0vGlRLKDUyFBqSPQ4pBojUC10UfxQBOQYE7IdF2+iRCoQbqX1COpzitjNtc
I47Pnr45jJJO4Dj9oUuKjIokqPd2BefTH7L2mATGmrGjrtjzzie+G3hG6/Omdq4/whpngIqbZWnq
t7Km3UfYLPHYzrmeBka6LBSHp94nSBUQYDiBW5+WP+etyYlSumHtlNmemaF7H3iYiKzPxUkTa559
buIbZu1e/8BzVxwM5XZONMFFtFdr7aAVzhWFjv1TXWSFKTsZIMtCXMn7Jw1G20iObxv0uSl5ow4H
7rh0TyE1QrR9a6Y5ebFVtoEkwYu/d63trq6UwEO95FguPxeT7yY7oovOgDl/gT8d6K5EMECVNmVT
VF6RNvFQP1SVHvTmhkGYdaTHE2ibxsXbgyn9PEfZ6/YiQ6aZFggmTt7pzRhltQ4K7ehLJIpW6j4R
xPzp8F665Y3OfNfiQcsa0NXOLlCVIahLITFfb+F4bG7R5herbp5My0rNZEvZWL3N4Ddt5TZL6mrM
JdNJtO8HYYJrqsKUIijweGWylu/e8zFlbC/f8saTmREP/dmPy6G4jm+qSbQDDUWU4Og9uHSwda3a
0rSfLTAm7FeX2FmVACgTCqM0D2EspiiLm2uqd4ULVYmjB5mCoh6KTjIDB/VPtjMKl8oeMU3mUwOV
xozrV7GgQiILhWeFMLgr909IOGuidBggqHeSYLOd682VDtUUIiGEcduDLAbOjpB7f1k1JqfFc0cp
OKRPJ7EHJvSlM1RN3aIztXIxHOvvd5E3d46vjKYFfNYF5uETnggsJ7K6x8knP+gwW7fyJ/UU0e4u
cRsXvbO5q2pfCqy1p/yqrUocVCHiGuFYl89HOaLHSTe1GmSMmYn7siLtTfGfYQioLQsVPhrbc3FD
O7l4gLu8BYNcwRP88OHrJnRTpDcZxKK0kM63w7MR5SPWjsZhFoV12Ko+j7b70v5H9ySVmbCUTnC9
jJ1b7wpsOxHk9dv0rOFygWzLYozfcKSiB6E23rMdr95hvOBWupnWY0rTDlZ6ahrxzGZ/9pNEfyWZ
ukbg4heTLBRSm5L+TqK6qqyE3Sk/Gr9UabaT+DaSWoev5a8tfJvSoELNmZYtcFgqTyO3z9ixhXuu
ahVXWszTSYdL3U1nu5tLm//STQUYUT7QzkdFlQ/2YyweIkJb+vud9sYnznBTdwDH8eFhBlgeoxHD
6UZHRs6osJpauL2WFuMovZ4bEGo98lLwktcffYnwwLO+UcqF0fr202DSt9XYHxMc02E6t7g51tE7
TxF2QnfOdeshgG+HgAQkQ8I/HYvRjBCQn/ugltSapVKK8WxIRX5aT9/Rs7y8Wmgh3Xtlrae1iIQg
yQ58SVKITsVVCF4EFqjQw7yzjeFQg/KpYCgUnQN1eDDFDnRSJq6ZTh86FEbJXM6Q1jfhKLAAWpqh
OqJygKmaAuf2Ejkp6tKSdQpIQAVOFaoAFlWRgQO53u6hLFP6B2H71uJFKDFIy4fNP+v+3ZpyPaR3
LnusxxJTEczlVzRhyBTN67R8R2Mlh+RI0hMbB8taX1wpwhuhFhvnU914mc0C4eBLrrbyNSUrBveG
Tw/QSeBXIwYYFk3ZhS00aJWnviEWR7dAs9jsFO8qb/gwxRSCbrZtMEcpWv4aePIj3vW3dSE89Hjv
fgDDU3NWB9qfAs6OrXNAJalN2C2gvxa2XusN09b+cMjJ/ydX23KKo8Ep0E5L3V5ajNLcJH9DR/gC
lwbDzYrn41ZwOEyEMHavEtSNOq+4KlhM9Jl3Wpc85mnbB0fv82Sw+P3Qgxo0Ux/hLdKUoMsAxocA
CG1Vzg3XFshPeow6u0XQVFvB+JcZJn8+duExaxbmwOnNvrTuf1yqhaLwR53M30IK0MAnTDENd7hV
kVnPb7ni8ImRlbAYcPdiAgtZSbC1btgJLqrwAsNaYJlH9lJlSorzb6Y2W82N4b99DLnZ8K0+gkw3
j+f4eGw82nj6Q4yYgFt4fUzIn9HSboqKVwWJxjd8nvflA96MVn1W2n9bGqRGBcUjRwSnPPdv/ak3
A6UTqDYHpLd+YtUNwq4LtLM6lBGFIlRksw1RORNpyfwC10rmNBhBDnJz1dRhKw5XA78ito2ZhKYM
YagH2WexK4cGLPOiZF8Zwz0SgCb1d5XEhkUbLfXUIOmSf2HkNrCVXEkFGNl0Fx1uQc20pNHAWw5x
w6Fk2NYxoE/DX9UshfoVHQ/oXYZdCdjSY95dkMhLukP4gohfRtN4po4XwHJN+3dXdvt/6xpk5U/m
ZwO7mmXyim52+NnSgaASFE4CzME+GTBTO0bi3iwOGDOiaSm/2T2S86kqQy2iAyA/S8TASzXk2JIw
ZHjeJGak0kFEt4As6rkjJFDuP+W+xOnede3zMLe3zhqU0FkW81k/riRRmXAr3JhttBbdtNm8eD44
D8sUgdqY9bHhXDYXyrcO8SNSGXrxCFTTI5k6lVPc78hmctFEwNJSToc1Q15zasywpsqwD/NKBk93
5KKCHkD03eDYlhzJJdn7LQ2Qk+g4M3wOLv55dgmFfElySG2i0kp2LHPylPe24imZqRI5EptdNCLt
4wdCR1KMVpHG4HiQLZ0u9yUKIiPNt5Foj+Nz8haRSUFek0EMXqcanYdWmOTUxY0iJXdkrHsx0CjV
MSpBIFMBngWQN0h9tFcqBRA0kiW/VeeEyEzqMkZf1jlUb80b4KVS1f2PDrMasTrnA6KXGnfRoD54
vFhaTK/N3qof8FrAPwYe65Y7oblglWBr/DBBVu90tRPR+cvpOeZXExfYXHizBNYL5EAQli1k3VCz
57xzizqQplXKuiuBHxTRtly2qd/MaejGORYAKMrBVZ430hoTck07i0mYYotXwxyhw7Vn99pkOPfD
W52TDs68flJ1RqPGzwi88nqvsoBG0MOHL4Q9ow1BhMhZc+KApCFW6AXPS/R+uNhFkfb/yBzVh9vj
Qacf3K4aV4s6qq4ong+cP1FvBFb4W6PQscKQVcY0G/pqTyAaK1hbMunQGr8KPJx8wCuQrRfhZxA0
5+aFUYTPiZejO4ykDlBz2lDk3CP+2NX4HTXdwo0aUkyAOe4nO5LhurBm67Sar7BXRqyoQvB+r0Hr
xsZAg6HMoSW0CviFykST+GtfNkG805QO4PkeJ/1BKt+LHuiYy0cVJYyD6fRqsiGWixmaRNA/fOsU
NJ0JNhPC7FXEJmI37RGXz0FSGPgxywKuVlm5w/9e9/ggnrW6HNF2y4k8RETapJq12+gwnO6V1lhL
/8kCx34m+yWDEnFzB8ZcS+mA4jX4JNKLUHwjE/rKmT5ORga7OTlW2X62R6FOgVGoftH8Fi0NC+O/
PvAsuxrKAAIf7m47JVI0eNb6tunOUoeReQYMv4AzezREV+Sr0vA7BAHdWvSco/IBehdM0kKJu0ln
sIGO5j2mlh/7zZpfHOwy16/cxMTycHEkh2nnT8ygOmrKVP0cAptBXw/UwPC451JOGJ/DDICIAfr8
xSRTIGdwILWDCsA9FdYKU1OMKptPSeSLahcv7tunV68Z/X+/DEbSVA0TIb2Viy2Skq+OLZsrhufs
cLZyRZM9Peo8I8DEheyAZvqGBbdxKkBkhfg+s3EvkfliothbNL+8R8OPAkz0kRN4j/2wysONtSsN
q6yAs/aFJjBhcNilB5+8YFLCuluBSfWo4x1BqjgDVMwrLD1+M9bXEbnKxPsllS+oaa+TB+pyNzgT
p8zfLatY9WHIN7la5/s7kaxcqVCANdnHNynVfzSJyvKb5qj53MSGzLU1rdb91OC+izqh4ehGqnBm
J59r5D1CZ83FBX7ZMul7xV1RMGN/zfsdk42BI9w28IRM1xrFKL2FjaOymKdxglWeGXEMquzBm0Si
dwNMCl/QhHBPvtIDaGa22Kx5+ncPUrATLxQmfCWzX7ljiZW9p1iSFxGg1uSbrywDX5PhmWT0C7tY
wuLXGvE/6P+uGgXMUqqMO0ikMi8Mzah8jgi4oYRfu1GYSmT9ySMALXv4zPaD/BMIZzaAcFDz4Nzn
vkT2oC66v4rFK//MdE7He9tnVgZL/biIsT0DYPnflp5YxDK8xCwQaoNZHeL4CckkJgwOD0jyXP6n
Kq5/70RjG8YwYX8jlo4n0HpcV+FMXijh2awJvWS+iQRFW0crza0G+atLNd00Drw/KPyQIE3fzKwK
Bh+sXGAI8IPUwcSumHQySGnEDAt7EzXwUXqlsqV5QREoLlW6Rbh/PVRzRC6it8evfVYyZ5IpQyk+
fuhQCHIuBP4qLOqBnu2qS1NVAawTso+68ChuwK/J3GZUIJWr7JHOmTppBFmKkrdu/HW8Ni+maONz
Il1DZKNSB5Gbb00DPOOuaV+Fj0ZrOSqCRbXntieImZllHX0ZJP3eZgKTw8fgEYLGXsSuGPLxqUdS
dScuX1q8q99s7P4qUIQcIrtTKzYcz7z3NZDFNBPm0sjB0RMYpt4LEKDBDkqS6fySdt5i3krg4zJf
V0xStWnK21+fNQx5I/bN5LHe/ejtK8fD9bC8RftR1/wx6x0omupmTVH5BF/mIew+QQJklX3AhEYl
nY4WSFZTfdtwE5UnZW9sc88oESZAHwJBK/7M80Smo3cznAeIC9PN5WNkBsDrL7GKvTuS0srGZTcY
jdCgn6zZ/Oq0LUWOzw8dsZjcooTA0kGVOrkwmNxfj7BBTc6lvHqtVB8qrsZq7Z3yOkTcjLcQU/Jz
KDb7yk9P0XDSVNRnv+C/eYRndpU3VWxAiju77lq2YiDc3YdkPq0ZYGsczMqyfvPmKJPv/EZqaQeG
WnHWx7paPuMW9sFVVffG86N3O917OT2BGLsAJUPDDnTmLcYMafjjiFi4Ew3tVoqO6z/gIPZ7idVp
FxueXPa3FF2IjcNtqOeUOdLNfm1KxG3t3B39zlLSehqmp913xo9DW5h9wzZVwVnJ6rZZEjKEyiDZ
p12SuRsHw3yWz8/WJBH2k6AK9hB4dMYxYMgaJmtPwLNttUOjP/tw285dqt4uC+r0kP7lslfnn+pQ
G5rZh2fXdC9eV7ssY+//dexzCNIuBB19dOBMJLZBjmEgHRA+WirNhU8zVPq0DfsaukcHEmHBRokX
apjQbCEABdNNbJER6ambBcntOGVfI9QOO3tVUY/4KgdhkhNf5kF5ziNvNBnPwYo48mX9+cAnfOrA
xrq1nF15Re4/l0o4yYv9nMc2gsTBiMSJTfGayDvr3Rzou+8vogyFv/6F+FAqzNA7DkcQ7ASY/Q8Y
8wselgc5leRUX+YDLVMhPBYg0RzxYKD4rJ9mWvZsC1/b9eZF8GEUnxTkRTOTklQ1FuI7eFsIstot
3uhkuZdKn7vQD9MwLtpJcaf+K3PNAKOoxsP9IxOVbwBbMutdRCrJ3CjMdZP1FnHQ7GbHcvKG6GBt
h4ZiymnDpFBvDWJGYGolwh4cdRmr934l19OQiO5l/B85n3sv/o167f+7DrZP/KUVf8GcHV4e1UYq
G45ZUNShHHu+XXL6EQMgAU7s068iqPHWfZ/b3IrdEbFUdP5F/lWAEhPz1VIbTRB3xQOFTq4uOUkH
kEGqGTSiQM6+Z+Tb6ZuZ5pGU8WLXeY2e+HB3EsTF/JhEoxTb4kKpcOtj7Jeu4/77oslZIg/VLSf0
g48INcRqyaExYH8RXvy+MUad5uOiv9l18lFlRYxrdhABvDwPylCuo7tH5/25EzZgOF1JRe7OrALL
5lyuLv3P7sgfYB+vrkOJgN1bYfjZAfGyISt637QUTiyIt6EkiSYTfRQDpC7PMp1uwRrY9UEffQnR
/rJVUDVXtdqon9lw3pLqYOYY7oqTcERRDWwxi7kzMajpLP4eaXRaZbAYS/HurGaoYk1NuuDzLqmv
5cioGgzEEOgVnMgyJC3metaCJvkZa64FefT5Ifoq7Jbvodbjbz2d0ghjn6PX20ZsJd/DMWfzZ/q3
gHc9Pqibu+FFEkU6qCMRPYpFe73h94KdaiT+oJPUcUbKmCupwwTtkLQ+ithh24dnUa4vqLwbAcKJ
pDymlec3TovoXsbVJFodXlkrFlJasr4kt6npWzTux5TrsEyobrHoNWJuNbqP7CcKtF/Var084Mu3
u97NDJCklWGomD90oHt5dM2v3sDo61j/B+4LJvbxl3gMulZC3Wu7wWwMGwxSsMryBD/fgr3JZaAA
gINmc6a3LCf7BmWyXl8L5pZ72T6yuFPM2MymOGdpVpwE/bVCBnriXDK5c031klOHst6ti6tn8cPl
YfAipLSyUGndRR40S7vlLiwKqP6+DkHlgLzisjIx0BcGGyJVmwYgpWJDhpUkcogzUPTwBCwWGgeE
rk1xxaITGI7yDYXGp/K25vy14sSf+cMxUDDBW0ZgTBehlDUhK7Vx+VaGpKxDbA5/2IYzh6Z7wVu1
eeAJXfIRz9C2oeKla8O10tXHp9LR3X2w8SSjuNO5EoT2IjHga84ZCKr1qbALor8nQdY6rTcQlYHI
So+mKrPhb3pBWPfk9nLGStzs5ind9MyWWtIMSfrhF80AYMFwsLXL+Dl9k5eqP1yoabXs9oqlResB
TxCHDc5tWSUAWAXiBLSecxFSWKHMsXp7rpgwFt2ZQGHUcUtjWh/PCPpzsaTnW97XBQbvSI3K++3v
gL9D6wivrSUw6tFJlYIrppHMumLJ5Hr2R2WmbbzlgJcXo5fsHWVfua78+kEvrzy9qhpD7Gra61Hy
4kJYT2DUGVEjmfhaT8YPLce43WU2dMyMpGhbl1dP/nZ3KGO3BcHIbwiQX4GAmHsLhlBQLeND5Ju5
eSOtTd1geWYmD4xWIMr9VtR5p+sOaPis9/P0ONUMwFoTHylNrb5k9luJ9LpIkb2577Hf2ehYpmzd
0RoKlfEPbIhYYOKq/o8ync/gqyRwgaWMdiQ7Bvg2aiAe0ov9fNe8ZJXC5i+kPObxKjw5YbVGC8Wf
/nvJVoTxHHpzy7G/xvhRSNl9rPbnqJK0pCoXTqQcfZnk8ny+7CaGcq5/A+fwv76SWYYIdjvVgOv6
jFWqA6eNH+X6EzKnpTIzmkYEHCDEU9Wgdxgp12X1B53aaJJRE/zoW9/goKy8eBBakJHoMcy0XAvU
BKGX2qtkKyZkUueQaEZi8/0qZqMEEv39egAOH0nQERRFtgxoc2d/JAjOq7fl+Qg57jO5DVyfzhcK
6GGCUJ0CMzouwbPmg5DldHKdSyzCWik1gsFHRCl2olroJCjHVxqRpCVpeEzlAF+9SSOAOd+NGmtM
pGOTJwSHD2RXI6K24EJ8j3He3M+Hrit0lCDlnsBMbn8LQlZmokHfUbtPXBlFnDn/iDFGLZYDdhwV
Zw8XwxvaoT7NLjoInvwiG9YZOHvp4tu5V3wkJUcgAqx7ImfwjFnC46pW3906YOzUv1ohHRL6x+M4
UudcV3F6ixxqzFfeL9EzKnfwylY4Cwmc8gpD3sBlEVUBZLh/Z3JIDDjZ34fRxqQQvX15748Nf4/K
GV9fwbiZHDWtzV+fvwsmWKqgaicBGfrDHGBqK2exteh0vtuYJQGtMyr+NIpD0A0mrMu/eHj+AvDK
Ql8zh9WI58KJpqdNF0yGGHbsaRw8kQfkFc98QylpwVrfN2gk2TiTw1TOvTQCeyl+xPWSHgtYgKqL
NcILpanxJpKLrVXCfp+Wx2JTlHuJ3SFY+I9ODmbWw2KP0xGOfKdUEePkDcYsxax9uDHb3Ew6Qy7X
DNaySaOXjrlKuX5EXICey2/LSIGNczQhya4cqgxzzqmh9+G3LImjBYOBb3xKZglgEY8eLxmIpRXc
XYEwLCMLp+IRP88r0PGAGJNxhL13tVNn9Xt0gXl6yu6SRJRhoaohiyCG0OZSWXdMEIHe0kuageFL
6tr7RfOJOULDNaKySPbgvtM9dTFQZcIux1dXP9oQqOzjxTJGJw1xO/h5g0DELGgpQp9twbuoc4F9
If4Uz6oyGQEMOLyPYb3fCu85QYL+0JcbgC2AhRmboHzj6JmG1GI6XKb25DDzXBKkzHxT6pzHRiJI
dOyVDsC2NKmppqo3CZMZkMBqko6Xw2gkPXp5WqKOhdtm8bpuFRCgrd086QBoBePJ/wTCLxjik53W
sKzP0s8maJ5iLFeEGVIijf3WdvNTPfNySDyuI07yykEXHh9IQXOr/AD5gu3c4LDc5cPqXkTJougn
prqHBrlY3va629RlFikE4kzk5XL8NXN46+YAuQP2sZ3rU0m4w/JQckjSB7SXkyW4l2CjqvCjM+mz
0aQjCXWDkELbEhPrzNWmE8i74eC30x44OfSJqJKD4XckEx0XzPY+v69KXNFCIk2FIPiHKOCXib5m
FuO3IwZWr7pQEyKNFCTW4W7H0szi21uvdyYLxEzBr+7FgqOKheIe+HInZgf/PWIXLy2Nqf87dN7/
0bDL0E7KUKyokF9OPYM+JCpYQbgYpbXtDQ/TvXZOU3JPXOehFks/JZ6o7xeyG2F7HcdsdVnZ3Q2y
6L6J6ODS/yDBvMVEi1mbzkviUjloo3czr28ng6SLPZnpMLSPXwOLC7btnPOnTPHlllq0Zgy3oxYE
HKWrBnyNBuikDEGW6jS4y8tQuayQtl308OlFnQX1bZ64BGKNVcIkxo+Xi1WOUKVkDs0Vu1R46aIw
Rr8307YsoXfj2ADDEixkWXTtcLH+rdPu+6+VFhR8vqpm5iqnAoUg7t4JH4V340UlRx/K3yQdpc9M
X9XtOHaDug+4yp7bt1bxWfdBRhV6qNwTBB6YlFT2EchqDkTZV45H8DkoB9+VwkdbOWF2mPLuHBee
2yVP89vTtM8m0kq9pQqs4cXJ52uUf5gtT4KifCVguLvLRco75kPEKjIDBWR03SYfi+EzVd735TjE
S1V/QlCwy7qkXep/f3w+LI8W6dQmBtmdVTN2IpRv3FYorcSbElnX7e05GHwIoUyUWYmkPl+B6so9
aKD7Y3dhzfFw+3Vuh9vDHpCHf/HaIuBrjsDgCfxUK5HlRkwAyYZQUQAwJX77EjoptPw4H+1V55y3
Aj44UCZBkf2oq1YRgB0NMEM195XkODL0pYuM5iP9zlTc7dz4Ly/7LnPFA31SSHq7+OChgAQooW3n
mMUC0tDp5t+LSo2YSJFCZlZD+rCnUg5r2ggBG56JnmIjZdjAMIwJTQgEzBx6wa133tBptNTZmGBt
aG5Nc5OjOkUjnxEnB0qjugSVRaqKgERiJ6LIa80hvBmDjaVzvIqXeOxRBeeADq/8oc94q8AMpP0l
9Pf3KwTHAOLoUN4RB/zgdSKlIOBTsj6teDukVOWB9ixtOO2uPnyVBXdH7JVJlJBMYdXOGog6sClQ
6+2ciELw2jAn84lqSF5ARFiippqxh6uQsE2mgBnwno77JQT1MYGKHkgzo/rK8AssO/aNLF5yBlJx
XD0dzb17ZQJZKh7Pq3Vd5EFj539oz5n+y3rh+VVeKaxSXmUOzMdI7izBN61g4mNTT/L7pHB8tUvd
4B9hZ3ohTRQG3uJ3ubeStq+O6Op91xXLNMy0LOO1eO1YPPw18svEoCim8+1748cOgNmKc/G3rzIR
vAqn3P6uCCOKvm/n+bnFYLI6sUhGcUa/ZLzDqHRC7x8wLH6nMl0YRPBdJ2bKQRXkJ13Xkd0/gZXN
GYyj9makpI07QPbyyL9p5tC5Vy/9GAkUpkYQXmExtBwNSof1UM2gCBUdV4ZW+dx0+ylzSHOFrFIR
9qeG7skHwf2OfhqDcS+r1tViAKdweV+RfX1Fb+3GDtLOI0yj3xaFgGkXMGDoPsEr4JA/TD6/ExWW
+E6/p6BZx8q0FanvlX7ZlTuU8Z7ayIz6YGSNFdwXBB3hBZ9IAgwAs+sR9RlFi3axZiDQl73TtY+T
//BALlZfHtM+0bV9ntrAtm7daPIy2ir6h/d7gEiTaOKUZamu/pd657Xd9v+xk7/soTlmi4kHci9i
XkFYDHimIse7InhI+sweO7AOqybSNcnL0USiKJ3JQOHq5ZVHRU5qKBN90K8DbFLJMLVI/wBSLqHR
JqA+GuQ5paxsaCb9ZCYqEU3Txo29P2NzWwSoUG5WFSGOBvmTdUDKivu3fcJjp+lMM5G+PMfFPObH
wbZAZWssiHjyc/T7B4o+jVKGSmcs7wKhOspwN/H0D2TsAAEV8h0LcXl8KsQ7ItjNLcTZXh5K3N3g
gPI3rXAfadcqcaeu1/FNkcphBdq8R8DTqNbDSbzPeE5jTjj/QCJpavG6F9PVDhhq80MrTkb601KA
Rho4OvBMkXx1tB1BOFDO8QQpADKTpLD3nrOvrSqDnTTOCBQmoNQLr2DHZV5KWRLxCO4EC644UIH+
mfEZ14AIJzqYAepHt8oHwfMXYZG7K4sg1IqdDPlofTgarBFvEoM2sDKi967fJNJUgsJ65KQR136Q
DgmnE3nOekhIPEMxopE4XgZHP5QHAv5T/BMcplGtv03iJ406/EfEGFhoo/fuMdVMr8CEmUFRhY67
8HfZnV1R+mUGAwgI4n2QLTe7tZiehAWtYuOgfr31IFUCVV73NvjB4EQeFLrNSqL0G09ZWmVSFTIQ
k0sRaHdvGyQKGGkh07YVTdYeN3jwjgBAdRpuxCf4BF8mnhJ2vFK7lri5dCiTBqtRVZeIPkF0b3xK
ry4CmItjzluJm/8ee6FkqvlCN+qQT3GCYNauIgIh2gEYZy9iEIfED4jXFkHRO0VwQfsGR5MIKOHv
jGNQ0CaC1tSPjAW1Qr815feqQkG/TBvN1KePR7PK6b3HpYa2lepCokwewpsxkCsHQMjUwg+6KX0t
oLPQ7iKYGX3/weCVaeWFPoNBVWT2vlUqMwcloWP6AZz41qxbz/H/BY639ix4S8YxRZIUDQf4A3Ih
tUyRIj3t2NLcpKGhk90eTWMpn0Du9LEkij5o6GhXspDT6ouMReEuHOm4VNrbrC0KiH+n2OyDZ052
3DybFJ51u63WTVEi2gv/pAmk6ClIHDXg201QvaZv5T/q8CE1E59NMPh9sSANrsN3HZ1L2EIIMtEx
f0PfNhrrg/YigLx+imAj2KzcqTY4pZQhrhefZTbSq+EfF/gcLMuTPBzvk7ysyT3qhLmZcI4lIAdV
tVcqNnCyogDyjk3uOWcU8GZxzGja5IU3+vQyyOoF1ze2Y1Vqe6KXpYt2aCBaICn7tqceXANgqLT2
uES9zjZAUCjy5196Kt9L/eTAeL+3LT0HD/6wgJewtsGLYC4as+PScl62uVXXboQBf+AsG75TS/Fa
t/EHfharXeBEANbBcuUcvYxKkzqV/Ue2WsvhcbAZ/7id6yUSQKM225XwyQfcyw19M7zxUub/aoDI
1Srdw6qmKigXnh018iK1XO6uXZOH9FqV4Q1LstwQCLOAhmUkFFUi7bUyCoecrX1AmzUoHLRyFZS6
SbQp4chza9kUKmAmVJsPWUx5kzq93ckMaR6jUYQTBpb/O0LDKnZI8ZTL4yWaeqHA3FjlBlVgx46Y
0mIlcwVX2dk0XWsEpbJV2zpUMoYOmurDniZpQcy2iDwvXfO+mhC+be2iQVxSXL2jPG50nIDJcAZX
wjEWLm9IZ9f9xiuE/kCOsgfLb500u/Y9nIwk8Qo7q6x9Ei72C7I8OUY4R+8W9IYfCP7qeUocyeJy
+RvTHimUj7NTM+wGVlDf0eRf2zPWPBT0oJFMUFOXOO2vGkHPv2dEyrEZPg7xESKT3ffiowIZMDQ8
Cpfvu42vA2acNpDimAUdVnAbvVwvS26ld9nxS+7y4BJZyI1I6O8DO8y9IJ73IIwxoOL5yqHVikE7
DUt+cmvEkL2aK8VyvY6rsk49IDeqVzWF3wHsOofOTdFJnfIfYcr/NgmxU9jCFgqw7DH9npXMTY6C
Cpy1sL/9kcPHtFBOHykF7LPsHdMVQrZ3qknt7eaTiisA+fhXh94JndgTGyF/vnXVQn4NVRcI6ipn
VMH0Ucf1PhAsBettV5GUIN2tYg6nF9MuIsTJncxXLQhi7l/8ApOewroI0wA04xiWUOgW1cKuv8kT
zMvbjXhFL6yk88L6xth91Rv8wvcJ5+cPqG2VpOqwHez9KlX5gl8fHsn0uWSX6iXr7VHk7vizQfbz
2cz/o8kxtfFMcI3MWgUtKrVMQ2a98+tmaopbBYJIpRmgRI38VU9d+glMloTqwExWxhTXc8aCILND
5ZwTsFtUkwO2cmo0LPonpQq2v2koS9Nm23Pu6oMFXWP68EhZQ8iSzJwbM5qvnUcdHvGJZK3MzC8x
8UNaL1jyG7OPn+QJZcYhKWKVtmvCQLBFad7AGXjec1Iq+y1pZltCl0P0Rlnx1Yt+IJc0Gb8Z0FLQ
HHAAuAUX0NxENkYyDrn3BKbc48lieN/EISmpXnIl/YSV63PLnxONS/drR215osX1kf05FtcKKef+
6pGteBiVxF0Dd2TOK+y4pl0XNGKBCQKXnd0HiiXwahrx94rT+jl2xAUpFd6seLn57oya+eDN8D2V
Cl93yjcWGqYx/Lc/l3UedtYzXLPndKv1qI8DhrtO9DowtUmSz7Dddvzboda+EIL18S02dZqCB8Eb
mL2i6Ul/tI+W/emLkRbICfZc2IL5nYMAH7ppg7CunnR09ciQ7VSwdByQrGTt2wp9wqtOPKqjX+vY
offfUMzaPe7/y8ALMVItR6mlrYEz/hkEzWaJmQdf5OangvsQOlUmzbSGUwPoBa9G8LKC/Nwifw94
sIyTlwGEFsFX8aR4D8RgcXegN21cq73qTy+tZYY/1m4zGvVyvwkw8PQ+mj+JqUV6QSTYkTOeLCTZ
Ym42BKIPAt5wtOTcL2Xy4/zVOUM8N1kyw0w7obCbOssDHM30uv1vUfuHAoXXKo9+jBhLxAlOxNnJ
CWr+ZzCJuNea1YOiiEBuONdI1ln5o1KHc4Q5d8jbY/VTOm7f9LNBtBP4dMlu/whj5mzhCPs21TbL
CPhnBXT4/58ZIZIaqJuLfigL19GN/jm3RTlAYgEWr2f7GfNoNZAkt7DMSSYNMlT1l8oFKB7B9Qz3
C2g77l0NAwnUIaGVg/fUs44vu7dOe6LjDc4YJfJfGTEOfKlzherJePC7abtosTGWjCXm+9ltzFTf
j3fOn61Yfxup/ZT90cbDeqC2WPXFuGyI4W7MgTWyOkwIAjv1DL/TZnOaRhXKAugJ0/Npz9bilBOm
ghxaAE03PuNiRMcj1lhJmdNGaJE4IF20IM+gJLwLlWmBdZebZbXBn/V7CKYzeDB9wmb/IgcKS42s
/VbUir2VSluSOTgr5VNphW2Ax9eRk78e473FTvOj5iZ7bN6djNp2kNCIPYtAxJbVEfIqlzoXkyoH
Nf36/xDqFyUm3VckKByVvjWRKjlRkC7QMBiK+wGhYL1fgXCc8ZmNBNwSpd0TNy39lXYb/LQbb9O3
AL5b6iK9+oaDUDLGSsCEKD6xYoglu/PcLr9ZDHbRCoxUrTosAR6mItAgbTmLPE/HhBwC7Tu60WYE
+FZ8y2ewCs+P9+ruCsOiV7X2X3zYGPAWFGxlWFuTuUwVYG+EmjW+cGk20mnO93y2pOhDXFPTP2Gg
t3NEjH+AVBb1CrLOb3GOo751BuP6JkLAHIXlYbalXLRV8+ypr0wrdxIgyGkFRMV1B8i3sTqEJHyV
oMnE4eRnrAqWlE4vwt/LhxKtx2qkAHGgAZW4vYWVWUEhO6KY8mzLVjub36zDvvP3s4maMF3Ec0FW
Sp/SP+TDn5tOcs/jzBYIx8ZEF6ZqSC1+HCJ3Dkf9mq3SQeyjD2dtMZO6yHiAP9rhjpIMCwgWXzzi
zGAHoVc3+Ul9FqoWblXA1ud+8XjeRZLLZbHcM9k7d2k1L3FqAqk9kaXeQXuV+U6HuwQs3hKxpnyh
peY6uQLHpSwgb9YYp0jHViDi57WBuGjIvON1KwFlXMKPJytyLrk3CISwU/145ppc7ayihaQM3J1V
DDkP7+Z1RD6haQbfXJrX+30iajWpxO9iFBEZje9ieBmbfgsV9Ntq7OdS1DRwiJ4mv4SWW6XPId4E
BX/TcAT+P0tn4S+AbM7WM/yT5I9/iJAk5oWPZFtxeLfz0R3AGeBTspeiu7c1rJ4jCxikdr92yXwy
6U95IxAHLa9GqFK19r+BINKFG9556GgIm11nmJTLpaGXHoTtqupkjKKBCCQehP/tq/1598OYP6dQ
Nf6ijL/prOD127WzGorHql7/thMF1hU29HD/aWcEkbdml643Sem19UEaYi7cuD4BkycGbzOzs2H6
bWcYflUsv3CqyS7LZytR7FcgHs/wyf/+8w+XmS4fPz9Q85B828drj2yvQc1uY48RRdV2wONDcpH+
IIJ9evVAvkalk/OqsbACI7MIUBuop7U14A4vToV7b2zt7/P9y0J0f8SNIcOR/6YFglyibi5bWSCr
KL7BXylsyRMYCSupUAzT/rsV/q4V3wakgaOQ+TYLTTVd6Ux3Uy+pDYtgkmjmuunm/WUJupFo6o2g
gnojcJLOyBigRPZxUux4QJoJq026Oub/n8sJKTAlg8/JwSXMpdzsH01aRDHBoyxDw9F6jR5U8zzG
krlpC35Ui1elZIyWkED7LbXzyTLmbxD6OfSmYsRfm9gObsSAR4+2Haeif/vmRP7nE+ZkWBF7HO2S
plsW8PlFsTnGSrgVR47omxyvk4H/BKLWw5P6LagBvR1V/Q7143oT6P9zf+JqfyHyEkQJqcXRRGiX
lHmpZTp0zXEHQYliKE5w5wm5D5PO982Rm/jGyITA0SHOcnwi6+ej5f/lz7m0uQb9jWjiOHEiWf0a
7Qr9Fh5Mjxtni/MPhEYhLi/U9vLeWMGrnrCg9FD5YTgfVsXOJrx7/iyGGZDpRcJmHzXOiwjuXzZK
bw5G6F7myDvGq48mPTY6KDbgpnHkdSrRkYfB3hvDSxepXoG7xVlhsdRJrENIxIbjtbe3RroKz3m5
x9ImfZOvFtc4JAsaZnwMH8NBFFp74YLxAKlkoII2S+O6GpdKy/4+cMAVcHScy7oHkTiclL1K5OrY
YEZGWkTdbj7w1GGcEG6nPoEO/2yoP7rCoxeEFjKOx/8t45JvpsCp47FOItuaxs3KED3pliaTzt3F
TKU2AKaT8N4MOyH1Ywe+cl1Fsqer6wWWe2lxA/nRteOTqT3ZGBd7QB+dHesSr9SopzXQZBIWnP+M
sUlvLZoGVHCeDJ/745HY9AvVMIZzH3lAvnR7STTysouMScfwq4FTV23PiLn2s9pNAZ2JNQk8US7m
AqUqOmfk6U4lbzZhTvafAmesQuE6ASAfv/nGGeB63fI6+XFprpYOyvpYwBADscGMSDRdPQyflRQt
Kbs4r9NvfKR9CymYg0wSTojQMPCGKVOMAYYZB3PAMU0lOYVwcV+cqWJ2WTcncVgDsHP7vU3/rW8Q
Zh4cueGyWz6Gi1AEcMi16kDDeH6uI/wHUQLVfjtSCri+gkACkUpir7E5+wVGztNLIcLhZrJTlfnZ
NR4rTDt9JGRh4/zJ5qVxo03MxMpZ0tq3jQx34ayKUU3y0q75PP82WPesW0cmZumAx7XkYG7RBS7O
DLfFz9yppeb3aS83OUounQ04jg4n04S6rcP1wRhMaCrwF6sjESkL2A6VH22C9Do7jK/xoabbnLGK
aF5lpHmup/GBjGmzO9n1/ZeifzvMAH602saX3NuQHlmdjqYE/csGB1Zy8akmY1oO1+T4/UnzKnCV
kkQOv458HfX0RazE7HHmjdADcr19ce3iA0GD/wJ/KN05fXRMmnd9n+dpBev6jBrlvFF0Msd5tsTg
k067voeTU26Xsc7Dr/p7GwPYLoVQviyitWwb10VoISojx0L5I313SnIH+hgNjzyIuUs/m8jN9FVz
LFoMwlb2GSXNdjWWfH3nl0I3auM/6rS3CP61uAknwG6R8xU1uiHCPPriWuswutCgwuqZe2MQn06z
BFtJd9sliFTBwG42AlLCCReqQWSEtjKn6TQjkwsxdHmT4oUVhuajUz3bltRM1aA4bzkU/yTcuA1e
29MjP74CtcdFDo54/1zP6TbrWuquTqJ7+G7tNd4ON++xN6N8Ky7Te/OThCPnoMbH60QuqFhAq21/
xujqn6Rpv5MT+xnnAMxLPofioWUVhmLkq9/MLHcEL2JJ+8CzMQXxxEFpufu0I2Bma4UJmV6AShCV
eIst44ylasRBKgGSTM1jR3Y8oJmchIUF7xp+l96Atd+xGjBdrV+x/NHKhK0+c4GHkqHPVIOLoVq8
N5NyFHPDkUj2FRAqR24+wqjlp+SYK5UhmtWkpXTnOmFOz5NhgwHvHi5so02Ne7C/6Keg++06N6+l
GbuEokLoLI540tIw6lqrH7aeClIglVW/8wm3oJ+ygOFUgkgJYU7c9q6ry9TUMwHKzK/Z/t4z4h/+
HQsT2vhIzi5BvssN1eVBiXzAYAqLZy9J5gwO4TaQ5e4IfJZtjbyEtJgHWvI0N02YIpg8Iatf/12y
+/8CZg11k6rLLXKEnBYWCHq34SMNdw80+6LYV3wISg3KVzHLcB+zniBntSEMSBBkUsSVOUxCWiEU
4A9/SmjYdn9H9IJdncGbAp3dUZeJKZQ7HJYkIV0BTkmwzx1X5S7gWnNhEcAz+VrZfOvC6KDQUBfx
KtZ40YFN3L7D+3X69EKddh/757gV38UI7nGot4kt0izl8zOCpTuKrZv1riyKeJH46mpZ3X7iyAu6
5kPYgsfm+46M8KX8IpAgulHTn+yRRP/5XzEuM92zRbp5d9EZqlG/8u4gr+J21kXdLfsftSWJPDr5
rPGeviwsmIuOnWjZPdfOV0Ov8iH05Sy3hScHlpNZW7pVrPX6001SnLi9saZYTrng2VBwQI99/xj6
pj31KlBNCePSfh20b9qJSuBTMQueUcMvIzkXwWFicSmv46m6ANWIHNgdKh/PlwJqIrY/uslN14Cx
bqeHJZP9EINankRLnmH+k8/mSBjUprMyWLzp/uu87Uq0cI95ncbJn3+pPhYpCIuA0dZIWpJ56Xcm
rvqoSuaUMT2Kq+lXYPeSzmHBpqUhM/fqEl/tLRt5vo4255n+YbmsPPLhA0Jt409ugdNU779VnJM6
08w9oC0xxHvy7udkOJvmYqU12dSHC3YG7t6071VFKPtVgB43870qQZFc2WnZ//QjEuP/3KVvEH6k
wxMJm4/6Hvu6fDG/Z8xrTm+CA8dsKmYk/alAtEiwlosAShTA9IG2/cB8CT/bgVrZAxWtTvphBbXV
mRy9Ai9eZwpJE3bQZ4+r9WL5CLIKMN/A8jpReyDoXDsScaYKW3P2nXW29cOZYjRnb6+zWd04jg60
OrEbVA/QcI5YCrEJqVsk1fKUp4ep7s4V23MeOX4DYgDnCh/Wmg0LJQ2EBqfRtf8dZxOB+PNn7usR
1rscKG7ieTqQyBzJ08rEdOAczYPsL12MSBSZjMN7gzHOBRGdwhrAUi+eyircHrNenHwN6DGDK6wE
WSu7RLcG3tQhZY+rohO0aKsgyToMiMpKWBpKAJ9pHqnkyNqXen/H+MvG7MkxbXNuAUKBKPb/XN74
mxo2KydbmHQT8CiZ0gIx1nQsE9aFfKHfnrtJz/VgX/CQ5WcbOQo5jwQw14Pkp2RuF5PNPIPU6Uww
rphZzzL1bDifsxmg3rOLR24JR2HUs3GmMiU4fXl9PqInpjtg6RWD9zhn/XqJC8zLoTvaIXfgl69f
Jgb5Ip0dmQu48i5PDJSziigAdSoxSls5Yj9+C2BbNQ65StMBHrfTuuqy9GrdjpePbhie0cOofA9p
jvLp2NDKhvFEJp1iu5funR3rhjeFF5bMzb9ilCBEV0hBy6+qmX/ewtmdlqUF6tgasa0lO3Swie+W
fo83gavgvLmi59nlYV22zeO/gMkBMf/VGoMh54YKred2NPrNJ2Koy8qiqGRYufVTDWeoCfBO7ikg
wuojN5fRJ20CV0tTJzYKFwaSllvhHwLPxZAO/K9hh5T7V4VOzj6OrsUwxt+krniiH4Q92VStgtV+
0b9Lv8Gbu2p+tfOmt2ZSimOlc8tn7+fTEUVSNzE2l0Udw7TkFWUm0E2prqq62zpkiBBAeUo/YZpC
rL0amDlEHrylwVUwxDgnNVJhDSaAgm4ajipoi01XLDXOi+AJSdGOlZakia8OK6OScbyHevOc11mW
6rlrfZSPWKWlE9RG4B0W085rq/GE3K4ZRP3uuuX2cIRN9J9VtYb4bqII9A+jI2JDwcja5XtFsEhJ
pHCra4gZ7E09pgy6k0E7B+X8mjwX4qdjj64hFyXgEpQ5htZs7xarHq0AhTaFCeW978o0RphZ+OOa
VmmVLKsQFY5shP6pYp+Oho7wqOO4XYhTnsnsIn0Ksl3mqGBzV737hwrVyCDkRBbe0qCFADyNh6JB
yHfq59cuyhSPwIdtLIpZi9upYHkkp9KPkCQ3upuBlRUZDZo/vP/NOUZOfqgi3kFvKrykW0TFe1+6
hNGxQJ6FA4KXtAPX49AzCaHd7QuJLeWm1q8CurEsvkHmGwLFyZHoUxzHluS2ISWvC6NHLWhZ73kr
aDFz0Nr5sy/Xdszf5btBG7O4StooCdwTfKZcpNBD1lM6P4sxxdr1HF2AjyxmnMYP75ZWdBuTvUY8
WCuWz9t2dkByG7jU/TPg9vLVits6s5IRrlgmXDpprPISSHkkZBn1yN+jWnIU3SyCcU2af3EcRZlQ
0ftGzqrwlvANwvhxymzNiohmoAyTEdawcQ6HtaehbouQq7LsmgtSSF1uzYghgnCRdYopR7+uEFgR
AbuKb+H5KK4nA1cefAMSovB4E7sXJzjqLZfcJD/ZTQRfR61oAaf6JruIjHOQCis3cnMe5hj4MMV5
G9AOE6ICn+AbLHhXYkin7O3od+ViYBBI7jF82c0VXMBKEGzz6iNVaLUxye9H/8UvAbtxBzk9qGpX
re1J5K6+o7QIY7fSi0mxZ0tpjp+TaR83EpCSJbOrFDzyFhQa/Dw0dsO82Nu6do3WFKwGL3fCP/Hp
eH2qOsUhmLZmZtigkOtqbGhdIlNmoLvaNDlgLBrR2CzbNepqaXM4H0fQoAawcZ5Zn7BGNxvaOMIr
TUzUaENNCSb1xgG9oTRpR3xvRGbcKe7H/nXvgYsbfd7H3ebAVc3OfQMYEmwR/SsHMbUklCn8O07h
WuHfzVs1Flkpln8DoCOU794LlLLJFEY3MH5zXlpgkmtsrt2QX8ou8tQ/Qw3Mpdh2YFua+7hhIuLr
aoPyWmDsl4jkiWPD6WqmxZbndnHf2P7xTVqZurs57QF86XxcDLEitidZvfBNtLQGwlzbVkVvWqIr
OqFrCGBPQZGsYzsWDC16/jxUTSt82pTXgijRsGsWddL3EBbwueM2Bp+TmWRWZZr9Zj9EcnBbZ76N
JYeoI3uOMkDNAAPXvRue+dRLeZnki4VGxqcWEG2VI/ebzBHQWp+CEMhBj/PoOzZY7nqyGxY/hRRL
ramXH7zSLFsQqHFdnZMjfABpCrjnrCdxNDvHqFBCGJOkx8FoipLsreKMTX/XhQN0J3x8j+ymcUJd
tME2X1T/RyjneocWIjs32v9EymAhSyfLZXmfs6b0Z2fsEbTOKQi3+Y8ZPfMWZSLntc5cGG2DIOpK
CPkv3D2w10XSiYW1zDgAZKv6eGM53DNSDy/f+/ffikYLmbFnkXqb2SIh/8+d5pPCqXAupdhGJWX2
aLiwGzljInr1hg5etaoodxiLCY69kkpAHoQAExv4r3TsrjdusqDhb4gh2PG9zD75lVTrpbZAuQ8p
fUXN8Bc37f1hna6QP8gLt32+sWJ4rFUd84pu9ClxbdR2K9VNdsS87ZYRTrGo+kSyEsAWvCft7o8x
CjWTCypZMkdrT8Gvck/Ybm1G9CPNuAtf0+3K9woXIrS5gE4ZINh+G+Phl276jvELowsnhWIn1fxa
qBJ+IsxbjdQhxyZfR/Jad/myz6J1//JVkvsTO3oAPWyl66FAnMHwywi7y/OUDHa5ZDdlChLeDqES
mRSjFlgtBuAytgJ9k6KeWSxnI70ZNj8KWI9TfYvEGL2dYIU5MOYsynB6oiTzhh4UrP46ziYKDy/6
eHxWwsN6+fbaNdorTWRp3Ma1tlANGpDck3hCCkSNPoKf5AUC/oS+fsKJcA/CNXa7HaAn71/3AWxF
Ua8t+VsPGkZnJNPIpf7+4Uia6hitOuHASUbc7uTzmCTBTI6/Tkkb65LttY3+KbBpsIChXwBdslhL
ezaLxMtVtlKp1OXpSI7m4mG5mDL/uOE9OxwVMYEfhLElDVTlbqxFhqMmA8vPKKUIqNlNVRuwfTuF
cqTIfZVw6FpLQ5vDThvA04GAzpmW/AASU83dQzwPkPfK7sx0cwM6iWXXmdyLlMlXk1QoJctC/gX8
A5keBPxQ+UaWkrhmWAeBYqXNhuycRub0I1OPYb7yrHEe+009bXEkIzzNxWsiFEafCED4pwRrq/va
fbWoq0OTLUkDN9iR27P6kZTnfmewCDmdlOEUTD7p4O3p4wJpIjEGOkbAdszbFJRxSauCbGrhHHDK
XAsxJ/e6NeoR38PtQLKSFQcbtv8+LqHsKVU0yH2fJI8Pks7K5r/vkYOe/MhAFTNzp87dwl1Ifw3Y
+LHfuEKkuwtJ7XX2qtktjFIH9QnrY104y1TUHKYWKmKZNKDWxjUlDPHOQK4fqnYE2WSnfvaUdv2c
BIgA0j3ppJ2R3CsyWH7nh1qDFN3g60lbxOD6NoAgivRmAZabGrloI5Yw/BqUGKhtjsF90nDQ/Rle
9tSVaz25c6rdHWPxINEjm6xMLQ2WnAIxGFi0vok276bRprxNan+KwnSqgwckbs4X8TXlch/6126Q
RFP9WNa/5ErQ6MnULBb5/zpXEfQorHRM9nqMKmL8sv8pvB86kiU4WG1ypRyy3UCa9VoK8+92AvCU
LVI3WOEa1CdDhMVtT0VJiywx9NPh3e2S1GpaKE7ehIGtdJIdcpOZEJhWRXzWSPWhbIGYgbVeF8Ol
gSAjVTLMmWHRJWLV7i8J5g9U/i7sGtcy/zi2k0MiwS0etutcnHdWrU5DVp+QP31uFl3t1S4Wdksc
J2p7jvgGu+KCOUj5s6SEEp4NtZMbm5NesGwyHqGCov78rOgpRXo8IJsIhDY1KHbmlV6QhcSRBpd0
IRo/wHpEZ6bn1IhajdBRxSSW2JLh7ygw+iCTYNtul9U2A53Tgbtg94aJBQCy/KHKop+Wrpi8MJQv
HMKZGFYh0N+JqrHcqNC2eBDhKPzzjQUEOyzOyHislSLV9EAoZKNfkmO0bRlTwKsMmRfOxRjZJWSf
6dBF3DR1++hEdd6QIJfW5QDn6vAf8fgsi9MoymgqjrqXAGkmHJ241fpxeX5N9knWWxzTKRpO6xof
rknvIeztGrCYASUGCsMdNqQP1JTERYpbTgkuH4FHObRvdJbP4mekbqRomc4AAqI8Qay+5teH/tsA
sfaYW+ijaRYxOLpJ+LGdjtaKhlwnG7gD1DhNVQ/JcGKiHpJCaj434KVFvg1p1++vhNS2nQljwlv7
JcQhZIXz20yGn3A7cj87XZpnoWD4y/5o4UVFvH+VSxp4wvVe0PSqsARCfFPvYxi0laEERK3kUe2s
cK5147/GpSG51AvCm59iCJ3OetWu1yfc5sewnX38xuw4su/KvRUDi2hT+4QAUVWbIShZdyU37I4U
KhXMFOm2/vakUjmTGKZWTjkRL2gLiCL4dJBotWFdSJ3jdhTd7taOuIuqsv4HeSHKaBEhnq1b0ONZ
2X90u30/Yu7fXeB0BGLKoUzQIfSlVtYP0tdKZyh93j+Ty5u6G4G4JOct8RHq58WwmAEzMG6mq22d
guq7T6LNN4wIJVf7lQRIIHPGvfwP+iP7y4kOnMIqZLBfsrrwgVWkn0VVvNgY4U7N8mWtW1SiqQgC
oXAtd4hR6odXFxzD1b0QxBumoeSI00dYRPWdw7AmKDTG1JBVfWgXvtTiEDj8pDGkrxz4X5h8csMP
OHU1zm8ICgJS8CYj3v+YEhRUycSmRCJAsC6G55E3dv6EMC7wfdOaj0r44KjUGd9pCDHvoB2UFeJ/
1Dwunvw74IDZd7i3ly+Qe91kCJ/RK4vmQ/wxfbKcnBqKP/V3wSbn7yIZ1YCBSx4emB+EDKjK9CXY
ten2AN2g/bDAp3z9EdzACxnwFnAdmsbi+Z2WDCQyaTnaR3Btbxxz8DERh3X6NLpI97Nk1WfGjh+J
DQRDRbXNlG+dsOdOED7YMQG0ITr5eW3g/0mC1TVGfcA1nFHxUjFM2ea4fhM05AJySYUa+Twz7W0H
oZdcFeQiVvJ4XPGotne9nuzfcz1ug5Pht2uzDwYO2ak0QTtyaksHrzwKQR8it3DsBLM1Uf8+7Jrm
rY0mh5Yki5fS/SJKHyd6ZGCJvOHBtJEV7Llj82/9IAmNMb8rsk5Z+PSxAS4j/6x4udS/H3PGXBSn
CfkgIKqS/kyt/hMbCb2xXJhq0twwZjemKXdpXbKUKN9IOisJ1CvKmb1bT6bW4vFGJHVr7ZKDpSr4
egWtuRGUV0u1wZEg4kQpp38csNlhLhxNJSq2F5tfPgiWW2HwhVdGTWHaIDAFNYtS3CTVmuqDY7Bm
BiemVN5UpQgRO4W+m/s/AyW9DY2M5RjeeAlkLXMdcFSUB6B3sEoEZ+t9ZZfzpKpYbvUKer7m/FHy
R+X/jRsnMt89ovwRBs6TDaj2abji4CZSTGDF/O6YYncys58S3MKp8fRDiRIidUXy4gWVOEOU73h7
EMhyuWjcxzJSusGbh3fFXxbbLUcv2cKtSbXu+B/K75/nUhu79vXJCONDVzG2vn301x4NaLZKkS3H
ziP7HXljixJ7wxVAiwpPpg9QkET1OCHW5KQxkW2ogJcSZ4EhLGwxEAqaOOEZB/kn3VvnBEyGKVMP
S5NDhMd2yZcSHPxKzKzo6MYh+aeRCj0+oeLNs+QSi82EdIFJaSf+dBwZUBgz4p5MQbt4VXsIyo1n
EvT7KWEG1ID97sUvUosahLItiL1uu7hT0BQwNJT3jxLufTlHn5OZaAx/2ROYrwmZCrLl8ssRTJB5
7XD0l5T56NRVvs+dcYXgZDKQ2UJvkweTuS5J4p9wMDJ2EvuazBIg68G+8s+XqG/ZoE/wU9psqflo
K7f5GSOzKzSFZwsfdthytT5rbOL5Ln2r8sW5aaKozPcl84eTkG+oILaQ2Q/pIuGc2DiaoiKWrIe8
EDXjSX4UebabgKCmy6lrZbDXO4jeaPMjYkLLJZximBa8KKDRI/K6dpljpJtPitwhpStosQFuorTT
r7cY2IGGwOQglrt/AJQR+fCGLr/Vpc6mkVQPsl9KjddkCnIgPxo+ki9vVpuA51v9z7h7EgxPEm67
2QPcyAWyFm4NKS9QOCbs+4eaan8ZuewhH73NYJc/NrKqKJEV0OSSCibg8h/AV/pga9Me7Aw+Yl4T
nqZ6zgYoGNBPMjcR4vu2lxIrpQAjYtwPCYe7nqpbs/vFoo7sA9C9AJ+XsUmRD8Uao1tD6w9EnY6V
c+JknYoerEbAuR575tSOaeGfOczfoA/9c1+FKKrW2mg+VAGej4Lsf+9ldlH28Fec/kJdQRFsH9SO
A/FoZjAuzv7100/Ym+9lpehvGtdoyI7DgxioNnCLppYPDZQ1VO3bCP7F26T8guAiuckVFhpw7ZMM
K7nny+Y2M7GFgeAtIHgXbBxw0PsCk7Mr2Y8sm9g1gzcwk5rThOdY4L47ccG9XRRdrlI014xOwwS2
VY+o8wB9FfjiC4a7WCWaq+J6G3Gy8C42uCRYkFSC1RDAJjkNlyG5nyfFOUavrUTDIsl3o2cbSTIs
JzXjAzID9uSia/HLaogUAo2IZ+DcO234faFn1heRAUNiPsMPRuh1nFKUdCZYYMSXvMwq2mYh2ZkC
f3enBm69+z++HAAwdzscoeK4g3/GM0EeTaOYRTZDvolKt/IXNh8vIH3TGBfi4S5Cb8oUVFg00gYa
Pcp0oQfe+8LFa37vD3oM5rtIHd0HSGWSJ+AtxyWO442sZapDswGfk2W/f2NENgzp6yXVqyopk7ij
eD2J74GAAOitT9AnQetTHB2cvR7q8tEdxaLFhhR7Pnr0wyFndEDrgYgnHijTkmybgRnSCG1zn+20
uZ1n0nP1i5u3pRHDQXHckHvCbyAvfoiJW9d7YKW+K0gmd/teba8HnwWo4OidPzNopJ3Urvf7+WmU
9E+vnuGGWtMlVFC9ZgE2bRJZy94olVoIEecDvMF7LgtlTl1V+5b9Kccos4u3UULB4Z/5OLBiaAUu
Ecv7Ri0IqCTqXjk3V0TTuJFNuoYAaX3Jhmbd8OQlozOTt7IDRI2JaN+0Ege43jWe4KOMZJbWVmnR
pl00qNlBBaiBFh/goO3P7p/70ui48zmjeEEo76bvQ+vNVM5J1TzLK/oCyzBU9csQMhYjHUvF13PG
aLQDjZM5BQ3258BDKihvHaJlSsIKgJfkfHOV5s/Rnix81fkbJWa3y11PAwQhHOQm3u7AzEG4b7/U
yhuimCd9mWOUCS+G01SvCyT8oz9LmPgQi+z//WgSXHIaaL5U5p/98rS5zBjq67WAQyNcT3YHnpDE
b6WSetQFb30c4OHtorNHFBtIFCS8sH1pK9QLc3LAzdcbPJcnKrdnihN00g1ghex0zvckQxxICV1n
m3Qa7mpsChOFc2Z7j81iqGTbwlTIhXnaeC92udBgI/jJhN8mQYSikwYxrurUMT793peCsKoKfqAu
njjzK4WsWWxkN2aX6mJz/EUHxusKgZ8W6vuGWo+UC+pjigtcaZAVbaNJ19PE93ZpNnHLF27yKTGr
xpcH/SP6WRtHPqjZWUfNtCdDLXngqZr4GFWeC2/baKjM8z4q04R/zMxow6//Z2nWtB2ZK0gGK3HD
HWembfkqgBW6IMHl7FFo6rRNq4ANVGvZJCgHIrrQqG+ABeeuMOVhLVt0DI5c+PjQ+/teincm4qlE
dpIEypuApc/4tG2lS5bjnwivz5pipWGyL/PxA15xY2/QtVaBl/ioTXqZBSSCCBgToITUMqbuUzfB
M6wdcqKqJhGda0u/UMZIgpmDiMiWzC8zqDnOi80J8oUjQAA9tK0FH19D3mqaK4EIDVUaw8WhtCQW
YvYExT7bMbhjnzQm1uuFs/Pv2JbFEuUGf4fDfK8kOenhwHtRiJwJkvmW2BCwt2EM98ZvnYAmbzLF
Th/+tAOMGrOB2mh8SdY9qL7c2kDyGpWtYsWMlc8On9DtgLf7xNXX5yb7VN6DZtCj11U4gr3DQOA+
doK9KMsBwWipqVFLP4M1JlMGKA0x3lS9tK8lFiwGO7u52JoBpD2HhD7YvvyII5nuRWNcHBB5qvpM
xRLbeBjj8Fnu4hSHjorhCnxbliVh64Isqc4HmHt0LQv0o+ZhKA9peP4vynyr6kjUwoTJKLX7zmCZ
aPJLQ4VvVmnw3QGKy+YpizkM2Rdh9tbA8CWyTYz4ytCaChDEZGhm7kfg3WOJ0mwlS3tjqD6qpJII
+4K425QKBH3FIkvuIWqvs0J9AZnxtR8goqDRh3Da0DrXs8FDU5ybjOvtis6i77+Y3wwEU4CNnpH5
9Lg5ttvxNef/j7wKk8lzavpTflWqpXQWTVon8X9g+bD01BuyqbTEByDEY9Dqcznqpkp819BwJHqn
jdhz4ET7QzjB52aOgtnxaDHDsttwXvoxlFTuHjn1i+cySaiWF3WsEO+9NUmnqnjdRt/ivuHrm/PG
OaRDgy//UVDUkIJVXMk4rUZWsDLFuWnPkhPoAcjAehuRvqn4830j1FK67WqxtVqbZTMvgGUHEu/c
D0Ah/DDiD2xV8Ribx7xiGS7FyHKFytML3DQUgxMhIY3L1TVPLtkucIuRaDg4aA5RRRHwrUSI/v5P
tbDkSHksA+hpw9YRV8mq3UhODAKqiY7my3lVQoOQcmoezW1NgqLk6dcyycFbl/pxfz0otnYKDqvk
NbjE5cNArRRC9oHn6idpyBpUBv6VOhI9dgIakw1HSxr5kfV8/sRIkQgxjyD65CJKJnOLbY7eiR/c
FkRHCNb+n8W+nhsAiNsgJSsTtT4GZxOWPmnkqLFv8eiAkVO4rsQ/OqG7Miwp8Aoq/E+vNpWpGYGi
ugx8tmIB06Dy0lbGzi8BCe5ZRZ+94LmEHoPknMH4yxjj1jlZ6kC3iAOfPwaRAmj0GWvFfW0B1dNf
fwNgF7q9YSVSzD92JjrzRC25a87lAFeVhPY5v/wTYf7g+L59Fg1gLwnOB3af/+ZCn6bfqZMLOJKT
nrF7MOpeb1rEJ3nJr8EgeBQv/fe9GpRJbCL/GQTleEpJjVuuH1S0p4YUCLr27q4UrmhdGeGtU2zd
FcUb2z6nVpwe9qS8O9pNp67R5Tdt8hR+/QOml0tZ0P5GjNOCH/iRyU+FG/IiJYCRWOydC+g0NcsI
3lJecrElkbHQ0zsyK7qciyb36zQnIAd/VCnlEC45xoZDsGoWE+oo+G/LCeF3gp0eyfBPjXjps2WW
o8EZX4ulDD3eCke4vNnK5h/JIVlxLmfZrDKSixLtEvggaPjUWt9EhoQvoGAd5G7d80gDNz8BATqm
6bS2bZnXQXRVQG2UZs+FsTI2EufISR7KahQxn+8/6SnpGYLh7D5KmcgZZ26l4GKcDzQkrse7HIpL
uGrpwMWOh2a1zS4UfGdCqIjOeVmM8KpfhcUd47DDtyuuJ1iuglyhu+oYrRgqrYMNuyQK3CuQaDoe
ceAPCGWLHuddzcHJImeqsPSJmQMdZID7/Ld1IK088JS+DygM2OQH4hWZOjfwTmPvICqGh1LbSzeK
4ZbkYf368JjnLst0vSU+KD6n5ffQGQk+WVKt1S2+QvzxjPbEk9JeSOaH4cvnDPAzTL7FitNdForF
bnGME7qONdVCG0Kx76lY/tHNRWN3bfIpVOegCAGqb5CNHSPUaUCK+0BekJgfhODvhtGz9vR9eFHm
vP39HO8SUJUkkb627HR3BDvZIDTnDWafdO9fEAeyEWzU88fNbH8Sb9BUOK6WiugwWLuOk+OWdU5l
Pw8qo2KhxF5jeAtnD9V4ajhK+F2vU6MK1I1vxMd/ELBed9pBa58HbcGphGZYFNOaeQre4j1bYozb
wHPNTINklb7BgT2frDYoTvCtBCOV48Kf1qdwhW7tnagHxsdW8v6MUbW/kXKOT0PA4d/jpXWz2ExK
CdCfGkk8lan2tq/awApxOi8muGELYE5SftuI2OUOzz+JVF2t/wDXpNNChauwraPKrI/TttJJHEkq
3hATIM6lkHEdLSk9A0XBxMdx/bKlDjz6w336S6ih+7103sBbDjuBjfzi80Df1xoWH5Y1kKR60dQf
EVqHzkF06pc9IrREd+Krl+9UUPBhLfG7qf1eB4haQPW/BdfS6wh7chwhvdcNh/A66vE1D0pIeWup
LCYAsznp3QoLVINCFcSjXBOtXmhbOL6ImaMg26CHxWZF99InpTFlQHCsz4JtA31M3uYiDzolPG6U
C/1wpvAx8HkuCNuuEeLn6bI1+xfSpsBeBri8A8Jt+Igq8QWkPLmOUE+btsRHx7/Qp8S+g5WCmD89
SyEspJv5W/IHjdkzfDIzNlTH8c83eeZDSgyg9As3K0sML41S/NivhcFy5x8cNazRJIXffALU/AlN
E/uo3tm4aXdDek5plnhM4RUI/GoLo/53gJOThHkELhTVn+QXmuwpPqRj46DvMHFBGIQoWes8WDnR
x5yxDDfI/6au/RHGYDm+NbuVQFzWFCzkbwxsKjSbOsqDuHktmRDI8bicGeBJrxkTCFeCxwQReNlR
QtkfWHPIFw8DP5hFhP/onQD8L8YvfMQtJQlklvqxEBlt4V6H9S0lRnVxkwqEnlfPo6WJ1ZiPn1NE
FbsSgdgWoYTU6Hg2yHVlg+MU5mdQfyMExawofOqZA/CoVQven0HZcIAiO+ICMbWZD1RWzBuYu0yG
YURbJGsmZPKHOW/wf2a3NQz2EFSnEvez3M/QWJekJAMPwNT+te+aPHAH/SCWyZtASyg0OIfSmQEG
9emFZmGq3NaCDFr7YUkpkSzDanvvSqOTniGNE/OA/0+3aMPMe/Wl+OkwqhXVG0e3zk174f+jfVpC
ZqYQB8kVwunOZJS+5pWOM3nfPuJkEOUCzZd+Vl6ZeIxVibv0qypXHn1vZq4PfKpIu4IYD3zUZVDG
CLkboyglt7ujWuzuhbHVa8OiKPjLOqfTMtY1GAInCAuZDzkdzywUia99HKzPRZYW+4bFITsNvHJZ
8JXtmefwau8HnJux5DEPW3vh/W484+DgHLbmGAYCGaG62MGjgSGSHXrY/cj+Bzf59nRe2mWGpKJM
zRlHV7XUoluGscI7t980ZQJsC2AHrmaD32bgkbVSY79bI9QBtbS9AmuDw8R2g9uvojwQw/DXoyZq
wP+j9tAb2tVn31STEO6HDByYGInFYL/GdqeZr6vAovWBio5jMoeksfw9TNP+JbN1SaFv1kY6w90w
Ocf9i2SVLFP+TgG1JwWDKpTWRoiJviqqYIrOZTKWVON5t72BAkA8B3jKGOuouJzZpQS//QeS6kh/
lHxAC/aZYGbnsW9yHYhMEBoCPYFy7bFx1Y6eJoHIXA/NXiByzkK0xk6U38RyPK6rqfkk6I5wSV8D
q6fEpovLpUD9r+r46gcdBpxAP+r1msCd3pJ5cSYZFkzR74OIVxDvHas4pW607hGT3NlnnfemzMH+
v3Gs69hR2+RhMNAsQ7MkW0N+QFoC/61+qmv6rcLwJLkOR4Y5qj+JfpAFF6f6iwgu04zIP7hZUWM1
qgpVA5dnyZpJKs3DYDB3yL1r0OpZVqOyxajlgfU0YOnO2wJAyoIp8MWfR6AA1z45l+hcXEc+QtL9
5cIlCkYRzsSjgTqXFXn/Pb8eNV+RLJLDnt9a4UmWpFwTruNrHuWqvTy/bQHCbjugUukniRW5Mz99
otmTUT/ISDx7mHRfZNIJSIGokpN3fsRhtzJ4Dr/tHhC+X73+b4TVPhkes7hbYXwmrXXwEGeXuokY
/v3UHYjE6iVOG3AVrJohnIsqLph9aCqFESZuREjfND2t7EcIpsU6tvL6w5h0dLbERmAGvyf7E3H6
tbi+pouaMbCbWPZ1n8XaPJ/tPJMf+BqVypJPUvy0wnk3WxPK6gmBdfBaLm1uHYtwMMuuOhY1dRYv
QZFqtm0gx88udOxAWyU7cXXBeOoln+LEpAqoxrmJxh6xPzQHtdzvv/FdX5kpHBoKsPLqC1NSJr9I
jAEWS6r196VlmDMCGX+Or7MaNCd3sb7U36l0QbH1x5+ue/f9SwZYC3AY5u+ZMCvfrPbw/D9aAFml
cYe8rGatDrvA7bcKBB1mJgjJGjquxMidY/Hsw7pLDrynlniKMNZqreqFGglDlAzbH9jT4Kae3K01
H5U1P7HYRNWbnqhqhzUdeIGnRcx4+7op89v1o42nbn4nfLXfUthQCzw6SbOU3yYXtxL485Cr9zQN
WKFhjqcoDEH0Wp7WzMmKaAva3mtxXPlsSFSsAUjPl1lbwybpBO3qoUYlrjUHebUeyQDeBfkvkqjj
UbioYwZYunWbdm/xY61Vw+sa2MSFWK8U528g/gmFeg2pa1fiSuPKZB22SdWEhcteLdB2XVSTGmzm
AoSuREStsblF88cX1d6JjeMNEZdt8D41QrfrvWLF8rKuazcbWT76di4+SBl8+es0m7AEawntKUZ7
3VW36/1ePMptPWQPw/QP7Qq7TklQtWkv32Zfu6nMUB4j4FeSVhjRXFXlVZFZPbSb9UNSv9sFqi7X
gt0/3NmFpfxhZKmVTZab1dklEaiJiEFXvPaJaPK1mm2jD+9YF+YlHwDAYHNT5lNdKthNKyNrpw8D
cGFX/679yhzX/PTMkkO5aroObHtE6leooNr8MUNduKjZgOSZWnviDE4fqPjIn8fmJ7Kt1gxnAcrZ
MDVz7qL97g7XaRhPmVX4Xb+ZmjYGjK5l5mCeLGg44GzAVTtMgyUxVPJsLXh81tqnGlYzBXlKL0bn
VgQxE/vv1/5nsl+SrS90w+iAYX1C+vwkELyomnMXJJahEZ3vC7GdCWK/o8CmqCwHDBYBeHYQDSM0
47B3F+XlbwHUNmGiy2WkpDMZu79tzcELD8StXlZ2qFU3nEqw4+YSjXbVHrDn5CEHlEo0Ep45ZUit
rtt76DolOwBnb8ZzjZi6CHuuYoV7AVh8LN7mCdHzFm52ek43jDHb6PDZzdFC6h7080GP2f0CkAEN
L8oDc8onbiEnnin5AvMEpUB480O/usziT97BXO0TNrX3x1pOvVNnJ+W2aagQmsfWnG3xe1cNU3I5
EYoVOOMl9xKijO1JhmgxZo/NCFRJcy4522PXK3k96HIA3V7vodB1P9myGIpizQV7yjEPSaNg8w1F
U+10uHH8qijlf2VM4McDzjD/e2q8X0NzrYnnB7ROPjul0jnLL42bInQgBbbWmM4iyNcU8qVFCIw4
T9lXKcMKJ/DfA9qlG8j89QP51Y94Mb9hs5sO7Y7gbip+0cc0a+BiJjPZZVcExajVb7aEvuSMRmOC
Cib7TA1lRQv2ZqKOD7zf7v2QwvsPSahlT+8fRMwRXbAySFKfJVc0aO3cFoQobvYAUXsdTEzfPh76
SoxQXII06aRP6YOwQ1Ey0uJtNXqvABiU1bMFhnWrJApvziRPLvQbGq/PfkaN+ZfbX+/tIlc4VZcy
WHqay/2vcI0ZBC8Cv3Aa2ygQ7Mzc1iheDlFWH4jzUzuZ6J2dJWCYUqi1Xt+DZ5gUoqG/nhMWFyAz
PzVmtrVWHb0/LvJbocljM3Bv6VAA2Cd6VQQ/QBx57ndy2b4QIkVPI6Guq0O0Fqx7EPxc9zrqIVXp
23/hhpKJAkqGp2lQ2Mfe1eTUCiS5sHhi4VAINAsfRk2CUPBRC1OO7VULCeIvo/vPq1YWjI3uoPio
LZ3vk2hPgVgsqEg29yeA6UuGewNdd/Fp9UTIN8Wk99bfaynJslW9W6Zoe8Fz5yg5Tp6XZbVWVTSc
N4rmDp5hztrmzr9KV+hEXbDnjmVB0hI82A64alx7ZBWfKDI48i1fHU5QtNro1eLx1pDGmI1Nz5G9
vUwj2sWUU2x5XnB4lw75PL3dwi9jLEeiOwGPsoF+pnEwsH7v5kI3fvsYMQBNEqWD6KQ8Niy4HsUz
X2GSzifB7LuCIbof67cM+23cnMKdBSfpdB0bwXYOLRl47ayKUb6aLEF4vTEs7Ker2hqT7a1NP7mK
nHtg2GOsShLr96w1tCPb4gQtO9adq+RVgOY/bi0Af7y7orsidyO8Wd/i195he8rAv7Ur5nKOeW9y
saK7r1e33BrUc7loM8DArCbYF3dAC7UBgvy39P54MnAnDKJf3mjjiBn3DL8pBhrgNzeE9B7nnxUZ
LolnxkXfXdwjRMWpffgYdzzfzfOAdCOffop3R4FYH7zyTAww3HoKbju4Whxqy0G9gXMgOICAAabm
t2zMfjMRNHcK8tSRnh/gUYe+heIzmtZX32JXYMIY8EVSKPYSP86Zd8ND9YdRID2MU4w6poC6YI8T
ZzSK8kPm0wItB96DJ+8SrKv9Ib1uEkKq6TlU3AQ7pkoX+AfnAHMIE18BL5eDLoHrxg6G/uaVPMEg
YiXC1AYl29gX6H7wZwXe0D1FviJEzGs5iIWWCO/j8nqpN93Cmwqhwbd+ga9XER+tjc9GEFnbMiUT
s37bSdo4TfWkSKIWhl/FixuDJBJvLTfzkPKlBC6DG4s2Pp59jt0rGwn+HXqeCMJprb3ofrD43+88
ruO6yCwLnuPkyMYL3sIl8iTrpyizFNpct0saDSrVy/AYAbKWRustmj0JxP0ri9cf31IV4cXEVBhi
+ezOuDCDyqBtJgxs4uEbA08ZClSP+Sq5S4Jv51R3nRiDvWqjfC9s2uz3MSZrTi6lwJMilDmwx1Z5
HTFngxyAKTHUug/rWwqadHVd797dpLEFzR0T72RbUHovYN84rsM4/W5+a9f3Xgy814nJJoUuuvxk
HKr6F6sujFbm7W/1ZNTTexYFHp9Kv8tjvgU004AcDT9iBf5wbzWUbEe0mIScNmeYO7bmBFeupiN/
KbRX1Ti+adAZooZHwjcoQTIjKHeB5qz1cInQmfJALTsrMyRUhh31RycaWpgvXDrPaBbrFJ8TeXqU
KJ66dW6CD9gKdNMzk+UWRT8u1vGVadMnvLk0ss6W2Y4fep/NDDIs/BgYfvXsmQNEjrkhDToGc4XF
8sAj+AWPasvx3mnfLIxTRS3MwxxxPbSNpUpIiSdrhiGbqmFtJMyTsthBKvyv5lCuRDtdC0RC2Wek
9RiFt3UE05zMRDKQsAwHXW/jD/IQ0rSKpQA7kmYls06kNdoieMoBi9H1BuMU04xDD82osKLcsJo8
mb8v7XfScI6sgPnsMV+9tQ1qF8oQfPbIt57jtuob7EV/Pdg4GLD2ypFLJ7jeKSE4NB8Iekl6E9ZL
eQh7nHKE99myvQ0mECkIau8iMLoGHqHo4Xnq5xHiFA6/n4ZWoxR25RlQa8zY02gisB3pJjwHb4qT
yfb6ucX8xLYoHskrM5qSZujZn4dA1Dfbzf9LAZCoLP9pGHzRbO/DghJfN0k84hHICI5C7dtkzhEI
aCxQXd6RL1xWWy4Cwn/wd9NbrZtabsvpTiglDr/gzJ8Fkb6fbEY0MlY1uo/Ogz+kcmqMT+1vCzkW
sz0jB3TWWcJp7oqmSczi2bMSeGuuRWinTHcQQR1QDRWZDGItHF2xyD4Eto4xwk8RaL8YzLhoDPZ1
2JKFb7UmiTH/mG/C/r0OuTCUzCvyz9djgz9CyGy3+mJISTwLDlbyqJXN4w7XHQ9XesHlrrzhd+JU
roUAOBrOyS1wgXny2cf1VUpyAuygTCNvgwVgJ5sFrP3yRqt1zqcTnyUSOVdJX8QToOqBxi2FATWS
bXXLo+KDTdWV5mjBIvehLavI9s6x41DHATOH0PXFO8Q/X0+cXKW6joS+hh/TLBoTz5HGkfo6B1qz
zpXc/rDWZwOmnWrKhRhbg8Kge6V1Zj7zm2lzmh4RR5U0Sf2CgkMUCZPlsgfwdazK1Mm8R1msvB9T
R7tIBufDjaK70J6k1mqfcKWn4KL8kQ9TxhPoYqh5gpv2wGHkn8VhR/mGNQO/ATXtgXuFbtlwkser
zz9AhrQz3WqpprPO9rRz1Ld1fs4Enh3WNfH32hlNi/Ct8H/XCUNBpsSgD0cXD1tCZj+Z6bjAAi6U
FoFycn6jyoeF1vf9hGTQnAFKbsXWcMkxfKdNdoQ84UHOQZ7V0VFIRjgo9W7q68eAqXjlDxEEY2WP
cMse1VUN8o04ABxVuowQeGJPq5xBhb88zmSRn3ze0qdOg5d/DR6iQ/iatJMy4ItcO3Pb/8+YIXJ3
YIdv/bxLaWSP5Oi2iLwX5cnaLVlOKqI1Nz8N/BaERED+plKELr/4yViQLedir7ZOswLTlaVFM0bM
w55CHOp6uMNIN8sMvo1fNioAWWvz6y7kveYwgXb+WPmmu9Xse4Sb31eQajw6sz+DNz4K6v1ZPLYL
Lby8YAhsTaZB6zzLnOZmS7ZqPzVBpbxdMYdjbNvpKUftsjB+mJ3M1h8nVhDBXhVp918zxUJSGZnc
GbU80dJQpROrutebIax9GBbYZg/MLT9xUn7su+cxHsY7KD/3FeGMFrLYXA/onXyqxSZDGS8ioGJ8
nBNK0Lslw49uhUaIfxXsW2/NefT8ibHWk5qb3LSKl5rqtMnOWaEzLxAUXvDez+SW0Yr1mV/z7Y7Z
tVOSRnWH3CT/mu9eLGz4MkSXIu6E4o2jTpOD3iBylhalB6K6I2NDBotSkhsTlsp3rpLsz5LFqQo7
K1gktWwmsHQRvtQfLHpZWnlLZYs15wmPCMXQVQ9VAIcyZbP+X3uHcyMBUlY07zwqhmVnsIIsjQqr
AVNZIUBQdMHhlWYNgERLT2azsb4uhB831cT4mUn6dX+jZos9rwulYFB2wkSqPCy19jTdOAsqi5fd
s9t6LMTnuTA2Mvns5IwctkT08qg+jnAQM1NwLeyGq0mrhdpMhT1htRG9Vv8zTtIwXmstY+SLXCEY
1FCry3IxMPKT8mFKUd4pZ4wNj8b3aQcCXOxv/cww249IO4LEJVVWrZu86eQUeoQU6Prsc8UmNZ6e
kQFkTvoBQKQf8qqj+DKqJ/TtkXEafTN3X17hpkkNeeNE2hYZxvn8lQFxqan2hXtc862hLGJce/jZ
kglxh2lQKUP49piVwxjSZPnIs4VhAkNNSIjUN82DWZNnPL3Px6VsCqSeAt5eZBpwuO7XGyLCRlmR
yNd2omyvibZMEQ4pGFKP3JM+7KAi3Evqz0czpE+MW0tUVYWD1hUUDC74SHY01UGuTjZlKzEpZ5Zy
o2wCTA8+DGhSqjG0vLlsj6z6hdnCfaryM579QqWfRPcvw4fj//ggkUFergELLYxKrEsIFCA28F6K
pmc8Ycwzn/VSFmSd2tQ99tYZ9s7hHcJN+D7nrsoDApck8QQOS9xDF6Uws0k5hdKNXBF8qKSsY3DS
kRG/zwbcj+mif+H/YdV1Y7NoEd8w6utdmnODBBRUKy9Alt9jm4NsJcPuR+dqCfhy+C/EUwKpqFc5
uc5wjT/LLXbMfoIAYIw/TX6s3gr2sz5vgMkndE06QwupiszBMbpdCo9uDphcFOHw3g95blqSWFrN
/cW6fLzQQ3Vw/eLgNrhxCnZScV7Cm9Lpnc/5caUvwyO78ZwZVq3dwEfru3e76hFVpufUT2p2BW4w
FJrvjPr7uYmq2h3SGNEc5WTMWGCSThtvCyViKj62gy+qaHU0CXwrIl2KEGsxWCf27DO6qkyPgURe
8Oln6s/OwoWKWe8Zy/jMlXi5HETFiy8/nSowITvsFKwFZoFOMicgPAis8ARE1FElvP9pBxnwzS/N
PwpUQJpssRT5CbX7zJNMjYwHdbVKloI/mGpRuWlsUmriIHvxYTqJ5AxK9m67/latHreyEP1avUbX
mCJfwQ5aqv7+c14FCu8d86SHiB4JZcxA66I2WZzF0P6IF9+6lN2/jyghI7++EgXTMvBfpLf/D8xv
SvTgVltXILIJM5cwYd00a7eQllETYM/6XuOJ/kRXl1hZU4q6MewMRklg3ZuhUKl1YtvssiqJTyB4
wQ+y4nVEkoZMW76gFV43vGqPlqWZzKe3riqP4mkY6Cmt+kR3qBVzSrNv2dDRDJWhBhxuxm4E+Iz9
m8ljqNBdOruNeDteNhH+BCkhCBSq43HotZSU9/TzmN1cHTYYF6/Bjb2W/V/t8pNbBOSY9yvjvnmm
hcE8+zIg5a1D2xmeglw82ioluuE9eR6lqUcDufOkfZjGNyW+XLK7A+0n7pzcxfSv3gTA/HN8VZb3
icrH1n0aLzYkzN7o+Iq8OEVjtmJidr+zvSvCesFJuY5LzUQ06q+RZ1ZmJpHxaSnjexVwFeXgd0qO
57v2F32fTEoJSmqd3SvMNWhG7kJy8aQlpWLnQ6tEoIwSgJ4ZO+KY+hrm5sYqa1M4nxjPVJtev+mv
7quqr3pTauPvHqUcUE2mYTav87wHy1ENDA7GvJpnPLTLgnMIGq2QMb2gph3dsjn/tUxDFspaFkuO
1L9rvV/9lc/ERubVMRmaalfpN1xsgaBulwFvY+HUhHdM+AZauhoXMCkB2xqghAcPblcqQNeDgDU1
hwplbWzZ/zCDUOlNj3Pg8jW1HW9k48ScAfKoc/bsN4l5yGfy1PfzxL69e5YPAeOvTRgUfLAJPX6B
lrTLljEsOxbCWBkQg3HPH8t9fbOlJnkEllslHa8B98kW3n1sQgCHKdDOEv57q0OCk0TWl6K74rD0
6SVy2oq2K+es/DxB+Ro6D2iKI8sXyY52nB1ApLdkbeGM1QZXv7XP/5Bu+pj6xKArrF17N/mLlCNG
E7Uzzk0fK6ZWxHNUI9CC/EdXioo7/kGIZraZ8T67nSuQjDaE+OfTEgmgxyflOh5ge22P3mnHpDin
x/8H3astZ9gDPHGNfcBJQmSgVADA1BJCIVcM3ONx0Veo4eDUDfyfUFEnivnF19h+KFjpd8YRBEnX
zo+VP4IFEnlIxRV2Lw92eVZHxXP20Wtnh9UyFVv6wC1E5IRUNl2WglIWwW/UcTk6RKLbh6OlGJuY
VQIxMq24rDoBV/IaAsNxMroyN1n5+H4LeONNkeDPGUIvGNtc6+mTKfuzSMyW+YG520z4EdybjRUx
+qRGYdJl0CadCgTdq580c7/mOvyJzzRzhINoePGxm9PR3apurvgNpzii0yhsLYyxM+oYYeWiX4sM
zErFvXMDrqMmcsQpiY4INwnQsXXRxoRJ7gfio4dF40wFBk2qHwfEdiTJna4UH/Gei/nH6wx1Tl1F
WNFHesicsygnhlspyy1FaDOKBqoc5OnmG2x99zyKFvN9RmhgsiQPra8x6++jHH2cUlfKk16t9gYL
gxCoPEeXnHepOTR9BtcOZUKS+dqXrpVzD/vKaEoMQfVlstrsNu861543sEo26llJsVWWnZiTma15
152nLxAooq/z98z19+QyV4xPcL8GMPe4Z4+vWupULbRvCyox9auHNPEEAscrvEqpXIKmp3KQyIUO
QtEMQ7tZs1EIsrwXeI6lVnb5XbsPupCRvjC8FjOcmKaBHwjXuXmvfMF5Rjc8ZONWC9S36c8Pk9EN
2QwI+3OLQtnpvY14zfMawUa1H2xRdUMJj31uJOAufDdKVv+tybFxrtrt0tS3KYGQPg5RGExQX6tn
LcNNf6/aYUQrnA/XrDN8YCvZKCWROyURvFHsWc+oRM5LiSD1la31QjEBpNP2sGHOvIw6XOFQtyQ2
WfBDVi0F26pK20b+WAcaTY8Y57h8EPxQLV9CFDUNhnVj7bM2rjW8kgp97pgLRMRRMlB9NNzVly/C
pst+56+vU2AyZef2esgJlvoultx8+EuXfmSCf0hEcj3AuJE1jkTHSwCJxsiqs0+CyMJqRLrH1qZa
vCsKeIjiUs98HAxCunsRJsPSeH0cYDXEEfnsdLtjbmYjE+UbwyERWt4hq35vMZ3IBSL5jJD280uO
OoZcP3S+O747cWXIxp0K3KLC+SVawPK/JSaGxbmLIym2VhjchdE7+lnUWjs+CgC/GjPeC0dB+LI3
fUnoYSULMAvWDrxaEDFGY8xHr8/tbL5mtb7usPsGo3Ku5waGHELPqkKkHYCz5l6LCuUwgWJvKva4
jOpP60QrtnAq7mrKz7qVMEmOzM+y+2BLL47dB3jOJRuUMvFSWc+dEhZ0vYBxd3NAwKqoZliq97N3
whf+oSzbelKfx+CI/vT6EcNfJ612Y6Kr0ZbtcqGmY1pTGpH/3abkXH0W6oKu8mV7cOpYJJBFILdH
NFbM6qCw/zf93WFHnxDZom/kYGL9i9bofTWEDHDyhFqOFHpjAbr5j/cRct7hwffMS8arnpetv76s
fsG9HjhDloAf5wWOAH3P/N6UJKHzUdvOcopbGcrtJHI7GzyyoBGC8hW5gleB354Dfam8+rPfKlgG
WUN57iwFSyIK/IzIbsXEuLkf7nmF7AgaxKXJEZKIc1GseGRRfxUT/EW/XT4c3DDKkKVTVEHwRAFH
0uBhojJc5p1B1xvJTjDNLKBcNoI/b2jjMK9bDs2WmJghWkjEPgCQGqCwpj9EDSCtM35FZm1iI7WQ
vfRU9EzL8wVUFXbA5CijWrEW73nPW0cUjMwjVZnFKWlXjfcXKmFvxbHTt0q5nHAB2HeFD8cbXSlB
Mo6n+48q8edN0mL6SFIXd//u909q4lnGrl0PkRG/kXGeDZiDXPDJMWspRmlN0+MbxPrc/BJcJ5H/
twe9eXDDPqOcRc9wOWK94fBSmsbC/dAe1mpPkThQ3rJmmzMYu1VZ/He5erGom/VoLlgR42ASfOzB
d32y/4O+nJJgALeLQAxccNr8lpJkD2dnvKn5n+ro/mMn6SrlmWw0MHpPpGCVYPwRyKwvFqVc0PP5
UV1y4slfWXwXJFrwvjOXSWlm2iGwtCf+sC6cBIO2brcT9E3l+XBNAhbf4fA4WL3NsLMAsY/Qn8zQ
2S9CVNqD5CP5DUqX5EtYgLlPyAt6Sxd7njB2sSHZZb09EiOUPTRP++7jxyzsYtwxDz7Z3+x30mF3
LVJtZZhuZPJVQMpJh+g92uLbRaERvS4SC+LKTvrmWGvweBHZ7LqYIic2fW5IFxkS4Wx/GMwEWqLw
7lExM83n+B8rKEGzlQjkWBGf64+knRPxVvuS8fjsysr3Og+yEjZX3OxGrempwklVXYTcTWI4dbR/
pCRD1pFRkHvdJN/s4m3DwbBbcBslBJH4yYSF7dnXfjPNgxCrs4YKwvdKmWSGhLRCXjfRWypyH2zi
cTYQwE1T9RLu/7A0cThsWPGjGd1P9Rf+F4F84PmuvqM8YjMKsBSH40eGb1I/ihDYZobe5ErqNSwZ
cJflsdY5qHLXO/9fuJm7Wvx0g65wRAzsGv5+3nroJp++UPbtmsvBbCNg87nnyRivY5/x8CDtZ8Jf
I35zFK9zFzvTV4xsdoyjcc8ESMrTA8DlhdOp4/Utgg7d/EdAf81xaKycpBlXhUsxAACJOB44iX0c
fbIrQqFigzLQOxZjvPrCE/iIIszmQtKDyi6/J+EnXqPgaAStbY1twxhxzSoyhKXOzYX4fN1Lnz02
eQzXbIOkrn9pXL72h2pafORak4onzx/yBqyRsuBq8J/je3utr9sJTnQQ127GNrBd6O4thY/ZzITk
KUo9pSlj/q2jpWOh/w7iXEBJOJ4uPolxnIJLZOH+bTjT94NATSoRbW7vhpYAAeThC/6BYArS2lVD
AT9RhhdK58AYacRQqvo/L9dKnY6S7HKSjdjHtA6vuu5Eu16dnjERZIOxWW48SC7rjvZUZup01cdW
IbYy1Uzm4WYWTTbTPgCYb+uxRuG+MJjfxNYF5g2BcBr7H1xl0QC3+SRcHKYzbH6WKbbzvrIDJwkg
rIIoHCUy2JfSKxLCEUA9p88jzfoHlQflfIh/Mxhvinpm3DA/n+5sWDa2eoG6Y1V1fSA8HGaWzgJJ
MRuEXh20yNFOWEuCrltx/ZdqT0NBfKiq3shaEaovq5xskjX5iyUa+XMHnvwQr6Y6vJS4D2GuNYZb
h4CmR9gKPpAiWdNKrOyonIzbibLtKehhWj+1JOBgEaNTdzUGkFwCc2ne0H4GEZHqBKjXLnH0bhwV
ooxu5zeayVvq4g0rvM0EPVBWD1HbhZsD3LdwHGR/LIWI79NcdswUNt4/GVCNswOK/AXKckCHdM8+
U/k08cC7VLGSbBAvrQe9tGpizW8NJjeWV5XjyErGMcxufQqZKJpxi9CqNWzFn/zZednhK/bzwhQx
a/hpshDgp5QgTq9WV2hrq/HHD9Jc95d5EDsRCHmOGkLUaFvXTs1VIC9RKNyQ2A9bfD2Jf3Uq6mxY
bZXDR2YJWC0bJpz0rp3SFjEWPPHWn3Dz8JlsEwGQ8vY6GrwwaeTgD6yx1sTAWvQHn4sVnsgFADgT
g33OJAAX1c9G9zwYPzMQSb/QVUoVjx00v4jBS5i3dzzqa1Dk/MDsOVIzC+zOqAMxmgUqf6b8fP/3
R69P1XF3mOc9lB74J45ovF6WETnu1TKktGpdhfHPL6yOBJYEWOT01IU94RVF35ZaNvCqd6QzveIa
64reC+x7ue6GYUw/5HsOBTmP3G2lOq6frbCs1XO6p8juydWeZI/IHRk29jCB6H/ZkdaUOADVprCo
ENv3FOZXL2hPVEdrzCnb3/ekxXCDvRpsubsWljbIOMqOyRp0Xnvg4iiEF6cyjj13qQDfvuOTHKGL
1ztu8cdJzujnlbF9Tbh7RGKF3jMI+mn9U84qR25aLg/dIGQ42B7ZTwvgriaQile8QJhgCxMXFIzc
ONLK8fsHw3l69WWbE8A5zzuHmNQBDgbELmgfaduzUZDhdqNApHFGeTa7HyCa9B4OeudOYtdh42pG
qxirVum0aKYJMAxe9PZ17JVndPXR1vzuyXucXRILFFOGnUE58ISJBuHN9I3J//3bqEjhRanzTQfM
hKr1ZaW2Naf9FPuIx1tSE58Ms21+x71B0r02dscTpD3wH1K3lL4An937TQBbp9VpfWGna5OULWXN
AfrWSkldARmSc4bSoEJhSC3iOjRtT/ngeNVbQjBJp3rcD5791aZlXrjlp4KNMipKfJlDgogEY8dP
60NwiMAJNTAiJvwYvhuZ3//XBV5ihPIgrp9kHu53IvUnXpBt34zZl1cc0WDvrXD6dXQIRwhD2PHH
mWiI3NXje+2e1M/Iq7iSgcngiQ7hNyKaF2UGQ665iOF74nU/VuCgaG0pLBb9GTHb+K28ZEiq5aL5
FKgZ7jI5I4Cf6D3pPRJWO8HgpHeVQIs+0dHCQXgWVe6HPJ9WZNUFa3YwtOFLDAGhWGdTtrrX07+R
tnuwxZdqWWWBSkhbq05UKMnTnzUwkdqG/dTqUSI6mGvaBNQ3AtX43Amv9FFGv7yzN+x24NmtCdud
xotoCIthzw1gdRqZSDNNblo1X9rGZ4KTNdwcgQ5eUGbw8+/G4t6M7S/74HJr9aqFzkmNSE1zP3QY
2VERTD/1kOLcpAdkk1/KDPwm8/wPJ2rSsxW5hWnzMYHQ4NZUo4AfVzYdQoaMpLde3SgXylE1vMfy
q34vOSCv5bzOO3xQW8yZKwK9epdRGcGeevLGq/EFNXkkn0E3PKO4NJRP7mmw8c9c6KXFmV06hmVq
t1ur7N2M56oSC5rdTNbvb6JX8PDySSNpC3NQj+kWmkPMAbMnP96byppTUzFA2YuAmSvf3HahL/65
hgYUPCOWuAVfJfpdN7qnyhU7c0aENQzSPZo8+FWFs6K2Iloz2KOZOL2KMfOCbYoq5AuLpPulhP2N
ynabFeKs/OcSwPnG5UKQI0CHQ7ZFiD8V6Lo17ooT6dm2NrDHUAAZ0z6Cdha3aJLlYO5Tc5eFmbq7
UkkhugEMZrK9PYiaPDh4NuX1t5kv2W9pjs28V3VCWXiFGqKkN97pmC4SzkWzzqAZJyERJWgzxDsx
PsedZmrJXyFFE7RFABVfweQwXcEInDAO+uB7Z82DOUCbWIaG7d+8zIOmrZGws5gponf+d3qJ4KbH
9Wc1aeyrV/hnF4SvQf4fNDdz5C1dKRNOrdSzAfx+7ErJkwNsjTwj/UCp/Oa6AR+XI5z04GjGOAAC
swaRzVMp6pQc+ah2aVvRdOmd1hK0kRh91b/auoBOvqY1TdzO/vSj0UkFDWrz3mDGrS6K+yL1GhIr
yo7XJZTS9h5PQpCHGBsPszg985oP/NXj8agz+cDhA7sAHvb0CivSrp36wec9T7sm1KXzw9OyYxc/
znb0g65A4Ostb/rZYjpNqntKTklgnK5x/DeSrSY6bPGnojn+x8zX9MBwuaJS77O1f0hzq/4YtDp4
18N5c0Lg3XZgTef0+MM8xwI4xUQgvjgAERdH+36EuAknS0TlWCLe2RoMK9J+NYAHSf/RQCsbUAc8
EuW26ogannOv0sAFTWzw9Vv/f/blIC1iq3jk4HbkTIqPS1WiLAP1bKrxPalzfCpqSNHryp5o5iP5
p26+6Ru1Kp/DUc9qtbOKQT/gtKILWnCu0yAGp13j8EQqAGRagw7DEU1umrgzmSkkU1TUvWV3Jup8
L3/rMxRMbc+FtaKhyTUHidhh4ZBxEE77Ph7Ko6bRg/X7tB5VO2PSR8dyz5I32WLGMYW9avYDbeOn
zhokEI/SnEkj+QVBH2gFjUaIJ3PzHanKXO5YFQ61yIDeU99HYWLxBnJvf/Y+8FTw4DMW/kH/ZbK2
g0TSGM/kEfpC+f07ebAMNay/folixUG/SSioJnikkimbrfCI83eRvcGNxhBo4h+a8+GZrCJ6OcQt
Mwt8uY/mIj9Jmv91jYwj5Hsr7SZuV1T4ziuywm/egBRWLUenEPr+IfiAo6Xq8d7psY47qe8XP+0h
vt1+s3W7Icw0nsPqxPuK3a4h+NXHv9Q7ZJcWgzXvUTSpOMr6cSDQwRjsqVVM+t00+3iztvgN9YV/
HESsSz1ke2TzxSQkVYcBEv1vzk3qtryR1oa1Hi29Um6UfHd7infNid+eUslyL4Xue68Kcq/uEeMI
yub9KStIEpQ5aG1u1ZA5ctZZV7U7bUM8KApTdlysoSmgMCrlStRDxAyrMsSUKm9pCgTv1gCHTRpV
dfeZWnfCitQjP0KWKe2Y6eNzhByJH6D0zEJaWC20VbxETbFi/ctf7WJ6lzNIo0DLcgSC7rO0Nrwx
vcOIwPffktQ1hFoLMuOxuws4oK7TFq9fG+adW591WTF3Fe0+61hCbMo8EhJ2XI29xsxNxPnqqpyP
SI9aU6ynvfUHAEexJjdV8N3slQuF8r2jPXNkXQSogMZNBog7+VoQpzCMtdJanVXyg6zELO+IDhE6
FBNgEkK6l0vEt3RsyGeU+Xqj1OXneroqIJQo0O30DioctCA5GZHNulC0tFoz+6y6BcvgSDnRxu15
9ZvVlVjBjGrhuKiDRgWBh61uZi4x1WalKJtLGZ3PZsJ7TcuYG6LIVG4EOQ3aK5yLEtCw6++3jbMj
BY3RDnCQQPIHDkAYCibci8l+7snDvaU/ubbBFpSch2o65vW3rtKAXzBAWBHpWFFE4GkY7mb9gnoj
75NJzJXNbSoPTZn9NTbhwTh9hX+mqASXEkT2Zu/KEDOQaDr31ASebfEwdDcyam2t5hyGqfA3Or2x
Krkr7v7GwJyHRyg+iT6rrSKzW7GcGd5ln7se52YL9pa7pmge8Qu2SwT8xOXUrsZtvo/P9B0tlr9V
HkzxYJC8qHIFjJnLsYpqqiiGSUwk0mPFzARvslqQbqKYV565eT+Y9KBb+Xm6FV8hWD6cSHrEa7UT
990604OvT1k9DvYSYOc604jUQwjYT9XtmJ+Af0+/1AjSGPEdj0UiqE7rp5CufCfI7KCHjPJatMJc
mBoJvJZ39g1TXr2+CdxWppA5RkWuW9POdgo8J+n5cqmY3V/MEO+7mejkbaTLyY6lIjQYJgB/FvW8
+uHSCjyez1rRu6oiAqjkuqjJaDsmA+g49koVk1hCJTtes6T6b8KEbviBQBqHrsMTG4HzXnn9dhzy
v7/S849Yxee/8EPzhyt8YUIUUGHL40KGZ9ObSMb4NBa602+WXpXQi6xxdYMinzamKbzNwJyfaOBE
gdlEpEP4Xl1dyh7Y/vSLbjWpVVzOWI4VWNJ0efpw5+RLyxU7mWIYCyJr/FdHpTeD5OFXan7f71tm
9Jgs3t70OmEVHbTRqROKEErUJR/ASQ6Khm7jIrhSy5175KG9RRuiFQReaOYfrRml1NKqbT6w5P2x
wmWQqJPeSjqF9WswVls3l066d9IjxNLuIDL3TiT/sTe0Cc+yvszLk8blpKubaFwL+M7gGzBnWjnS
/UB8WxQ7eDAR1HLq12Aw5CSgBUnjTRhR21Hg/VjgbKkNBW0d1RGPd5OwnKrz2PkVSC91lZ1WAq3N
jsZSKR1M+H8gmaKA1SxwkVLB4g0dkBJJ7ZvhsMiITu52k61gOoOpumMz+x8LSlq7GLkFiSfKLlR7
AMLRfe1aMLG6WEfirzr6jOzO39+g5oIW2rn5goO09OLfKH0j5W+4tuSpl33dshZYdtbrqtcWWMNl
dTVt1VKUCiuuM9D61X0mQM6hTwYX/SiUXFR6tBX9/kyt/ZAw7LoIcgC+LWF/KrHID4RgXrJywEuh
uGZLnxXYX81YVMHLiFZDnYCG1dtmRns3w/X4lO+nFlc7RsgP1RYyplu6SOp3Yu03qDNAMabhoDZu
OjFXAk0M1SoLaOQGcz55I7+hehrv2thzwd9HIlaK1CGRtou/6KYYvCODmeyNS+BRrPznx+taaeWp
okl1tD68Svo81/F6CCSscFVgf0VKTos17YhRXiqNL1WNwxdYEAXQa7rsJiE6pBb0Z5bWtoH19Tj0
defCZJpYQNXbCLrSzt63ewou+blEB7DxfDcfoVO++KJ0DubrwLs3IXzJFKXS9AF5bVSt4/iaTv9O
Dk99AxvdJPIPkOTKV1ryOa6W/lZ9W+2m3whnqjvqHbp3zefbm5Ms8Ir6/kFl8HXSPjk6VkvC/7zY
D9vk9lgvGVHtf0LCFCnWIxZFlqQzSxkmiS1JIRlUlDoUeUujfZpYUvnjYVgHtjdOiF/NeadUn2MB
mDvsBefrNf/ANZ8WR195pWblfCQjJdtxhqbwbtLnN7agdxMgk4CWHBnFaEFLAs7LAv5mYarRnYY7
YdU+sH4RxilclivgnjAs4HiegAtUNxvMYH2uX6q0tBAFNsZjV+wNFoOlaSMHHnNctFD8qq6y13ml
CYBHhtu4CoRzAriySa+AKLrliliflxKvhj1bR2fSG75+/S16Zfs8W4U+qCaUG/QG+wJMGRnSxQWU
aHHnR8p9drUYjwv9TUbM+u4CQTbviGMxdkebp3fg+OBDkHQHhMMSmwvhnLVNlJ6vPSBOjRF9E3YR
jNpL59i6VUBzf/x6QP8UimKziZQ7uzjcPeLbpFMiAOAarW/Vpg7oxSTQx5N/2k0k++GuR7MfZd5Z
wkwtaePsKNfJMzMO4B8HGqpPJj0muG3kVJ0FLQbokzmR1LmfhdGT88A7ShzP4yFn7/CO09civUls
TIuTksaT2JJBzjWzLGeoRKDBgUVYobog1LNgSHhglYHncreW9c1o2waAcOHx6Bkvi69G6tD+KpZV
KWzHzI/7lj2cnMIQg/rZ2Hd4TqURiiQCtuYGs4OETsA5kGkABZ1BjdDBYJroO6yvE61wo/IlLwTB
+VxJLRK4qYLT+0ikbLZGv1wvIcDGHiXbi4vny4biAiN2dHh2XED4rlbXIIporoCpMKZ0gBiK05VB
zbATSABYgtyKRKgnYRwjffAa5+EZ4/AUHOOvvDU6PeovTJIB3u5MC+OJFhJLMvq1ASZNj8oZyirn
l1T5m0jYOXE59RjCgODZRKETzYaff+NmU2mvEaAbF4dzhB4opzox9967Ng80dDvo5Pa5eqtnyOBM
0kACPuCh4zQpEhPzGGFhZmbiIADBC/V/lWg3cUsb7EE988algZXSSQIrSHT/e8jqB6j1O0cjiamF
k771lN6IubO5REIwLzecPKvol45AtpAH7ytWOZOcDOmuH5R6AXo6yMURrau2+e4BzNYNuSn/Flz8
qpNBXJy5CNd/ZEVP1kczPlq6PoloFHdQfrN2R5a5WfN9u5WZNW7tXoH8B1fAAyIDw6uLB6yKMoUU
iA5x6n9RqKD1f8Sr56vVYVkwQxI9veNv6Cq+Qpf612cgRb9X5z1QBg8LjuH710q6PWBFPbq2vSE9
PBaRxP1N+evKFJWtgjyUejva6wH2SAuOeHTig+gaWswx5xI5tl2iyNQ4ez24IyzLvAgXB/uRiKdm
NFJG7BGXWpkawsi/t4dQamEW5XVFW7aa06jHOPNUmanJL5vuyxjMshOu4tzfyghNSwRizurtIqW8
uO2AsU/+zRBLUAfsdMD/oRTDpBfqNspglmcOpUqe8kkmnyjLEZnzT6LY8J65NHEiyz/zrUI3xuxY
BH3VgVdf+WMzgh3OwdYZtrGD7PMGcup128X9Xcp8yJiWOpiWa0sBJR/byAwGz7umfqnMiZdksv/C
mXMuON8f0PgaDKX0FedDQGNJXFn643AO+sor/mLCcJ4EAxst0kD+rnyKp2CtpdHN4480I40H+3Bh
QEMbgpf8XzOgQpUhPV9FKg9qb6+slKGam+TATJ+zcmE6CfAQ7Nv9isXdpgBAce78M9Jyb4jqi9Sw
PeWXxY8Qi0palzMBd9UAisjRc/+TVZGhFqVZs2SpG8Ed60J6CKdi/GvJ0ttbIkUnrGafQEBRazs4
7/i5fF/SPDKtfvHcupbBggZnEPvPY4mEgiWg+AsI7l6HSfuO+hyC96N7Ufu1g8tMndHIidQtmwYG
gSYNx/eYd5fBlNFNrtfn6Ci757DmkI1K/Tsi3a0An4YWr8B815uJuqQetMJ8yPpE3QHJx3Ka3DvJ
juuNHWQ1OGQ5dlf3AkunjwwU+JxK3eXvFzgP3mGqsIYg9qvDLzEXfNYzycdsghiPRaMrgLFH0/oe
sLz77tmDPixUwk5QuE8+J2xSCR9lUCupQXX61BwdZUEzmbWm0C0Fe4BjCCMAmwLO5lRLHUg2MsyX
+e7IqBZFKBwUiVyLx8iAGjnBaS4+qaq3E0JjYD8PXeFlqJq/lBRzTZlWd7pTG7KrGEHczQBtdf4v
rhZFkqRhBGXF9TX35Na5RrokgHfVcJozhgFHJ/eYgki+PgIXe1vaZEhBco1om2fT11Nyub91dHPN
/+oOCA0FQJ0gDvAPh4T91PJsNVazs4QMH67DKts5MOaEmbiAb860b9z6dt8MHNqljMnmYY49/Rbr
S6FGQh6219bjh5Rh537l2iGw6WmuomI52WqXFUwqNVak6aNlaw/L0/jYT1ixDrrwE9mgLBOKpyPn
3rwfnKQAYytHavBY8WK5sno6wzUQJSVNLW7xxmcKnKjn66jSju/Q3kzH9J34suemfUfDChyaS5zX
Xl2n6GQTit90j67mJ2uEfBvUva9RxeQMBBfKq06vL6nBZftG3Dh2/21CkgmbLGOv9bZDdsSGLM1I
QBk4vc/gIwc5y9YJ3DsUJNdcaupOZYEThlNTC3g9Bse2Y4lJXMMGfdAVMTqSRoSJA8WHujwPikBa
4tu2xYjgJ+PdANFTjfgJdpjwSEuVLBu0CYGcGXj2UsVePbl9QT3VLgwJkQC1gqXdHFQhQz73N/CX
8rDlSp08T3wJfPF1zQrcetdeTOBG5Vygi+hH4w8/LCoAUMQt9ketiYi5wLhZT+BCRDttoaEnsmJs
PgBhpF+446hRqOQzwBRWvQ7zlsgkTjZ3/5nLnQ80vhVWbPcq/5pIvT/+9RiUGrmyINTisJTjuMIo
zy0Jw5yNymZhw/GfJUFoKv9TN0RKPi36MVMP+DatHnO+A0gUtmwd1F9QogMPRrPBsCRPjVWr4GdD
8C2Z+ibm8ptQJ7QW4WQyKyjn+PwEg6hF+YlZXYokNdzqWTnMMGf9N/quBiqyZLTuSD4Ft4X1j9NP
aRuD2tDr+1/PqIOzOR2Ky3djvMrt3xEP3WYesdV5Blly2MgES4gb/uz/YLMQVjaSlp2uDqXhrSNK
wYx0MGqvAfFnorF5rhW5CVIfpZRifODLeJ7GGRqPSzJruMrTowY0lNIZbLri0jb6KJI0hmX+xjZR
lTLjdGpzNNuUP4/XbSEX/lD0tI98rNYFW8FLSK5SayWyO+8og3EI8+CFqNq60PcgEylsjWudaKUT
tn2yZswoaIGOe0N0kNX5mUUARD07tjiW5Jzgb/U8WKDYfkkoc4BFYAB8X/L1i4gDmtc8MQ5y3/7h
HHKu7tTZ//FFjLwfa65KDwzAaMkz3aCPfZzcvARMYS4H6G4CcSob4btORhuTsDYFRB4eRI1u6Rvo
tCnSr/vq4+S3hhZajqum36FW06W2neaUsXsK4DkqodeWQJVurbHQeYbAFquX7fbRBErfx2WbomJn
zwFAaGcrEW7NG38VbekahH8KmoDQ3Je9YFkxe39yvugjr3p1LNwUgX/ghXbpaD5eJQF6NfaeKCQA
uKRy0sBJOMuFeIFLk6eHSbU94sx6a7tlHu+MAeZm6wo1HImQeiaq8Qi1C0rctzcj/XgvCLQcj/6e
Yl6Y8PSDZUjHh/itfK2ohevznXnUMe6IkCEn3jQbTEj8BFAR4fXjyvvbQ5G+EdSIIy1lh2nwLMnl
+XAnpb6rUOBPyBsh/QmMrxCJAaLxGb11gA7512uUe0AajRj3xzz8lAjVDosUBAlvnITvqNXk4th7
KajMkSJPjuPYOtOdBurrtnyQnYhB/8SIvgvowSJtf8hLGGZ40MFTB6UXLO3290e7ZEN36L9Odhki
AKPuz4udR4hDTREHV1K/RLZzpHb7Yq4uGrB+pYl+xxpG5oKDBEzrIR0BnW9OQQ63/FB3QHDZaGtO
eT7WCYAekHtg2MKWlFMf5T9654fI5fPTW/YaYLvRIczdTeQkmltIbfPtRm+iu1a8rFOKRGWC82SM
5Vtxc8kSNIxx4HGFh7gtqQ7KijTidENLScvkgar7Vf++SnbQON1iYS/Df3AAFcW1+NuvQucmnXHX
/SYqoA+uEX8+tiuPZCAcUN7EkKKXIkJTu6B9d+OsiKHvo37uwJYTsBRcCybkrHtA+QIekTSen4LI
YTkOCb32niBdus/KJBwrosVcv7KdY9ujUmFZ+8LGPQwuuJSLvFrF/tZY/YNzMCaThRaQWplFOFXB
j0rSiFavrBT/cJAHlQnbCxpjf62ss0SEwV6ku15k26/p9NqETVkj0rgNbcCUfsXYdOz/it3Wudi1
hOgYoTGpkt/BiXIfhom9hICWTn+6U+0D4zX+zN54ymwsGjrJ9ZAoGh7HdPExaONihEkw9QPdBRGa
U0WVn8jPvmBtmCnWmDnyZW26ex7K7Ybui2qs7hruv56VEh+ARul2byq0/Rfkrr6zUl9FAyO1NNi+
tZb3TZOt0tU289FSXbdz4KOf1WWLXpwZiqUkybr41EIj69XyDWhsw6teP65KaXZVu0oaoeqzMW1y
3I9G7WWDcLOp5ADJGDf+G9lHHQZrWA1OEjCFiESwCfubwKEldryiVOYe60bU2PkJ9ULu0xg3W/CY
lWjK/3szI3UxMMklBPxMLE41aqDJKFJLdloylo75kJZCsd9YB/wdZlVdROd4Ck9btu/c6VrgCZ8D
a5d6lmeeJXO0LZF7NfznDZAT07LwozKUzrOSNx/px2VYGXWmSXjjTk+nvV11VCl8Q/bZIfJtN2lC
8Bqc08GsGBN7rPdUEhYkEIWE99Z0xjt0XaPLO6FPm0Z8w/JetcavFYnvyTxW/SdR9PeET3i6g0PX
W9NnXVQTZDQh8bJlHdfIAJfm5FJrt86uzegV9AozuMAMqHrgjkK4XqDNo4NcbyeasxnwxaWaQnK5
wkX+VfzMGyoPI5T9U63+LKQ/SFW7c5Hu4mZoPnmo/rFjDBLO9+CivDqp2R2OfqG3/UhmoiKu8Itl
GT8Cwk67vf02IsMKqQQ2NzDRI6uZBxsQ0EhPzxiHfVAREK4l2EL1c7rjLOLiV/Re1VmIWu1/mgWb
AHXsEWisP6Kux+aDv0Xz+pdA7b2PqWsJsaHt7g0pTMel/jbJv9UyGOegcglyoVxVZmBY8lK7e/pU
WMdXpio/LhJf31+WSwXU8DDs2s7kkyprbHLcku3q8J4TB//zQ41buzDfpDhETN7nz+1RsjnAQMvx
JVQEZNcsSJCuHh/vk2VYWZtUv0Kq1s38IGPOXG4//tvtX0EZjOWAjG1gWnNfCrIne1W0UZJZd2ot
MmP4YCjxtDKEtN40JgldmiawdfCYhVHeEJtGKttt+mCxHMyIWDPmKYh3zRt2RyuvC7fDFJtEopOE
tlHQ0PNVAp2nBKNlt4kT69uwZuTqlM4g5q0qYTzKzkHUa4K8vkh2mwL8fWYDhbeXIgJ37J9qQjt1
8XJ57v+1w7VM+HUZD1ILWNcZAX0KeWVehm5kgO3ryT0kPXSR23U2/Z/nUvcvKqWC0d4HMP5A8bT5
x7M6sZrJe+xOcj+0rdBYzwyPuGB8xSM7PJFKhqOpGeox0akYOE50HwJHPWEY6Tp5i+1k9em8XO3p
QGDGypAizGITpzwQcDRPihvwNup0if9xBP2bGLZGcFVh0lMs7MLuCjkKiiIshmNMtH4ge+qHZqhS
yv03Ta3Wc60gLX2v8YXaPgRn2tbjfk6XyYZZNL8KVTW9Oy9NLXs3D1WMMHqPZZPHDf7GacKZmCey
eof9wZzghF35miU6im/FFogMIDqMWU3UCJpLXzdrJLQGu4CA2+u62Grj5k1Yv6WCvC3VXbdGMY9Y
0iAIRylSeNCmoGzT7/rkS5fQ4HMsYOrPM3UCR4J4cIEMsyNMiRZQIaJe4kV/sfKPsUuhmnQeGZvX
BCtSbQGkTxH1ExmAAE/bZisxCadNSaAYnbaIRVwX/U+vYgZrkF2GONG5tUjHiJllKUCwIA7BWENE
YxqGYv2NEg8lb9XYE7AMP1rTISdH9QiyVYWn8+kDqH3soaP1VLwBNfB2mM2L80XAMUz8QMIQfN/Z
hWQZ72QGsasahQb0bmAvZrOcrAymV+VKqyW5FY9P4uf5tuBK/+I8j2B4NDdnDx5h7sYLuTAaGoav
MIkqmA7fKAVqgRg1XGp4YDAndv9IHzl62aqLvPJLdaCrn/uBi/kMCBJiWb+zvcBnFEXswbN5wZXu
QYekCr0yfKFPRZnRMuPDbHe9nD2GMzfwCrm956uU+5mrnLyJCDW9gXLVayK3bLrr3AQgZjDWknS4
OSbWpEn05gKEEFYFt8z4g/RNNRb+ShNlLdKgW9rmEzvEfwkN7dca1yl129d+1ECtWnOkEYZjQK/q
hO7xF9PfxySorVAGPYsED0efPTadoQgT7LvpWEeNP8ZSlUS7kJNDZowhNVPBjxqsV6TqK1DbjYkO
m1A0WvfeooAPwOewAChmFViQRzdpDBi0AGBZHejK7xDhXPMtekD0Jg2HZaXs6NM3n911KGobjgT/
KHlVl5MJbChlW/gh06t8EprURiJThgzEoDXayAsyMrC4UTOJWTKh+LdFQU8CJOphtQxv0MpQrChH
uzpIYlxAR7cInWCI2uXK1ebLq9yHKMJBgI7DK2RDN8pnXRnOnvYFsN3zMgVUfzwt8UH8hGTHSQOG
scjI5Ght7nPA6kFC4V9/5CKN7xhKZ/dYD5mBOuZZrQBm/+8DVFhWYHeF7N0SgcAJ6SkoPUx4dqG4
hivx6nm66fGuCoKj4mO6T/ynRKREfg3hWr2A+T03fiMeGvU3ar3QA/U3dCt1J8ozJc0JCA4yY0Vg
V7V/W/IyR1dAmuVM0zd6h17ps7sakvcA/HCxxc+pIj7WUz+dU6R6YHWRltnlkp+C3OiSywgXNt0z
ky+DNORRNkH+Tl70X5wHItLzJOlyjJP08c+sAfQnsCTTcWGoRBBC8muwQqjxxNYb9BYKvlBPhwsx
Z9qWSAShVMr73soh33MaEwypZEz5GIKmBYeTue1lS+ex6/H/tCHH0lrxqzQgZhwXQDpcY7ebe1XB
Q4dBgcgrzjZR5CKDCc/itL0lTQ8i04mCX9VYuyJ4Hy4MMOGq2+hgwg88hz3qG24+OXirOkFl6hHr
aBB2JVuCkwrrCZso5cdYr74q1xnArBGG2xp7A2q95h64PlKfLyPSAJ5q0ZBdIbQIVqK4irBVjmpb
KhUv5FBzm+FMKH0OLKuehpr4t1QpcgqEyCLNuCGY5Fj0Rd9f7rvr/vTMJhEJyz/LbDCAiBURWJ7g
E3loYcOhP0UxCvVgR8nHyvjKW131T3/h5IQaFQDVXid4jaeukiKh9Qv7uARmb2ykhb+oFlWLx+3/
/lsAdLv1KzCn33l2d7DFGOCVOtl1gbvRiBq2qU6HSSBhXIEdlFxGRUGfitekJI77rJoLi2CVRNsr
lGyuPylV6NLfOFVNng5a7Ovm3UQd81u7HeDsljDQGw1RatVzwCUjIJzMVLVXoEr/ZcjMNJ4XChF5
316+VAJIz+0udqE/WpndX37E9uglj1YF2FPk9GpLbdXYmnSF1Tbv8f9ArBDFBxysI3o7GwzvBB20
/NmvjAsrIlIKg66QpZzg3f1l+V8NmIYT3EOnOz8PBhR2/PkqvaVUBOAuGP1UEhyF3keMtMqXPikE
02dSQndBocHz0rzveGsfERrla6Sue39EZHtMZ0f+z1BD/d6Akn/byzErUC+vgn7xKq6KZBv213AE
qChE0gyVYoG82NoTc3bynrGOeNnUStW+LvDPkEPHilCmLnls7Yq1Ga5vCJ1YKAH0UAJrvkAKsLjk
R3aiIbX/Pd02CDP3FZ8vzqrBR+f3qk5fBH8phdP7/mdWugMkZVBZX8ORPMW91c2TRqxjm1NfEZu4
eCIvNqSRyIG7L9J080eKQtSJsAbQX5Tem2vQXX0mCGsBmJToOVo8kQ9OlRZq4PFmjWitVpYxO/A6
NaImhEbxls1iXbu5EEESZrSKPhdwGbgGJoxTzhtK1HL5mYjQ+hnUnP/kTX2d9TZCIJqgwOqKsyBj
C8j3LqOWzHcyfgO5lnqIZJ+JcMYZdBm7UYO+uL4Sz+ZkGsbgpz7MM2MoPtoLRzzyWNqISP9pl6xT
MnMHRBisJRnF3hfyxQp9pStRR+W+cxpy8fceTE1JfM5BgPMShY+mpPZdMDmuxGDtiFCWQ1b1siuP
OHXCdVfWPyNnPQuZfSQpb8XVYeTHDCJJuIKYhFUqmW3K3KE3VXq+wPorjcCID9jcKQ6K2H9yY9tK
1j9adBCcq0pXB3IFuMQViZeF4/3D4rtwwOsy6gitX+o+5Zy+rwBiUOqY4civFypItvgO8n0e1qY5
UgZ9vMU8VUrP4lQ3gh+RDFhYrXKO0/z8yNiLyzt4If2sg4h0hdRJl/nZc4o4VQoT5U0cbVsXlxNS
tKtp7S1F7KdHwMOyzVok6H0u0NjXBmgv0cMpsruJ38EBoUUgDvO5cD3jFTtt0IgsHyFnBcLKUcoX
l3XaLYPqTzbXdSrhSUXCc6qYwn91m3CrMZkS0bdZdJprtRFAo2m0zfS/vY7mc2imNSGtaSkL5ivt
0blN5brvh+rj0JSSSC/itPaSkZWKFIMRBNP0zRZs02wAsCs+brI5d5BmFabG3a54NxdG87jNVPae
hgH9bHq9WLDRin3fLv1Oak+B4Sn/MqFsY8fpOPsyxMotbDFnsELIV2lD9PPBKghsOGK+KncLJhvN
agJypnuW49V/J5n4ZH0McL+qIUCbAdZNO/jH+DCSBbSlX1nTINV3ZbEO18RXqE+mqj3UzSCNQiTy
JL1KItzoJgzCyoyPlrS+Pp/n5Gjat/lGeA806TCFDUhzgNQyLDSWn2ekodHKgo0AnNzbTxnfZnvo
YOGNB6Dm5mtIAOK/dpQu8s/mck+taMs5sjqC2rvGLfptRxsFdm9dnm7p98qn49XtsN45JUcgHhyb
vIBfiG1HQF8X4Ro8J4/MqfiIiyQ2ncqecAPg1YV3xXtb0AWwcWIZODm3ARM5ouBsMHVNwEwEffzQ
xw7ijRvUvpqBuSP3ayNPrmbQ4/3MYEraWMBrYHZNZjGAOvK/pdfIX9yoQcSBnvCczDKYBay1AjjB
mTsfBsYCE1r52MzOtxs/EvE5JL3zGq8MhE3+84AVqp8A7Wks3Af0Kc1LFlvuJjMnYbpDxqePQF4m
RisRTRX4yrqjb6jjK1m69wEGBhAULoythDLeS9Rjshd6n8jRiBLiwuWLz1ElJpsjfPLn1IMidMp+
XsxhlRxqrDzGMjO8pqBzhBHs3VhDHOrsQA2UZq2vhnb/HljjAaXWgsGoABlS8fQw74sbvzc1uF0E
lBK0l5M6p1JMZ6cz/bZB+Rg3mJnY90M0IAk7tKgVm5KT3/8t3omh4c3ilgdRDPzJ55i2q6ZgQoKU
/R5zlYqyqRD2CQrgXEup04QOaCuYYrLnXs28Cqtu7kFqzyvcI+FoAe0n0MYifxXQxhwLPNigu3tn
mmdxvontEQllLISmrkN+/fTNrhAMS2CchdCNW2ktbRbpDci3QDEqX5DTJev5qXj00n71Zl8RELRS
J9X5nBkm4oFXaEfCmRBdMKkE3BxY83pFQT8mCBdwVV8y0EughH9ayzXhtJ7RTdTWJ+STWU+9cGqT
wHgVvc2F9FDT80EJxsbqqOuO5ggB0BrNIapBk70dS9elnp8rKEVs9/kYar/CxLTjEVkAelBtrDa4
mVEGn74pnkraQD43S1dFz6gjScSS5wnRaonA/iE8mfCJk0AM86Wn6Lse/5Vdnx4dZ4g3RA2asiqs
53MZWmt44IShZUxy1CiGqQ2IVl/fP/5LAd5xXFeov0A/Y5p7jZoJmfFquXC+DB/ClmzK1v2d8fAa
k9cw8muMaKMOlsD1Uhmng72vPB/kG/zR4PatqCTyYYQzGgho6GApswbGUo0TnKpkntPcSB3EUeWs
uuBicbRBR3L7fng96jYMRf5cXjV2+peChx0UgFwQFabR3yHUjpJtX0rjSjVU4YZx+g2p5sjEludw
0oXHhSHX9PE47luvPOoB5i2GGrkzAMDPHMwvTj4pv/Sx02gXSL9mKo0YnSzyGa+t/JFhV9Z26w+z
jHrNXTTxo0btvpYtt68wjy+trYP6Sh4aBX59cRm10OzRE7Gh1zX8B11ZrTfoIzUZifWnVrMeOQZa
yoT5Lwo2F7lNtE20hsAGpSpBeCIU2Tg1Eqr1kHfx3iYnt5DnxU6nWwmC2sBlhzVJ0epCjNo9z860
ZXX7klqVdl2Za/NDzzrl7+wKRVAPpt2bssGsdmx6qmgAzv86tk4747BTWb36GpvGK488YEX0vnPy
EG2QCKhSVyHfdPL7kiP0jqfNPdPLonUSz4801hBOfs56uy6hQMMxiH5npRk2+nVRp8HU1FpF9mdC
5Gt1tqusRmMIAp7JxRIrVuFlxsMRke+rZka/jHOeW68I0WZkgtrEpLCQONR8q8Rf8kW5CLsyN/g/
i7sj/LZKVG8aEWQmNfR7aTxb/zP8EYqYcd+P/91L/GRwfgSE5POeuYJ+smS8wwWdsR4vtn+a9hR+
apq9xZBrLrJyixjVVEbyoA+tA1eMsqi4kOrNhiRDL3SkLZ+bTMEAyFpjiKQUE8J7oakYYl1cHU7/
QaLlboMq4vROH4XGMlkJNAwSMeIsEHzVGGIqK2b8TCK+Lqy7k8I0B1ZJDzdAYmG+P8B57hxoaShF
tfU9VKhwF7Sewk527Lr4VcIIXYGDqVe0PlZfQVS8WDTM2WVZYSS9mH5H1aQ/RBY0MoitmZivrnCo
8CFFXd4wzJUj26M3WiBwOsh5fwq8t2HNwgKToxSwHJtJJJh/8FQvPQrdWp+ODU7L+vGcghobVX4H
9DncQBm2h5tRovyR3vdz6xbpz4QvrKcvLXNsVDoWBfRI4h02liHfp6WuS55JTflP6v7lRfPaHnjl
72TLyEhZjxxo0hISg2qTrwp/dBLOGgWITVLlF5Y9KfZsZkuPPEzZGjlYC75uWenOIvFipF1bEyTd
ZkZBu9xzzYEnOT3zi7d0q0YNoxJW+9PucEbQnriUe1SLypgE6r0+Q6l08dQPirla7joPDQJAafky
7oemF1qW6h+em1FKXk1ywpRllBlNn9Xb+ze54Rj1hYPClZCmmbeR/7PWKQFPgH2cRvXBdyvrgyMj
Vfp19BCYXdF3bvB5cflFQIZY8IxXv3druKJL+dm/MINpNHW3zJqoI6U5ArAHMrwvRIOSUZaadv+o
VKf09xks78+JOzAe3YzD4TSsA+igM/eFfwAWQElrObb+GAfbLoRt1Ti4H6UZxhGfaP6Z6Dvcz1fZ
AEH0bjGkUczhQEZSyxcdbYww8wK2ZKK6XhQQ1MmCCvBKN3t2DzBvRjalX4qMwODCUFH7JBIaThwR
1IlWw299Md2T00c862w4+saydWFj6k5iMH9rb1tRUSfK3d7XD6UjovgxY4oofsrIpl/XcNNiMsB6
aeau0Ce/pO35rsaJdWl4WJ25KAnrE1AeOQRjZ1xS0BAJIEmQRiMQna/PwVVsplhL17pBI+yb5Zg7
2zJW6toAFO1mbDElXrk6dN9ge0S7wX+tSY2jN4xll3h7zAbapm3OnMzOPHSJXFT/1DuCld/Cs6ox
ke3fncVzUywAB1jtFbQJIs/pxvZjloinRNX/3N4eqbo0LUyvkGLD4YjdyxkZxy3kykRGEI9eOCh/
ZVSEw2Pf6IrlX/3m933IloSvYUWdrV/X9W2uKNnqSLzETH/PeHuMlu22z42cVWcoqNpViJltB1vF
44/mE85LJBzN78okO5a7ysV34gv8mH4mKaTWYZnbxJ6JQbnl3EMEqpJ9Cp1cMp/d4P3yxMnrtuaY
hiBErSQkUkh6ZjAumKeiTkmcW1ZJSuXvAkTXJKa1v3lj3DtQoqGzPw0b5JzzgCZaQODuYGpvMbss
yCKjHbL8Gc+UENIGd1qopPiFJlmbjdclpSVXR7ncMKrZg+jovkGcJMNxMpOZDEaisvJuaJVX8dz0
DNW0cvokoPt+3vd+wX+oqsqP6IQbUXvlOYtcSdT5Q0EixSTNvwoz9WksFkermUCm1vFxeasy1NaW
Gy4SzCwyZgYQqmu9DeDPvYYnLAI1v46fq/3FP6RbWed4+kARV3M6PWFkzD9baeH7V9pR/zGIyYeN
O+x4np2AEK2dAtfrN802xDQ0Eb1Al04WQGqCjarBSZGQf51LZvibjPR4yWPrcKWlqmsaYK+ULYPC
PtSwy3vQlfaKfkTeDrLujJ9AaerFnGZ6BS5WT7PRxQ2ym856YAZ/2GrH5gsHrNCuD7Oqm0ABhNx6
dIH8vpIbcnGCaCpw/4gTtJCkoHdk67MzZpTBsrvco2uyiuHPZGeiB7Q+d7h11esYer6qxilzuJf5
Lz6TuIwe5wszRzURXlizC/OLUKRSad7MUxeCvccC5mXuc1tfpROMZdhUM8oOFP6N3rpHoEOFsSDr
DiKRvxUk4Syyzg2STcJz/vFTxkbuXeQSwqWz1X6jjp8giuG3VcPESEdQqkhpb8YDnVVhy2PPM/P4
5gzCEnbWoFiRpsztFyW93xKoPu9QV1qb9qYMRIZ/2pGTaGzelPxBtVqJyiDEaI3zWd0+o+opGNjX
1AzLDHyMa0Wuu9Clr+TNSRtbRbKV7Eb64Lx5UpoeUXV7GIPRBQHSbcwo6nGE6+fwxkog995Mrypv
rRIK0Z7fx5gO8jeNaDKGRcx+CXDa41OUSn0HIUt+8YVnEbHki9zJZivP9e6e3CEGzL4D5kuVlkjI
MH8sDLda4TkiqE6xwogFXKyALtPvn2QzKJs9G5jSe0wCpkl0ydZGhXJ1NQ/Mmuh5bFCyLeKhpdFt
OsazZl/ezrPa2frQITdE5oCBHDUWvkphO+uw/a+RVRSeXELsS67RX5tgapoSK3N0DqC0Hy4d3/Hk
3yh2lPFowLe1WQ3F06yMtF/gSvZRbLHmt2PC+qNyiKC64uprFu9BDg8AXq7GJa9CBreEXcxGTUSo
ET09DOFoakydYmxT/ixqr+uFioOr1QCXtYV+Lgz8XaXm8sbQ1oHvtCC0g6Od0X69c/0lL7SZt7ht
CEP6YIfw049JXMrwA4/WYJsZok6hQuKr2xjEbrdzN5PROOd5DxKSjQSVuQiN4x1ylZtV/PEGuGjA
uA3osl9v94n18BQIZS2+rrWRNetf/HXlpWhETwxYrSaVDuTG1clv58r5ooujmyv0ZleYolFz42mo
Jv9D5Kk8x4wDqOlysyphFdPzw2tpn42F0sLX+WumaKDezMNDN5RZB56KP/k7I6oKtZzSrYU6TQFn
gUeBb7EqDdtTWRyRs0FC8nr/YTCz39jr2bIg5l0UPG15vRp1ZIOgYgDwqHKa9G4CHJ+vS0xkjRh6
E5NtjeUIoDYbheoiy0pCGocSnhfFquqmlw63T5zRm7zlq8DVQ9L3I1osb72Pwf2czsfsZiLrxQRe
jGe1gIoZVy5iPssMfSmklehGVQR8duIfzLZN1eRO/M93ZmR2qp3bKUSG2vFikiQLzFabi1ldUy4A
W7xgY1DUua4boz233I+8LztzrPRUkko3U0BhVEuutFUq7nbuqyNaMrhPeKA52SlNCfJ168wFgQ7Y
o/hUoHkyFVRc5FzTFIXTe+GG0bC6MdrJ9qTiT6Yi7euO32O4KBEeZhBzhr6bIAtv+fhwPH+20yQs
7IlLQJfD8z8LIiZ8llCNuZAfvUpjdsM5vE6/fGiLI573d101+W+3zpWLe3vZ6qcYkXpAOnp8F0Bk
lGtJE6gKxANK3HFrexk+5DSovd5iSWWZBRtfzXqqCgppJmHGUpkufG15a0B+xhGqonIQBgFB8yDo
zq0M5lzLriLLlnl54i8tiF3HB1VXVLIjqhuB4l2OFI7c+kZfQuXw5fdU1vWBbbJOSEeJ9UdaaLSD
3rDxUl0gMrFVmDqnzAfN2Xbten5CITDsClQoFR2JVGlsWdHewZd4rKqvK4sC24y2ryQEf9ZEml+m
XKyc810NJVwAA5IfdI+rtQG+rIcP31pJVk8GJjbi2E083bo2w7PC/D1M8lK1pmFMyQBfWKOxUSqY
3xhehy4PpCVULEouXkYXzwaUb7S7/iXXDb0SMXyFq5uOdEMe/5eUdTGEh74bL6sqMPFPDgDz6TgQ
IUCCrIKKY0iLgSc+4jKwcE4p74z9kMo83WeiknM6rDE+i6Av2VshM0iQuwL7GN6PJVrJs4wgp5pj
UeQwGgUU5pU3dL/+Ut0JTKgc9susDhID7mG6CEGGHSWpLpVZ4ublE38bVnqjLLT9JlmpXynAdWVd
Um37D7jKvzUSur1YRPb2ZVJqjgTXACjFKxwRt1XDFD10mcJfe5W0gVX4ygUBjBSdMCvn20B2f1Lc
wCoYzWAjPItu11EXj88L/fbiHin2rL3CFdcyil1/hSkw89rIaVSRO5vD4gqsBgWeZJw/IVNozKB1
cP8oBHo4DZQuvrQxuOnf9F962l8A4/vmoEZaJSbLRe3tvHXkgSD8p3dXI4KN8YFTeOhRCF8aWDmU
04YZWFYb7rn6ihe+hZaKvQE1v/drJsB+sjcxYo+dOt/zBmaQ1mv3muqBW3CrbEyDdKdfx/D1G3sD
XwyH3PxMsXthneXM2yxvX5Me6d/u67iJkbADIIhRObxjUwe23/so4dMQLgvFoUtFuZR5B3sPDYPY
l13PGfH4x7Wjh4CY1py6KIdsELhCo3AVlvUY06/uwIBUQLlAovH74nc4zt8nsbvlKdDMUQCpkzmj
EDQkUP1TKxw4QPI0i8R4/LGbZvgtBDNG6mpZJo73aynelaiQ/HLxChwXZCxDuLUJyeLEpvM3uOpP
8ySiLmWvEu9hGbekkz8wY+UarrFCnf2ici1VugzVwCBGllSGs2m+/YqSxupLofHdpIRH48dK2ceW
yreBVwkc//MUe0lM8DNk3z11PGELhqKQLFj9Go/NjtM2JkUCP4CkHI00eOd9lxsVUIOPykCFZEgb
QJun/IfABMDNNIDM8Z+am4rRAtQ0/W2afN9k6wr5Ra0V7c4hTa6maBPysUI0rjedAQJN8mv7riSN
E+RWGiWoOHecjl3/xhxJcGioHs8YJnZ3dESEoAmq1ZpNZ8oe5d/A951X32+mOwLfk5YqFMrxVDBR
WK8mQY1IsEiIRWv/FHYAAaKPeX1pzaV0+931FGv0ZC4sEs33qDqoRoaRvTmd5OFz6RUTP56Ya01O
e9MvVbD1lyZ9R08LRllH2mwYibFd1w7wA50tUKBY0g+f3GZghLc+o6M/uXyPpuDz03ROk0iHpASi
7xGNCjyl1+ySO1/U8F0OQtmxdqCbxY03l9eO8ZTE+IBjaEYmpv0IZErmjMcpa8qtRk84ZEGM5zG6
fLpY4p4zb1x8/nEkAitCR9ysY52Q1kozdbI9FdYHbCokYBEYtRs5amgQF7INCOW2Bm3sPyFjfKnq
Q3lZNxHU3IvA/ffBuxWtYyXzWMmOon22WuNZjZWOZXA5VjgUG2rYY9slidrsPvsoXBUkK4AzfsYr
/ruYGeVdkuIwnKYA+ANaL0jSLN9eRYMWo/VlITaNVvS6dJySEUJ3B9tPO8Frf3px7ebFp8qlX9uU
hqeoO6PlEKmVrErciHjD0V0CeIpSMvCHNgvuWHwSaXDcJRq1QML64d/A2Q6fukL/BfOg0+vQs76g
iRDsYZXPTHAWXQxkN7Wp5wyQr40eNFpxBKLiOrelLXsakiNcNApMK7HbTLoYbUhOmYe0ERc3tYO0
h0fZxCLz3yx86Y9j/qZ1Nv4x5qDb0VC1DIsdD0AwIq/DJeuQvhKwb5RHn6TnpzEwbpxN0DG7eUOw
FkE3e2osVayYdCmdhlPf1wm6SQdhZwd7LPeEFTGht0FbT78dafoQ+JD8bqPnGakzbZQhD93Km7yO
DO/HqbQwG8S+ypCpbCobudj4HoF3NjaRzDewO6JdkTt18wHJmtyQ8HiIRbdNz4nhwxr9MkU6VHAg
HCZH5OJDpzcpqj7lSXO0Bbu33dE6Adfl4un8fRlE4vDl4lcN5HoGGajJhX2EpK4LlY8fRGoIKPBr
EcV5cZYt/jS61kHi9JqJFUJhHLUGF2CEr473qqR6nxb2cJeNOo/cmmqQFBVPt0cJ38iHlUwimsnj
PPmuiDoUvTkWWaXjEF2W7JEAhSFlTqHJUbqRpSM47vEKN3PUrFGNH7K/Q5dSoDTp16Pk5TrDZpTj
5SjZSn8BeFX8vMm6iMPH0iu3cy2Hb5Y8bE/ceuTcWsyq7QFlEeBbw0I91TmxCcw33TfhTDJrZLqW
VoNUoMTmKv/FOq4CNYQbW6D1bBwz6EOL9XObByvWcaaioTJ4zjVTV7vvSRWosJYiN32fP9zlkVQY
Q+QGemF3Jp30X+vOkcXE4hw+QEnkrPlYRM3bPoGzFFJGzKTO/aA12Zdzd8yQ+RC1NGy5wqDrwgPD
Ch6SzhHMRSwo8IOUDgAkT/4e5gHWimtMLBPpZbCgJsA13JhN3T83et+CD4pZbe2Vj7Qncx+OdEaA
II+R+7ABJcTnMm0AP6U5iW4nQ4Fy6ukN6yddBxqfuy1t58fzCCFx6dOXCp6ZWh+c0iewFGFgtTLX
tI8cCS8lx2UHgFLPZHty3G9h2oJ3X7jrw+HhB/t5xGgpqv3zYQ9KTQOQELgzphx7tCDLH0FrfD5s
Km870TgGRRCgim58YU93NJ2EtERVlVUN/1S1aeDDbX7aAP0C5+pW0qsCynrOYURs1nuW68o/Qf4X
vDs7H5so+sg5e1vsm2HcvHS2ZXeLmWCYi4d9uQvUY2TRl1+RTts0A4/lS9j1krH8UiqMvy+xCZHy
wjgBZZUwpFDGPu6vv5T4/3d+1QjjPGnyUQ2/xnmPDwC2sJPftX7blF6Bgdp7YccCI7wsWR1c5tzN
xLQOaGf9zkYFKODpLrDznpNWwzLuf+sLSQ5C6e8JeCtzoQnnkM8PJnAmxUMFIZZPdf55pAKRIrFg
p9rFVozSSgwSURsu8vIwlpXe7rSfDN1yCdkqWtwlIpq95Ner5hYbqYGyd7SgzNa5cQdSjO+jZekK
CCzV8O8+Vh7G2NnEY+Hkc41bndx+rgEbMi82pQx9nbL4gq6sLM22UcDs9voBpVuhrZ03SO0QRbwf
ezMPC4fv2OsQXAMCyYgs4EPMyVOg+95WaBQ37lTyKILO2jVWEXsUW8k5MnYa5oCzmrrJd9ZgmgkI
1Frj9VsDRf4TVprTe8aAeGMjeilASjZTFuYGftl8Qq3fa9hnZMjxN0wqqFzy5iBIg/6j7eJ1IEUJ
7DMHhcJUwxJQJZQnZf07o0ayujgQrtrjKd2D6cC+vplxtj6zk60XQkr9+wq4ZAKtYqEccawiZAbp
aVVdp+Sl6YF+p5qD53kFndXMAMusp0xOUJUfVqcHm59ANYChkQDSXQJcMcoXUjz0MUIQYXnW8vAc
oU+KbvSpXuNdt2onMZEGALkBNTY6rvzq8jwVA7BgODehs7GWrdVXGfWCenjLy6G964w0Ye7eBbVg
T5a1nRphGYUIklfk5bvJ1nG2W6XGlNtjvroHcC3rL+dGY2beWiF9PAZ6IXWRpxZqlh1J8brlu69Z
pAVgXODZEC+hgvSBhxt6+UGoNfr/gY6PxkVdhZCrIVMYR3TDoPia3gQM1qeF7KKPLdxb1OQtcO5f
nmCgtonF4d13MK4o5qJNoKvqNYknywx44fVs0gjyNzkekcIYTmyth76e+XLTEyHJcbLXuWH5C6LI
F/Pye8cyY7OECfTKFXr0VPlXG+tkdkvS0egawmwGGSSpF9hts4t/Bpu7PVVMZNh2DvQb8OZoUJNX
dvTldzYerek1tnn6pDI42ZQ6QGSZhQkLEp8Vd/oOE0YeKqzrFE6pIAhmGnHYnItCeL59n1I1BGI/
2iaa03QWjaJUDSW2FdAw/PvaA3MnDQBzBpgUXTLwn53V7V/kuEC2fY/dH/JDlz6wCdZMjrYw/azT
WB5ra3fHCFAsXiw5N1MY10hSTYGC+6U65cg5xNkFdQFwayZ8gzZMUsAnI0Kb3C7ovRkYlmavUxPZ
qEkcoUOXtBfiR675zD5HF1ljdZuZ4gDJEFmsrdilGtIqlV/v1n0RoKvFHd3awpkCiOSO5tTxAnLz
LxyxrTutig9ohmVOdmC/9DJghvvztecXIr6RDKICkDdy26gvx3FMItkvREGP09t4N8ZqABFP5fhd
PWwcAPlGZq8iNCrUBRBK0jG+GcPzXW3A+yShtrMGOR+FjcoM09/hRoA8h1V4HZvLUqdbwuFXep3P
vMrw4ZQulqwLlZgajnM/OIDy/ASTKn2buEe4Mym6TDZi7JUhAyjmMh2RF3/OmZiB3oOvzjsvOzeJ
S2HYuMIAyKN0YQHRuscbl6cNsxfCiDmsR/i9juWNE0/YYhAbfXHyc9BtT5XxrTyUtt99EOx7r0TU
1N1F7JXkYJjdkob2d+GW7H4xASCzfrv4TMTpuDvsrdr2Qltsqmne1mPCXxbRoDtYksRtEIEWDCFT
uko/BCdmHEMCnI2BXBjYcoYKVcxxq6alRIJnzuRkwKqT9FVDnfQxdnPUfKcijOpkckeRNSvL+AAS
wwQ8vPa4X4deFDAESbfTkWNi2QvlnEmzB0AVahdRpWggcJDCZNjbHThSxDvoOLToOgHsnisbFlMt
Qs/M4RzfmSdjhBm0bPmC4jY/kwmF9bOuptxrKsHm43ah8UcPgEQ1sJYhmMkmYDNM2praw+fHP9Hq
Hdx/BBiTuoTr0tYDPRcSQbyXEjH+E2bfQMsXIfEIFSNoSCJaYe1Dnh/GM/dL8pT9kG0YLMmYZfxx
d6/fJWYJc0cEOUIrXFeEKy1bLPn+csjGhQdcIuPDuLOypgHMKCnJJA3I16tN3TEQ0lEAxJMbuftw
fR7uUpfCv73XSdeBvSR0mG7goF7ugfbFfd5u/M4+DZxXqMvastXHPaZlGFF8DGEJsJD692r5QkDz
BhA2eoowm7xfFcW9CM+gGI3U3bGJc1l+owm2hYV/7oBINccYvt2nZSY7izTtZd/Yuv0p/S0HVnoS
JEyZeRgOJ1uU3Io0zyAUWeNV3BVNr5cTmionM5wsqVhZNGkRV0cOrVmXddywL2r4kC9kdA++V5yD
+VSv1ZX/lxsaDOQrstY06Ae941Frzim/2jubFjNUUG/+lvp5IIya6GZ8WsH7fxNuSDYpgkkzTDkr
H2PNaBDztDdgivYWr/LPZMfevob8XcHofGjnJa5n2Pw+ATfU6wO7N0kqzDlc0XnT5IBYN1nxhIy5
8eOz+HBlNQ0YH83g1h25GEWNQOQGx8dknit1y4aNBkw+hV8/WEai/XVILTkzLhEFqy2chDYvR73T
xZ7ieSLlEiMzGAd08pkFNKEmcsKqgR7cL6QPg0Ll0dIZndZh4vGdTX7aLB1Mt5xEK6jl4XyTqX/c
bg+k0xYsjNZTEeTM+tbGB3jIibUaTmJOJmIiUAIaIF8LmSo+yGQWCWCJIKHnvyLN3erpwfV+BPtP
h+PzOt406n27WR96A/BCuJsqFfkhnU1z1sN08uaILajI9HwtYPvl7/PC3bvC0GBVxi87ScgASDVy
aC9cRcIHeTG2zBS+O3ay0eTd2Kzwesv4SaDbsZur+4qFF5SZl70KZUPpUAhsK9aYEul36FJeYVAD
SsKUpSwHSNfqyRQRDSa68AR1sWayxPwvHL7/qCX95WSj2oG2sR2SJTF7JZIgEmRbkYnwKv95bRVu
1I7Jv7sBP8QY8XW/vbFGRI1sjyt1BKefhQINLsPtWepuWMikn3eJcdXOeXl/12S3iGOGAnt0isaL
rGkg9G5h0J+eiSF/bapbZqcFEGj9dVsUHa7y3YzIhQ8m+mcAmefPWsox2muneFq/WFD8dKlOsYf9
QEhouAFaiyqorvp7Z+xOrUqroucn8bK5YRhL8V49lO0zMiLDh4XARS+4PKW+vCG3S9oYAfjtQK12
OeJajCR/6skVwvWYeGv0fQ7rn1R+knPCeBDPJkOhqQxHXpYZFu8Ew7n5hV0lbzV2PrjHWDQhUl/U
onKZArzj1umyJvmTX3Dei66mOlSlTvzt4r85JUS7FItMlgQd+a7Gp9VVbyr6WnDEY5LB8G22kgvw
qTUhj4RMbdPXJZQlfnHu34uIZHqY8dOO+XUjch4lPJZy3qmtWTNd26CITAG7XBZ3cJngMtwCTumm
4DAwLNSZDejhvgNZBE5+8pBirVy552ppzGht43LTRKMoko/kCvjLPXOfrIqtRue9qK1bW++F7cWr
yY+ds9jeYJZw2jFlT6jBthM24j1yvpwVTPAx3ig4rb/2jHJStzjg7DaiSRuhg+ZGg8Q2FzKR9FJn
URGMibox2iITHTcwUvpcd5yHVcrBSfN9OHn0PYWFQ2PkO2k0B/WZ/gor64QrxBncjqLYZkyugaWI
BRPkTwyyg+aILezrfkwPSzmOu1iPfXkz09w89uKkL42CAiqb0bX6JZm+KnTIHm3HjUsIBA1t7a21
vhd/tihI06+EYgHgaVsDXridbhpNpKcgC9S3X6zTDFge2nqnyQeBqzueVbi41Z4iDyWfzOZt7tUq
ij0TnBiKtA+4ROfJgPbGYjm4W4R8Y69vORQDvoUnXphaTfwNnVo3ehDnMjRy57WOUbUM8yj2Ofqt
H6ISRLg9Mg3bpsmrZJAyotWFWJAExNt2ujFrMV0CQ9pDknCDxjdkTGezc1N3W75gh1BAiXDu42rT
suVYadI5ONi6J6AjHsSj3Nu2dYpfWLo/WAjMPTieK+cRTmr2Lh/mMfSBoGT9dHYeHh7KrK5KXcTE
O/fltHOkDptksR4sooo6vl1iA0Wu3qa7gXZdZ30z6m6D88XclAbiU+Mg3DGAhPrtS+sd9HpkTSif
fqFYbivfVZW3FbHly/0YfyhCbxKzuOnu8T5xdoe06w5dotJUf4+MaUTpLY9/mQ/QxvCIVLCme/hJ
KPZHxXAQbySEqFUYLa7/yf7yjNduV1nOj5OOR8knDJWgHqltcrTrUtWx0XldDmakBplYK0dWJyCv
YE06c0WWPEnGCKeSskTOqqGms9FciW2BHRJ6PaFJWI88Nr+4rjvzpuCq5P80T7reKH6FBCXJIKPe
xIC2jdQlXkSRM9BPiZHJB0INyEmcVqNziojvpEbRSH4UJxKR0qby1oEPOCIzgJkja9WRllsvOLLA
WnOsjezILJfDnsG87mPdR4qjIM9T0fp9/KQixPAHbIwXUrawHBdnAHceqwuQaaXsEOmfnISwmevW
UEVxZEbaIY+Crk2FGXaQBMxiUVQVYpmJO+xfBiEGZuRsRS3v5m9rq9JWXr4VAGP47HIS4PNS/eCt
Zur/gQNl08OkgHdNf39+1C0UtBuIZabPLlJf9qZCcrNYJGeDUq5sTvxUd6MrjNJke8t7XCgCLUlt
/G9DVxUIur5tGFlH+CKziGzqkf32/WgGQNKK8zg2dVrf8VR3FEh0UCyCZZbJZLrVqH7uAwugsWKa
AsNoqgbypsdDpHR+BfiX+jCQZRfHHfFlhmoD551mLUnWi0WxMDi12E1ngThReYFiPrZgzIZAb2xg
rSFkgUQMKoC6NHwIqp680dI59Sb1gQ4wu3v/XHtf++UArplA0hZfOFOlUJ99sBMWx1R8KEucbelz
jgUrmokSEc3Tc56Ih8cGijJbPipguB3ImGdwazGWMYJhWJuHUnUqGZ9hHzO+9lEZp9P172wcBGns
VD2WoOncL10YtyBYqGOreJnsnffR2FDc7Lx0BqGbqBe+EpKm7PxQTljmXPgw1E05rj9az0XmCZQX
VXo+xrbhaV1d0SxmmLRfIn0KCg3NPF6d5r1N9Tiiff3cdsDsNPA9soccUo7/7Z5JbxvbPQtc6+vI
InkS8dw21BxsxLU/jnprfieceptMBMrV9LED7HNBBkbFd3Ou3s5JFmFA2slCT6rXFOiAVzjMQ4QF
BV1MCeO37qcDHhhRNwQG/Rbk2g5hkuLirMhnZBLbjQGx9wuWBM42vJkv0zMN3wgoFDEEy4NO72Wd
E34jo/lC8psvL7K3VTgvbeUspbqjHUekiLdP4UrmaUCU5gkqklHGdJla2EF315+8xlVaujPlF2AJ
BcBOf6RGQlYVqqzeEyWyZPCtfcw7EiW5HnxUMBeiqupyM1225RmlWF10g48b3/hJs1FQtpEqtCTY
XWoSF1i++Vqpz4Ebfbc5WH+JM/KgkXr3lCnbmaM+oH4Md4Ga3WNGafidizrBvkpEwcMcPIS12Dfi
C1mJJx82u4Rm/vzSAKm+5PB34PKh1ZWG2nr3oo0+EMVd1VNZR3TLu0GzOnt1fCMzzf15evJdxxvj
eMt6dmTUxUG+hcY19/p8vYudq/D3ZTvw2ky/toF3m0ZS2olXZutXeE+Yb9Br1E0+TVZsrRb7Hk3b
z3G6y699xoiO27isTwhWguH+S396VzVN/91F5hjRxKFoU6TtjPExc5QPv77vxCXkA8TGSEIJntP/
IvWPZ3hDFq4TBbOu/If2qivnAZKCrEArUZkhuUNdwVCaTQcHqxqxjKbboXB9dOZxRWUppRVE2Mz7
oKx1Zo8ObqHJrN9D/dkJOOso2R2vevrwiEOAcA91/x3bNB9G9P+UmLsetzO2ckFf46st3Y7PasIW
cVpV9jK3Hv4jKeI3NwHv6/Cd/mFVlPvKxCcz33OX/r2SP0NqYmNtgvlRyNzJLU8SlIBYvNrpqqz4
2dcJr3bRjoj/TcDTb3m6xdfELqnDGeuvoTQnPaJKWzX7/zHc7Y8IcimBnLVh+9WU+dUMEHKxESNc
DPuGpH+rKybmUghhEW1qjyjWxj+h9LCWAxubdo7PtuIpvUIy+IFUxozm04tpqMr57K46mixjmfV6
gyCBhlAlKk1oVpf1DTML+nqNv0yBnnZW9L40a1Ql0lEaynryGk3YwpxVojNm4/crZwKNXpjWoyFS
zv69zRg/bv4yFr9SUw9f5aDilcrlQdXZwGE160DslMUxy8NMzLI2nIf0odrALv57/jmP3gJriPdT
fptR2aA6ZOSZlm4kXNLX45Lh9bdCN13CzqZQHfU1ppnwNF4kZtObr58Dpjt56O+YYBjv1+oghAhn
RzDQP7qSM6kAjtSYuDp4NfU2lMCxnRzi+OHD5bDLuZh5pKINRk3PpgFSiK60lv6/OeGS9iAhjNmO
B43kR2TjUgmtzAVv1olJxwG9+L7t4x4ys72dAKLuLwPH88vVyMOTtMlremiLSz9aTr1UeZ1l7LYS
t7cKH78rGXHkTQYNoI+LLPtnq0bmFee9rm6Q4+cBEE9rsj+uUAC0Bmpy801u6FoFGog2FhLTpPJs
UVELiBUs4OncfAmCwkvpe+nxLsVP5zUyCJj22/MDKMsim1u5tskjoBOL2I8W6f5CTkCp28D/x6jP
6YgDwFf3/yUQw6oS16kntQo5kObHCHeki5ZOoepNqpeI4+56fJ29xBAPk4i+EKtgTUVdvY/gSMCu
W7laXonUoOLlk7peyomMKmFjfSFm3KZ3sGwlEz3FIosWUiGGWUlb0gRg+nwAApZLjEVaCi8l0t8K
Lh4lTNWhZiMRr/GymczNL5NtqgpmyL650apYOGSUjbYuicMkIH8MWIatiddR+NUUYt30c3jhzU2E
LYHFoNhneHrYh/y/jeTOYPQk93B/WUjBVVbzISzakx/7Mk5Ko1G9nUgHinLt6mYOLrjBq3ePARkl
9k/2rJe9g1tAPE08SMxcKhto4LQ3njWc31KAdkqUxqUcqRLdh/1H6DCCzMAvOtPeWngKhOq7lsDG
N3ik70UYPGLxS2dIEjV8s5WoAil0L0qIuLG8zplQIN2qccJli03lPFhXpnL0+lgCbjTf5yt0gm+5
5EZlN6uJ1D87ESc0TLIECZX8GFXQFAhZwONmE4NZWD4nodKGAvPom7ZqUaO9uO6ljEiP+8rYb5qN
nq3j/wnyv+EhZWNnEXT8dy862fs8eEFHAmd6KbOpKyXxiMCdy6HA/7XouO6CqSeplXtEf/PetM5w
XUGlUsxXNH44A68SLjQN5mAJ0SEL1xBcrf+pAhEfb4UzxtkfaRahySKLrHm0ZxGvbx/oA5gUH6vT
kLJznKnIhQl4uyzraY4271+ct9HN9tTveOaSGMihKzJGJJ6ac2Tr1gkcdZEGzZisXit331Exj2z0
zJ5REfoyLa2aHdZc1zX9m6iQV1c/stp4Aq8SwRTJ4XP5UAki5LNMnSx17fYwz+ia/qhOsiXRRYQE
nl18m5J13qNpgr5cM15tEcijUvkX7mzLFDZlDzJWyBlydlhnDvv6xWvTXSO6dFicLwjual0yqkPz
Y8+nGpztb7mNrkSBZ+5ER2uBS4Hnj8WwuGN2dmtdlzDzp0ROYJKkj1sfsWSibUNYhSTUWw8xpHrG
ATMqVDhuR/RDqu17qtLNMp1hnuCZDW9ozGpEVQE+9cQfLHIDw/hoySbrxXzYxIqtvpNbX+nkMYob
t3uKclnj9Ok7i7Z2wfmrDnHPDpAgEIA71CT32vWHYTGOz+Ob1PDOdIcuZNB0UUef8xDkRwhpmvzE
YtO/YEWyDCPPckTMQuUWVvpzLopCuHmHJ0fYh5EIfpN3vZwF4Lc7G4ddXvL8L3ElnQFV1KnfdTQP
93bDSCIQAZvp7CugNBU2qqxLJIzQLO53TYM7pfLy99Q8HCF42PWTZVY8XA7D8KwbgDyyO+c3l6k+
GEJQxX8UcEvXW4NxK9dA4qityqM1Oun/gN0KcFtFWqt/EbW/ixH9B68H/RIbnIH15ahdYzpMdeES
JFaKGW3Tlal4ifbO6XBQhlitpKA9HgDFjr5h+8QOu5E29iE06nXPU6+untuJxUlSaR6D5HZuhe++
ZYl+n+iFARgvogxD75PndIYY/GtsULZl6ncMK9wf5lBQW93gqkzdJYnYEa6Eayj1xljd4OaWBRSe
UpbIpQl2RASUaFgtMMucb5zbzxa3K+wtlpeVlLM53V1CJqDPqxhVBMjEzNZq+X3jxO+N7cSP96rs
fe3ulRDyNrxufo2wC/nsFveV0KYDjadU2u7/vKMWiaiBkucpRLiEu2erc7ghJ8sqzcTL3FAGmFaT
US0GJ+Yoe0ss3beAGHN5EamrBJL0yA0L8QOLorA161QHaaNgExUPwGS6drRsHYfHXDVo2mdXtZAN
aEPDOs/ML+9EbWRa5xYQblf3ECXduSW8UjEUZF2FNCwMbrCUgVyYb0RbO8IaqSplTCuhGZYygBbt
8/EI0WxqcXtWW5ocmLvGQR/Zhi5n3TYCoIy1y7TOoDGHGoIR++akG2WVPMrEjm0PHbVWkimVb5gD
fMzZePYquEuVXyIUO1uUL0iAHL04DQ9B9gdnqDGlv2Khj7P+VrTycimRZWspheMW0Xlu8dVXai41
NnQ83sMlWJwxhFEFLxFqfh4twcw9zIIulPSxNJtoF45naTs2cKUppEQtTmVvOMv99QvtaQPWsw2Y
ST1C6Sd7XjljpOJP8y/Y7jMrhziSBXwe65L2OCQ8fDKoXrOk2MHa5EYm8c/lNenTucEFdqvzDMnI
8zffAKqmbESB1RMBXzprztNI3TCWichI3h+fjo//DV5efdcsMyef/0jhdjbFeKatQdWwFZmzJL1I
ytRuBmj1psThh6fqFTloXJAuXBFWPAtkh9auxd+HgmtngwKkYnobev2wFBIPQVbh8oscP7+iZ/ct
lSlurcuC2IqB9FRt1t7WbuyAfxlsauudi1wwGdfuj0XhhPDa9Dl0diIbhoAvZVv6W5OnRn0/sCyI
HG6xviZQKLCguaMFJYHR4iQPVALxKLLwIlOgJCixP7yl4TAS572NRm38wuF4dTVrUJUdAGdrjO7H
Gh69q+uF4sHxdvPlmqSzehRZNzGhlh/bsgAAR6+NLv9IXo1OM23ijljxRYP2KKG93ZDum1VyS61r
m8trHwIpaIUdyPxsqjy2lDtbAq2M8JTbGWcR/RpUrttiZYxKSoqJvByVD1Y6U81nVMJnWPPj7OKL
ZaFDDMUkg0aQcq/Y09Feeiqrs7cu4gV0pGdJmDbIcPf65gk76PYjpf/oZYiMA+7b3KNo5e//WCKv
b0S1Fo9WEesXuHmPJ1qG1P5x5bQgN9qnn+esrvutaqEVvKXRFksbVSte5RRMFZH3HHKUIHhjiESN
TfgHgckvkg59tlHmhJIPdjRnTVw+bBxU8TH1+WW186nKHZNem/PnRh23YDA55uJZfQMHcoJfZ/oq
/E8VSgc3BmcDlwammoZ1dtv34jhidxzDmgiPpj2NWOGL7RLUHjLYQWfOPDtoRewKTxOKkJxfKWNj
zqwimneirXaN73jAPEomQTPZ8BFStWmGZ/AwsFDuMi55bgMzE+VVV5Ah/dhQJH8dlZGT1ZWLG/8I
G1URxqlYXqDIr7CSoW+8qVw2NXoncJ+qI7+AVTJVhOqfc7LKvWsUSmuWvynB7nyzbyRC+lldN8k7
HPFy00DXjDcJmompN4I/BfQL/L407XBQW1oJqTJYCAdQ5edFE9QBFXs8itIZrC5KdC8c9jjUYXnc
Qd1O19r8RxD/8YGI5sbnCb1aHFZgHVlrhA04ih+mdj4gDPil0HA3b0e2uguPeCaN/h7nFudfel4w
U2YFJHiVfVvyVab6ZNssCLMAoaHe53C/w5gVEiFw/ukLJ/ZqggZTcuzqqWVaS/T6diG9aTajukyk
6r/7thxj2Ky11ivttgnoTxwN6/nnFyjfwbJaaJdgVRZAegVSGbnRzHhjjkU7E3XncecMamJmPXZ4
BEb1vSsLPNDhTaumRfkf0LCBXh6fr1Y5VDsUoItrNjPXW2zsXbzPw2LhhQdUQPcsXrnhT60Zvd2K
54OeX+urdpyhURLs2PWRqfrcdbhG2iPii6UtJVZu1xv9PZhMi7jeC5J/eykuWDxaesWyL5yQo1AF
qB/ZZ4sRIJsvRwXySnie5QD/ei6BjmG71V9qoWOUsm716/JxKh0JCA1bJDsMj5U/P/3owsM197Uo
0DQjs/hHbCCPPpB7zQtnKXY8681X75kseCqGYzBf4aB5lDcpT6M6Twgm5xUoY5X20VsoO0p/BC7U
BsCLQdjJ+At8aVQPoxB2S7y+iiqw+8xXprVOFUaNnkyktwEKnZ7hFV9eZmBY0RJvr1UcGHm6QKvH
7FwHZZwGUCjlKOIP8f4UIvpvVy2sZxT09EBEovGOq0HZZxM/4UoB2zF0l59+mmTPfbFmpKt7Vpnr
l7s4woHa20Ua3XWl3OW93c5Wq5miT9LuSmCSpEljdUUsO/Rd10rBohFzgEr+ZBAzzk18LVFuMqti
A6IUcJke7kjuhGCsDVbK9jEuTv28iVnHLRHvJBRRKAob0D7W7hDoLE0hu/yG1lIu+EmiwX/+YHZ9
ElO95S4biRo6jB5F1VpP0QGmNcF0UgKJN9NGupyN4/aMscB8C1KG5XbgXJ8YPZx2WS4zI3h/kL0S
DWcCTXywc436eo1KPz12v3KWNa7ZwfIc0F5zKRnZ3LE8Cd/G6FL1+I4/KUDkB5qMLWz9I16G8359
mSzsdchQruxu6tibtYYO9x40/T41wdDHx5yUMAf6BWnswRSdD0hdP7aRiTNcTq2/QfGtRUvbg7bx
bp3DoSttOZLgddKCQm6jLxvIgGg7CnbgtdNaFAruIN1xJvvAQ2a7wsEaA3kJ0scJcUFEn2osFPPg
1K2oJgOOPiPecexmhR6r+M+9eqrpG7IpIcCSiTbxdZSmxJnjin1ZsjfHP9KU6z6BT7P3kW4HUbdz
XwVU02uT8S1FHF3myJf2dO22puA7T4CAVl4a7uM1cXcnkj2VdE8HrW/LitnSJnPrPmf+YjZMW04k
u/vs+EC/74L0FrQelCYjs6wMiQzmcbxl8GOXDvrOYdjNPR5xzYdA15X8wgy3/ShAJ/2B3GvPX2i2
0HkjpnI+W9XsEFEg7zjE3+ownFNwDJMquqFU0mcSAGSb0eBWPj3StFDwPxol2VF8Hq9oxYBQxrAc
5JKTtYIiOYlDOE7+uZGd3gSujk7uQ4goPPy0eWQLdxYhTcBXNXOJ9fJ4RnNTvnBaAFUGWzKTNyNJ
K6EcTzCsoiGZWRJsd7eEVZj9K031yx9xWcNb1uCMep9nx2JpqSJI+dwDEs5rXmDxatYif9UYq4PP
BugolrSmbpXMieAovmBokE1c7visZWaDrvf2J07wG2FKZNNeF9dY+fpJsgOpoMdVkRfSFbs2+mUB
xqZJM27pM3y3wJVG4q00Hp4oTeI4Qf6M+aNNueSM2PV/slf+ALradio1J146rCax+bOFIIlks+UX
DVtFbzmE1YttbI9j+0bMUX5Ga26a8OH3dbr7UVBjf6jYAPHYzL5pDPTi891BPQApCNFfN+ls89rd
zUQD26u5ODF+thN3v/5/XpKXi0044av6ntnqVKHppiCdsPGtoKsMW1tv13uGdE81ZpaKOIMJrbeK
7gB/7EnxYGSmX9mHwgfGxL5PLG9EfhNQg7Dvsw3g/NTzQsepznR2kcwtMqDSeNGnakrjBoKcDXTn
mZUDE/HQfJdbwAVqSRyjvQoLGxAjn2hnG2LyTWsFm9mSsnFQ23CYQN9X8q+/lC6zkfC1hZuI2vsJ
uixH8a6t5M+djl/mEwFfd87aoV7sa2PR7l6kJfIpYhzsTG5RWGoEiqh2SsjOrQnMfhqdikAAXj70
vdCP+34n1+pPzcozbgEVFFpFdHe8n3bmCV4wPItQ39rfiMtZim2UczRFrdq8oAvblgMGhtb16TkR
sIAJzDCumtIruTcmtYMojbeSSPcUYbgWFJm4CPlllxx3K4CrqjaCBn7nPE+niKA4Djae5qAyCkqU
NSQLERoZFV3QJwOjH5LasNMleFXlHMe4FvEDkQ+NiFK4I73+FbUWoidxOADUlrkYtK0BO1oBLRkJ
bhpY9y0D7Gssmu3blik/HCUtj7AKOljx5DURXpritzn/BrqO1AWiKc3rByoZEim2IBqivMpUwF3R
6PUVXUvVYPz5tXefpUXn1Moza28JQ728zLNW0JfOThThJqdn9+xAiD7BtWPXVBh+Fn5HyW+kcLIh
5J+lXQ0LkREzd9JiWI8VxHoeHFFgpdPIbPiR+ybb3E0+M9EP1plcQbU2fLIzum+WqqIM2596QsZ5
yTgSEyWYQJj3wrEWgTrtYdLEBOCZje5zmpB7qlN8OPkz7D038pLLfKPm4e0GYA22M9avfT531801
5QpSGlZGCRJYxk46Qb5z1P0GqM4TYF8KqGUw+zwyU0XwsRirBRmI8hoyDtDgxl1dCu/UhQIwgPBo
KxiKkHj0UjnwrwWAxbqdsExyyQwMBONlF9b00lvw9zRp5YrrD2e/y1wVkUFDSV9sr8ugMsqobGkC
MRMzl0AAdEzezxVmQgIeW8oEKnldRQ6r4UAMIOaLBUq3gNMZJk0nGC7BtgamadTDT1shIsswt4fr
zyatN9tXBGeJdoKooAn0SlZFChG6/BmAKpaxxWQCrLeT07exTFwBySTeUbLspzZdLLR06qRT5PiX
rVXT/8Y/PyORnhgfuL8xmh8vG1tW067GCIHRR6eP0SdL7zMAKEBjD9LYkEbeCV8D4jzeueEYOglY
7M+V1OK+h7MUSR+96BoGoEatEiyAyAgNUuO0buza5kSBoaiZcg1FDAkAtkczkfXVDZKA11JI309Y
s0qojtOoNswMGKTH9y46HEtPPsLowv0Hdym7t6dIOkWbRndNFp1E7LEiE4t1vBKb2qfdUez3Nkl4
rIB0TrYj0hescSNldKeGdh/7PtgudOj+GOxbhr9EMCMvWl8mC341CWTvrUUvbnvjJMVLMfHa8In+
NgfQcVxWFYAtrNHLCBy+V6+XGr09pAhKs/z3o+CmUoQvw14vY6smUkvV5LiQH5KvOFObqdJtRwLj
TBKE5m+7fb3dNiz5Vcqk3NFQnEFzEe8ynbCG8VHFxbgKFAqfpS/2SUQCD0T+FjEv9KVO3MpScMmQ
1O2py41JWaxpBbTj3YwT3oAgdr6zT/66sWJeD+yq/6cbjGq5I85ZSN+nfi67LGrkeLueIBFyG4Yh
L7E8+44QUGL1J9on99Fz8lfMsX8Vx/9F94Xt11LevSgjO6PD3ZiqR87menp38QoGeEMgeC33gNhy
KMWWBT1cx/vFvjXG+gwylpv8quJ4jsT+C3HggT/rVhEC6m0T0lfShEwQ6rsGFkRlulXXZWxhXR2D
NFrPA2XrjUiJfETinC7ZT0UhaHmnZRbpPt7nSFYZdGzqI1FD9w8XP9R29DAaTYkcUanxq8A9edEj
T2d4OckiZUZpwiugR5hV2UrjcOuioTcWarVfahrlh50LbrR5p/XWQoYZVeaXzS+m6PEHt43AeK27
0pW2Hlh0CrZBL0xTYBvY6vFJX072kHFOx41R9K/hYEaLauZRt0XFOb7GxYLf+Ha9GroZQiGGkFTx
+5L1Cz+FR6qXuk0Q3n20TFu/5WBctgnngNDZXQEem8vBu8rF6dZ0ADWIsvh/00tcWa8BPhI+qRpN
Umlgu0wvwd8UFDY1mdWGsJlw15wMfWAd0rUykb4CjsiNOm4hhhm1npu1VnyXTkAXrDZLCj205PfP
E2/MSeA+WLZZEZ4Tj/yyV6aqCRi3GO0cz8/jf0bxIEEw8yAaSzpyTJHjqtldr81DG0lwgS2DGgQT
HI1lnAJpzNarcl0lkUxDtXELYpFH7oShhucyiVMex2WlUt/fLRLYscyeiqWHRGSRGVeLlA8hsn0N
lSO7CurBOzgFAKc+AHTwTUgyAeIa2o4k69xgUqxh6TNT1+siyY7snafF4eowed7LjEjFCZXguwur
Va2qoRRaxiGYHFDR9cuv0GbwyADzoTYnxRcuIkN8PRpjxhEEaeaQ93XNeuIvYKPLGN31HDZPVmC9
8LmGx5NA+9Itz+tbVGUwOU4WbPPPYkPfsWi+hO91nwxhypsOVwF0fhUjZiiIzNCySSUzswmHVziQ
ImSB76s5MaFl90OvkJexgM4nX/chEuD2ubRNrzRhUZo+qJBzpoX+u7Ng8XzDtBtslv8SkMTnJdzW
wuFtqX9e6V0BQmrl/vECEeVcFgh4w+M/e6XZw0bdcBkAy1a+NNJ4r4GVziEwyRaJgTDqlXiEAzBR
Ajpc5SdwvqEBSaxbKl8pjxVSxoIRL+gCKDezFeEv/wZ1h7J054353MFbidxlJ3M/TnaKH7sqAjT+
xVixnCt0BR4ptDOtEFKseIZ53wSzYKpmDtS42Igb+qHuc58jI16oOOksil495G0GZqWGQhfTFcMF
cPZ67wKW4cl6VhcPqkoDJnNJu7zrs7vr/bReKGpwjURevalrOkWgWZxpEXiVoekoH3wg9cWWROrq
S5vMy7himZBQnog6HRjx1j4ujzG2PvIuSYd1/8K954nBrzWAtjVGrWLyFLGInyVh5H646WqbPGCU
M8h/M4HCi4JZLZFDV8MMQLx+vv45mfbMAgdS9UvfT/XjaFIqO0IOiPIUKINCp/D9IsQAaxtk3czj
ZOsvaOhKm4OhDUI/pt5vYzRWrO/56c6Il3zEqITqvW/PB2Hg5c++cXjWwwSZA9OdmQeyWeEjyae8
KEXp41wmyesnTnm77mjWJF0Zg0dpHwUpfEPcXVk30rU8K5jwfJuFGsFLkadWFLMwoeLCLT57/hdZ
2LmlWl68Z3eWMRdyYFotMYjpDQwVsP0iPVxVuIPEzYl6njQJMTaE+jfT7Efbgzf+wjkhUwFKR2sU
le1UWDhlG64U2PIiXwaNqyviA8Q7av4TAVnIDrWOequZxfTLYc5UwkYRsDMfc0VqSq9R3HT74O85
hMlB4S3X0LYo0mT8hRVWapjELOzRZNKGu2ZokUV8QcetfYyRT4h49As++YFHCtTOAYPE62t5WX5K
PIOWH314QBOlNd8KrEP6yj91gGujPHZjzmhwGu/cBiOKApHA9C086WKY/xPQtogX9LvuFhnVSbwQ
cM1+L/o+Rpwc08N87fGSDcrnOzMZMLxWCnUaQZUDggS9dHjR9boUbPFaJEoYZEXcORGlj/nX/kwn
N+VKXkO/HUcScVsqCSTvePrAiDW9a/s4E944+TazqI+tmKToVtjZqhITstecyXsxn/1IWETs1qPe
vcurQDYRrMh242kOsReBr3L2Rs3t2QVEsOkUBzE40XZWJrlo0TcwkIDDwvIrRNF79xMyNFFS5yEo
AW3PmdkfBEwFhKprpQgOnNtEbTKnAQL8Yq7FyyTW0GMXslVNgesf15F2F+ny7zc/uPoh4pJ2mKAM
KuwuQ52UQD0sxEXSLERBnr7qiLxfHqYPqJKD3hLkgrq15xJWuczCxpr8rgXwm5cKXfwiAwNbMGmU
H37SLnKq4ayUXxHD/l5CnW2mIfjN9gmreO9srjgYyXZGMjWxQhtT9sk9X+Tf44V+LH0LXkvBOL6p
ugUm6yrpj53EZ4po77I8aFAGOFUzkVCMpLFal1nfMzDte6uGZuxCleg42IDgHdnMrFKhamy3YOIE
B2YPUT1+0+Bau/vHAjgG1oBtEQrHury6Zlz9IHE7AdDcp+ph5FEwxLgdx7uofaJmaJpzsokrHr5E
mvvJxbqQR+xT1BhWa7YAY+KCzJetJll6TRWrqwAfAYnnXRn8boy0uzUTDHrJKSgBhdN7SVvdFS+a
0O/yDBy/kQXwf/I8fgK142YXOrGZBxiP1RQMNtZit2afiZ48AqJdfaTvGIXvmjMkqn6rEFyEkvJO
ah0/Gckni3kAp/FDTKsOG5rfefabFibz/OlxY0SVsDh+vnYgV50VakOj+ZC5tN99oQWh6m+qs/Ej
zlc0GfPQEQJP/TsuTUIsJKTXH8Vn2HIgEh0Uhc8X9DAwKX9yX6DOmMSNQzKCKtCUR8ZfwmJeYopg
xC9xd8vpHN7H7EcR8Pjjq2XWXlW1mqTofwIFb9MxQ13XmQe1fvQn2VonXKq+GsXlRuK0TXfai7z0
2qEn7bEg79SegQtJjcjXqAlgx8Rd+hl4czcx6tZRruAEg7tCk05o0yMY4bhuaYj6knWzJL8393Gb
QSAAjZJngemsLlcbQQaWpytMcQRgKD98netxG4qESSi5H2nYJUXnoFQcjgj3O/YpFs8gsyU2SVhk
2mLKE4mWGqR8q3GtvvhsE61fQbJ2VzXRXl/JnjL+2jNOPzdmkqiPMepufSAdyRZiYAVuAcqJnn4n
X5z3VIDIpFFcWnWOSuuB6oRPJAO7WBUmun0B5mTfSkk+5AVUChUKb4U23eifTRLL2fTqKPzb1pKV
JxVawkKFEmIO9kJ7/6zOKqB+rk2dFxv0LXY7r+rFL6kM8F4Ayd+fLW0HNjWVxjjLKLjKhF3zg1TY
aiPK2FpVaRgQzH9a0iXA3IcWsihHNxbkeD606WUB/J1ytsu09gTs7Hu5BM3zx6Kbe5LvzVe3/tJr
+4CzaDHheHE7XZtuyaVh79rBxpnfR3g/+Pw4XcbJhgrQR/R1hLY1F3y2FhTmXRyD6s2K8l7anSQ4
DSoXCWkM/zByLsN5uK3FsLpJ2uTe33oRKmxWGuDhmvilJzVJ9yJyCf5fU2FUJ5w7lt7oTitIK+IU
n3oZkqv8r6SzTVaQR8fktdZPKq5z23R8h7b76qdyuQsafVz4jPz9bjRnAVHEHwSmKPQJ71gAS+qV
mQ0WEJMuq5nawG3R5/g0vbN/R9hJ1HjnbDRtdX7tswkU2QjdLqiaDp7uNBKNhUVSG5DaN4eUBosh
PLPJbe27Ik0kK+bWMNhP5tMJHI62mvKoNZD/Nw5dURBRtsbQG05fDWxXqk0+bObHJBJKbXGxgLYE
U1/Dbe/uN2WC8Z1grI7BaQnno+2HTzlbENhPO50uZNEkezRoaTxGNPCdI6Z1Q2lZ5UnnyzaQ/IXH
8rNFC+bols755OYPGic0GAOQXOdsSpHssUi9pp6Lw9xUfqyixQR+LcCiWkCELlup8WaI7gg8R2fD
EX9eQ2+I/gIzJpgOTlm66AoOy0//h3ZTVOliXTtNOfm2AInHVSIepPU8A7oSpgNg6vAS9WRwy2IY
39v0FwpCIy+0qLkc/gLgkkQ7oH+NB2Uocjbz4vxLnSOUMmXXW5IbZI0Kh//ePa8MXRhGv3w6YFLC
84kctHgNAD8NndMVvlygtC2phWQGUk/su24m+6+u/uiyU5asZz7c86kQtU6nqINkMxl+gxdUypYr
FU3d2sst7ExVaYcZSyKFttzeQrMRI8TW2EA8bkSFZf472WmAACCZnd90eqykp56HxVnVF2aPCk9y
RQMOojkizPKq3rg5WW68bqy8YXAsByRU9AegONULisI15EIp5QMe8wseHaFNcO6bU4HrS7PYhWQg
1fchlfaIRgSxEO44N4FALNqUWGl5JNPL3odStbmBdACkirmffE+O2KH6xzWRFnBMIk3aQVdWIiYP
naFoeNgmTueqHGT+ULKtF3PRyGa/Ene7vkdQkdCQgyUnOqlNXLZbuxWV9kCZXXgWIMbxYmBaINOq
9rFDNaPUtOu4wH415+4piHU5vlpXdjG6o0P9b80xteMnz/DJxxXa0HRRj41GFXcrFB3XRUq7vN2R
R98Snlmqm3b/5T1c3q/iaqz83EHcBmS/vErFVrgkmmUYGK/yl9FRKTpnf8kGh9DxNxBPuavyHpev
GLN8FfOL4WPtPhDBWNc5jCUk4CyZGQU1fNqwwI76PsG+a7k3+3WkPsYuah6pelT48kx8lZHbV6zy
kxSfICHNga7JJDw91gDPcEjFo/gMEj9FVgkA1+QnP18IQiTGPI5e7QDJF0OAZwRPQl6KLb20R+d3
eNGk+la1O3B/dfnhAobRXVITSI18RHAGH0V9qgBuisoXgJQ9Xauj3OBbswBdbY2obh+B8T3L8M49
BCrKfYLNDiLu43pYf6f7gKVEsdv2yOejUlf0xwgfJDPW9tcloGQEmkFrrTrwk2WrNw+YjdzemUQW
00+hgwBxg9gHyCkdhlj2kQe646Y1gFybv23Mi4a/Dguv+ziZYRNLcFiFAehUEmG1Eu5n1cmNlG0H
hRHtOKmvJIHjf3II7iPW74SD48knRpE8qD5PKMjEFHL/jV35uRNVCrtJLmzoIqBhYn7h2HrBquJ9
ZYn8w58UIJtXGXxPIwvRUV29pYEIM6vbbkICXcJCn1sloTY9LZAsbvgQeCeNeqGcYf0PGFC7mV2k
oYQKUBYTnmvaqJQ/9L0isRvFgnZ1caCWCMf1VWUV4fkIc701qcYZ5fTwercUbXhw/MUU0G8yUncO
k5AD51eccZZN2hf+2tAwo+y5aksTzD0A6vMeLdBkTFsFnkP2yRqx1VBOE7F4Go55EtkYxLBf5yT3
wtuxs2XeQWWmo1NyCu1FvxXc2gmKVYp1WJrVY3G8eU17kYeecB34czHopKnRlLYpBJJhH8VV7Rdr
5QhBxyMqFR8zsVM5om/Dq3FHPDjVVsaTOZzyaQGnC/Qjg0h0RtSPCrZrfvqpyQppdBG7TTcpHO1M
uNATjgUg0m6/oTJD7+025n5LQrbn9G1q7W3eIcLgSvIilOjS8K1DkBvNK5J7pmexwrwZCIRYzup+
I73koHpDgOFkvp36hxXMWmqbE3RuQNAiPlzEuOQA8cvqZ8Ib7PEeL1xY2eOa5hz9IBcbDktprh1y
2XdxO85oa63ds9XGE+Yy0pqvKh7crlpkrhBoIYPz4E+FZ8oqCGu4C4gSveVtJ2zIa6j5AvIa/HI9
+E0oZQfCIFOPtZ/8F+tvMqzjD/OMgImP4ix5+yDd/fDU72pQhL2gI6FBzwA+LOGRx2MrtbvlHlat
QkeITSgDRZRQGbXS0fldPGsjuDlbkeOAUYlMJLuoyjIhQ5JkaK7ye57xY28E+0Gqv7ahaBILjs1T
N0FP3IhNHlLVfaCEOABFQejxKKc8AmQ8wvatnRHxTuemSB4pa/0NvmbhkISMYGeeWypVv80UY0ab
WHeQ94YU5c7aO1yY5CnrNPoVbqQR2Y5VSR8gb8SZKBaiOQBnoCA7U7m3EpccF+YLRoX/buNo/aqK
fopU5kCmGyvdn8PZi9Gc4oFWHIheUkXzvf6u7UOHut0ZXXtNFQHzb2Tx96DqgGTh6I2K5/uJ8TaR
ACvO3yBwMvFtH/7G3f6PKsxvHQBxT+vhmrQspdMsuVOVBfs+Pe92CBY12ICw2+nCGywBz6bjhFON
fb57mkJs5A8kJ207DmoirTn1mVfg3Fl8KDisBOMoywqPHwN16D6kR/xoL4oRLHgbqaknY0yD0mak
Sk7G+AcgbDczRILlxGKzTvPpVx3roO5d0M13HVfh/quz6gChHfgc3b6PSOZdGljXKFJc6sTbqYzx
RzZh+zHqSc+XjcI3g82s1ge2Knu36SznTfKFIREqIbhW9qCOEaO4FMeHXtaEYjmEsr7795p9aF6g
BC1jh+3ZyBIPEu/FjwLKWB/AqxEBW9LXN/EoDzVH4gVH0ykoLZiO637fXk/o5zm/qVtKxIIUOtP9
+qMdPFbgfoKPKq/em2hM3KMC3klaF0Zez1WXL8slBMtONcoiTSPhPmyrOydHKw8b3BXXJqzwuQgj
Nn5o3ckIv5CPsEgv0NVS/OL6A9dg9H0TJsClqpugmpKfwFoKkJBungxU0jUbrHkII1barsEBAJHo
VWfDDQMnYm+4SQeZcut+gQ7q5sU97uJcHfVOjaO+BKBkoy4dqyGDxOO/stisxUmHW7yHUvZdnqEj
EKGodm9iSXbkJFEOPJaLQXIC5QbDd+FJUyJdEVGp1kVO3EWGNBWLTK3i2D83WtwPHVa4LwxVHwt9
a4DOQTSkfHUaqqGXuPRxU0ukqQTlLivNMeRsg3T1kowOFe3ir4WRdgunwwAy6x9/3cM6bL07ZzDj
cDrrfKoiuwzz7buZI9SF8oh9gPBS/w8vWl6JpYj1EAA6fAa0QitiYaqJ1BTiokivQEh3SEm8mYAx
v111+ZXXzR7OtUH7ziJomiEYeMjFApXvXlKn1PaIWr8B4+iaaxluhZWYJ+tyS4b4EEfYCdhq81Yj
8u0H0Br/YaXXCy9Qu0yJ2kJiH3m7sChgXoeSvojO2RhiheVLQsYgb57gERkHNzvd251bv1u4fIMP
3z5w8g91pO518PZbuNi2PUFCCiCcXp7vU9LjFwhwyIW5X4uNHAwqGYzLGDEOkIn6vQ6+XgWDJOk3
OU30YDIvWr4/JZIQZiV1xk9KYjGNY8y2wCwHJPueBOFk4R+6U75QCCQHNXOwZuGXTKh9387IhkSf
cuDyeGTTY4eegZFpSboMIZReCd1l5Tgch8qo+x+2qvYSgDzRUp+tkWXpDYB5Ad8n5BtbZV7BE5zH
M708nHs2VkEx4Vo8sGJrgHjf7gB82DCSrcQvlpKiJlKYn3GwShshBMENT+SK1B10h8uZwlvt8Elj
jV+pwZ7wPq0Q/+Q1GWJRPLirM2WySPxOINeP7vEOQOdHG6GQlxDSgspYHPWdUnZY7laPPMtUmaLx
a43Hru/p0x+hx0guV9NwocOWWvYW4MGNf3bcLKX1mks81pf7so0bXB/tGzw07WY+82LwpLwbM7xE
8kPg+7JRjpw28yEP89FmTqekuRVMHQkkiNVs9FGkCjHU6QK06pYyVAv4VlqhvOE8OA8n8MBxJEKf
ohNWPygwaaAc5dFM3dW+0kJI2V36BbmoEvf7GTgsANTvQMq3LqmTHOGEiHhQ4v6EusA+vgGl6Ghg
FFh0rhb+K4Uw9plLSumEiH/NdZLE28fQ9yEg26bqpb30m10GTChNh0DxCTRZbx7al8lLkqaayJLM
e98YuYN97RIQJawgnoOKRpDyB8KZbQw95FSqi6FtKejIZcC+tMc0yzs7CQVisqM9Ngs85KV2X4mx
nSxJG/c97vvZ8Y1t8mguHM/7uRdmeXDJaEzndNNTg6opl1yYKdmocshyfBZu5K/6bdcXJi6WHEpn
gJ9peule1oOq9zSJ5MCFsRNPIh82rnEw2v8ZSqrntVl+u+MKb2rXKHOd3/WkaupF5RLGckOki7iS
r7Ga3MOVa6IROb4alx5ZrVpr+6HLzlOKkBUERCIQqe4RpPlGYe5skX8EHaXkPqipPsjAPnQV9aTk
7ybW+5As34W6u7dAhaBpbR/3po0edIsoZ8oTRHwb7xoVrSeaYK4HRhcaJX534ZL+OMhribbV9Mdh
7Pqpba494w9zUUAj/cFQDUvSsUpA5R9yE8nrlR3Gin0WQLHiuGf7jNScbpkkmMHzIKX2Mr4OiiPF
HVujrxcE6O4tAdl0oyOEt7omhBjynXeLMIhbhLrj1JweOWKcoY8M1ERCH7oG2nWOpVO7bW9HBdnG
03sObpC/Oa4xTZCt4XL4EndON9HU1ABkNHYt0GC6xNrsOmqSnZta4In8BPPcEcY/yVcztFqxrfBv
NSYGUH+w80Ra4+LgVqqzglJkKOTEmpc7dDY4PhjGmQFcoPdUSn7OlQvtq4WDJllPaATltPH48F1W
fi5nqaS6YqHLmeNuXDpOL8PaX7l5Ll4rlkgrhZY8b9wyzQGlhf1kTCf8U9T0WOG2ghuBNz5BRPu3
a1c1QgYwX+kVDwXnyCVlK91FQNQ+CeX/WnsYWC3kFxSCw5IPf7cfDFSZhMuxTQf/F2S257MkzL8p
JVAFp09/iWu6r9aHoE4atBoC3HwI1hYci3n1Kb7GUxoiNafyPdR++fDXCbpUvnHI0SZrrlzGsnhW
mRLFKwadnzYw62A1zvEoF+QxoIG83chBWo9tG62ycDJHz5zO0In/lz9E67otF9IXmmkyjsmY01gi
zRWPnMCBfXp6DWmL/JCHtowft3NzU+8fK4VEXy4+8bLY/RMyJOQ+KFyBkFufwh9SEXCAdPDo7mYx
Hc9vnq0R5+KC1ftJW3rkNIczQfpQy5uPogrps01E3MycnUjhlNbhsGY+kBKTGIF1dHWWZNtTWyvZ
eTYLLlqC99AOb6pY8wCZF5u0y8MqXZdLDTYiWwU4YRPzcaSAuNfuAcWB5dNzf/M8sO9VfOxWsjiv
HRxqjw/Gp0hR7bWC7bXdezMxhjOOZQDUCzjRsr/uzvWSSYV0/pmG2Pnu9RTQk5GaL5p7erMOKY40
zwmeWQ5XM+LrpAeyzSXFlozfiDl/rORqOOwaile9z7wXUUDVYC35SlIRjUw0pePm1emdUZoh6rh8
Esv+h6BaxZk+JDmAgy5nhlNfZtP9dkTyjru5ZyFXLsSEbkE0UJJdL3TuQ3bgsW410G1f0nAhkX10
EiOu88oQ5Zb7djArLd7rbg524zxDY7CapUeMS4MkS+LbfJjXwzWVqTrkpt7yDCNkFY5mlGmAAKnD
ZFAaQVUHXd7//0262ZMnJ3UtTl8OB70ILOxkYNogldZShlrx8f9RuBX7kVr4H8hBoG1qxLsIDj21
oIy89ZbVMEfdBEJyugArOrTwR1jqtyvmm31hJUySKf9dtPjj+kHMX/2KTYwEFQwYc4rFi56NxNYl
ZppPsqabPsFlg0L+Y33OtuA23kH0FJ49aKeNLUiTtRa6LA8/OndynfB2DoSInJ0JcxNNXHLhKe9J
PpMGjH92oL9Los4SlAF4oWKx0t6DEYPTSDzNlKRO0754PF73rsclkukPVMKkLvS4WPyp6a/iEUqF
PiMi5FWatwQtCC2ch28N0Tf6ubWV282XkPsxJVt8cZAZpdxY7qGwvkkorIGwS3oAo1ktryrK+0UE
DEizyonHiOqgI+5JypQi5lm2slxNkIbKO5tK1OkOOYMaxfG97exgVJluRTyons9iBCOQuyMyFb0w
RGXalvexlMGqJuUswIe1Ij5a+6VcoF607OlugPoy9497bDC9scOq4SmL1yVKXi+LZeGie2LHNADG
C39RJkU0VCzOg5Kez1+QmbvYXB+mukp62KYFlDGVuy6QhXfdqKczrcqb39uNE2LfUgHtfFv6WxEN
jNk7J00aEDZxudJoQKT0D80pl6GH0xtLkUu5qrFNiH++I3o6zd0To700Sw2YtvGJq0wO0qFxHqmR
bmtXKp2kXeEzq3YD3DNnzNZYSjVaHnue3gv7il/wfPBDBHnVWuOgZsog59SoR1T5COaoQDM1DvUC
RtgW4HYpsRcHmmYf3dS1vZZXlF8LmKyrX4Lpl21ipG1JqNxeElElMBry0wlUwJX13kUMBzR4wcWB
h+bgZRJ60v2eQzH2+lg9b0Qhzm4IbdwwHXC2VrT/2K0iV1w8QUXw0UHMKdNuOeMbRuMdofMImBPM
Fqei+Sz2H3epYJXuHBmqKye1FHkomVDXh4jvmfslxOT4vfmFfLAPcUGJJ84aHhfhrGhCWNdmipYt
8xOTt1F4I1xKnLuHu+4MIIIelQqFjn+XA1pwtCfFjC7h3j0zQWncIvGcgyZcSX4lQJZiFgBYzeSf
cfIKmm3Bk/q1LQ29s/SMHjeYhRRN6jvf3G0rGzUdvPT1/1ZJ1m2sLJU78btsujRo8TDttftpLvgR
aZiKEnZFl5309k3PzQJNuR2pSj8ACubVjIWuM72jZk8yKWvTomBlh2Q/epmWpTuYWTyKZpht5uIh
GnZPBydG+C5yqfSvfGQAF13AqAO1Uf7yXtKUsWbMEaEBSjnFPu4XZdFd1k0iyYjVeRO/EsOUpRWJ
d1O1Zq/Xqko26VE1ls/RDbxPT4OQG1Vs1wUFbtDt6ghNCmlPe2n/diZF4hnJkmZy25WpxAjFnmX5
LPP4Db7gxlPlT44/4rIylgoZQ4ox3pUZIURo4UxN1L77/2AQIkLnIk2OHkkpJuxAaBlcZll7x3vX
gfmEiRWlMybXNaXmk4EiiOURtLsuXumLK0NcXxbYxizKPasa8Xz++Xwz17vuB7AMHQoNuDhGNnoV
bH7QgVycwmWaofXOez1+BAPeRpHLIw1m2K6fPrA7pZjBMkzLiqwOcVdIStqD+rPEZ/r/zYO54bTS
vj8rd1I8l8t7R+nGGx9hNokyTQIdV+0xtnuKmwb70iLjrOVXf9NeWDeyN1CcV5I37pbDI6TIptsp
wg6xAQAdbPG7MgsyfstGTuMtFH+bVox4mVqIxgy98BkVqUAntPPFV52A+kdtf/4q6faqUTAWdurY
m888L6nQAMp5sBSDHHYl5/VbmKQYN6pstsp0y3VL8mVpHKQQr1Iets2EqrP752djRjZ6OYpM4NFM
MuOQ0DHsbEP7sMfgSY7QF40w0Bhlgh4iU2zVRQ0aY0n9S/Jhu1jMWfi6fhUTBajNcmydlax4wijY
w3LGGRAOz2aKLH3+q97NE1guJshVoEoD+XNQmGLEBWHZ+wkRL/OjzaRZeXdsgFwpK1UdVqLIoaLh
yIg3PNxxK5Yg5ozQQzFLJfG6HWQ5eWA5Ni5NHHBF9BLHduNimiH72+rUEmwVARUQTOm7bAKfJ/aY
qXQ/XtmUlWge6nI3pv+/exedlIHW/P8iWrfZX0r2SJplvCN6xFkfrTarfpqo6GQiXbJiMj2ioRv/
shIsh2cwW5EYcRvm+46slmc+ZC+DDqR7y9vq6EPnW5dS/2KNPTSkiZbd0lFuSQvtQJ9ZmkNOh/w8
GcbfhBzqA/LBqzMkdZQM5u2cDY1+LfG8rkWEhtxhYfP6syMNGStKI6LYiNoyTEhcDGvmM81NcSxg
TFyTKGbm9JgfuWoJ8SUBoyilzpTZOCUEOuIq9AMUQrbaxt2MSMBKqLOKt7r3Ns00M+e/KM5kCxqp
Ynfdz4EaVkILk+NBo2Ylv7CNA/TE5XIH/yR72CN4UEM/0VNZdtRqWuIQ8CF4xN/OttUVGi5L5nzm
Hn/20nc6IzzbEO9SL2WIUnVYILD6gd3PDeCaR/2or5qIBJiY+aR3r2dwYjg9BPGVJBgoAIJhnibh
H0hZ/JgZ+X/Cblml7K9/c0g+qAl394c7y13QkZMw9damaYkOdyxUZhWuEDL3Gqu7t18UNMtJzKDQ
Qt+QcDPSgPdQ00jQpn3N3MlUTfzs0FxjzkWz2G2VHJar9P4mk885qTc+o0gBIOyqgaPNbg9NDJfs
fs5+EelTqLbxDxQV3+ZizVA8CAtNqRxc3RnZ37frruvAqyi5x3BRZ68ojne7bN4kmqqPnGLhUFjk
DJDQW59S2OTovBwkPY1xQhvx1TSKKhYySEKz4/kApfzigIUKTX/Q+P+q/yzJQOjbJJW/pLHUdvsM
V5DoCpZb6nBu+K678YU6RWUAWmriZ7kBsMd4P4McFtDaPbWWZ1k3Scft23N+ANcgGzjnUj23TjGo
JV8O1RfOS1dfBBVGzn2JGZffeLxNlc26JVPncW//yXhi8A1CKi8s92Xf6YdMrWbjrvErTolMiZw6
rGXp4jdLd8dSBl8jgThOVfsGDfYM+dcNQR5QbYPXuVbQIPKg4j2VBor8zKbnTPIeqa+3Dx2lujkJ
dibaWbF4ZBD1LVV1+7kuWvZnDO8lobiG7bk7Z8tElJyfvQHH+3a25FNQRtduT+Pm3xwYr3QDkIvV
YQj0Nh8/c/ZTuX4s8TDrhym+cD+EwQhKq8mWMqvyKnfDWstvz4+KjAXRe+D1PtnXgl5v6gUfR1qO
+WhTd6dV8BM8CKMNFQgNmBR44AEu1OLKHr+7KLv3x3SNunrbbowno2Kb1VkT690D2g48fl8lrsna
pF46pOvm5qvBkDlExv997cuNma+CJ94zlnRxKCqJj210j4m8g0Wtyi7Gqc1bPyinQZg3sHPCG6xr
6AenQ7lQcfnd+970ganSov9HI8TmRpRv6M9q8xv8/1bLlqOubKG754ZzLpNH1wRcrZY+e5/k3BXO
bMrdz+RICiZlXwSo2yfkwhiYF+eIbyDMe1sbhwlmeANg+EizzM2qwWLSbWh3Aq6aetoADlqPVViC
TEBtOaLSm9x3FdgHyi0ReITZOxIaolTaNlRHgzC9wVYYzNsFrTnmJ/bxzrSPuxs0FuDkC5MmDtq/
sS7FjI8CPnAkeZ9A84U3De1FYzlYzZFXfYea9ObjvVQZxBY8NcLO/0ziBdRL2SZxgIA1zC83cepP
7gCSE00K3wup+waGTWJz6YIMWATQpqg3GZ3G0MgJZYG7DHjRYGjTtajjhzHuPzr4Y8frfChoEMxa
3CRqTOLUDRq3XBsntFTEXZmPSs3Z63LytES8St2xtzPr/5eFV0YvxY8C1IV1232gRusERnC3S+Ni
CZA+F8J3h0AM5xEri6fyeLJ8bnCnBPXszfxnYS9VJ9U13euRPeApHGCC6kGacRWVPkA1IJM9cDAB
y51ePlf5gNq1/IHZySRRQZNX+XCspu5ZxcJqb0uvqD236KTr1DZAI1/pO/jepNGjPFTVclsr19Vo
oK20GJ9c8FqK96n/hcwZiqhdrZq7ra9Ur0X0CaHvDhZoKW9D+ykc6VHb1pvtHZhOKIv1LMOYGEMk
dGk9Eflw+x0uMAbK3rpKuBtqvYLrARC0380+18t+JuTJwSngpsRftv3gewJQcqFBK1mr0mtfQPo2
2iZrSbdmq5KAPvpBItEaFSNhRgSyRkq3waiBbe+HHAh6zV+L3V1JBvq8zSLyaFDfavNxgXBfRPz7
bdJubfXg1yD9ZX0JZUwgxTAuK1yh5X8T5kze7AflDnxi+0qJHM6qDTLk1ICdD8OG9VOfpQy4kjTG
/qlrQQA0f9fGvMlEOZpQPfRgJurktdq4BkL1T2LkKqprq6dH/m/VfZL3Q0FN0dJXQa9WmSXiVozm
WpMuMoAELfHaQ8CoDFGqT1ok+VgXxsnbWdl3dpapsPcSMsn3fB5QWqZ8sYtPvCY5nNUpSH/JWnj1
YtAR9eLq5YCgU8WVcepMD7NAXACjzmYd6+9ape2BQKunnkQThg9jsppeBzynxrayAclbkiKs34Wn
aX1IA0bFQc3REYwpEatOkgEsqt6Bwit78eIoN5ctFGRXS0K5HyZ10u8DHp0v7rEsi5AxKummE/O6
vKZGeg7oR4yJ3ifioivhepqJPWZuBhrrL75eWyqomI6Fv2XQA7247nodCSltYV1MrFXOrUBTyltk
WW/cFVCwn56jGZt00boNzFh/aklBz75W6kDSG86ce9F01IqcgaMAWgxEPO1M9SwUoaeHrxamrWxf
6ninx0Ot+QZiHX+HNlENNZSRz5cA0Ng1CJneX+PEHumpfL/622pCDF0ZsjaCAuPaGlb1iPMJE869
IjiQ6DA7zy2OvsfrJKrvfXZbqiDuF3llZ8AVNwjyf77QjG5mLBCq5LA7tkqezw6/9XxKLhg1r/Yc
lSzED3xmd8ByA/vKHEFtLBPU+iJ2qRK4dxSnD5tRdJc/H3vHvbRdx2sLUd/fgiyRKoaQD6BSxoAK
zCNdhVvDVgUOTTCwKpCM2iv585TCOs43NkLDdpgQq7y1L3SadGdfAVC7D2VyyalvO8KW/G9iPiuv
kp4oX6Q+AecN5KqO72W4vOzBKz2aZg05//Y8jzLkW2JyXP1vPc1XzQ1fDk1WM1REXIyk41UWMhnL
dMHMxM0wJ4LhAqNO9GVALcuYz80lMjX/9aLdicZKTsJNHHxIrrCm9iHnZL7z1LGIimXXyatASq0o
Psi7II4jF5TK03Ns6jYTENrySWkSv6GgMI43v9uXEJz9TqwbHmEgaJH7CGWU+pBzfr1Z/8/7MaSV
A1YibfHQuVBfv04RTs0C8jOxkWJILCFMcXNWpCTGWAvej1GDDgpjgFmeskJSqnrwQXdy//NY6f+Q
tiWNqcEM0Id7Zit71PNw1mQ/sxekCd7UZ1pCFCrzlWcTdNu/3yfK2v8yaHQsMX3C3LFBzz1Z4rMC
/jHPe9W0fV6i32aX9hcxDwD0pl9noJfnTpmctdTDf9JGqZnQEdDiy3O0F+1fsuP3cgy6SxA3AVy4
nVLCO5Jk/lqNB9lnTikjzk/qLDFpaRrbwab8FGhlCaJktVymPSPaPzmH9o49ErfoxHCgwAaHM2Pk
AzmVGAX5VvrYc+nOb0sBom7S7u1s5ycN3WayA8Z5KMcVj4YhEEk33SWQi0Ldx9XblBuJ4DLlNHYT
Hd5GuiihvRIAP0cww7q2Zdtyw9knPztQ8qP9G/XUg2kUVxOrPo1MFDhCC0CafGGo0tYhqwvugyKn
+enbO2SJ6O7A8v40CFElSyzotNJNIL8Dp1ua3hsXGcGA9I577txQfdQ5PR+jwYH8Yy4dQfZD8/tP
ba+Nou1m/AWUEYVntckqAMKem9FT/F1tZqASaYljDkNEkeUhctmvfDUu8+x3EynnCJ0lFVWx1eGx
k94fbPvI3YWX72SCdg9O034blb54/50Qx4kbLvHxjig5e3Ng2ztNnT3s2vjtR7ezQlfrQx0IQdCh
KjQWHa2qvoBCNGMYEtsK3Izbv9qEGP4HqFiV6O7c48V+wr0ZjCv5e/X127c+jMZfArT8h5D/A8r1
CNnXGBWTsdmthihsvLGLDuJgJuuAPmOEk5MXllDkApaed8E/RAeBze2cgpTEW8OmtlCD5zYEnIOg
+myGNbzjAD2Yxdcftndvc4jag5X9H5E/eveBd91o+OLf32Ai4FpEcxf5WBIpLGvPniuTT56lt7CH
NMOWIWB1qCs3f6x05QMuWOUpaPg+8LPELSPeN/rPv/FKP6HsjgaYRWu7VZQTy88KAUaVdGRA5Oa2
a2n1hVFs+sOammdiQaznN5LtmQOH600rRMtkdWP8VEOUC9T4x2Al41+Z4Ww5rc/abeFKZ8OvmBTn
SENc1YjYkJftKPsPz1Vc238psao4PjpuEDnUD8H5ikftCNjZh7ZlVoAT624F3xGbvOgiLgDknctQ
Gy9Jt1eKKNBNuxjKW1ZSdplEMvs+trHCF1m1phs6saWzuWAQUnIfIbcS2S3Re4HVYYuTmzHYjtn7
TbOJGBp/7/bAnYqVQBcv0nQEm/qQoIoJVDYMe3D7e43/AOaYEK2zn5VtNqqc1EhJnHMS9sdCbfRo
gpoeqqLuI+KNrlM17zEOujFX4fFkpPHdmq+g6EfbcDxrZoK0M4HTLVxEl23tIbqQzvebAUmBWc3z
o/nfyswGyQtUAZU1CQTYKY0rrNFZ7UtYJ+bOP5i0olvj9Gn0S3xBX4/Mgmv3lrIZEaivHgkrepR2
o1vH9m0TCixf7i/HxmO6ujTrdbweEb+k3dB6d3sAoELXr9SnEbHIIacjhw3ePSlaEf0Q0zWIaev8
9mYHI94LzcEYH9c+8gIRhBYy5AEQ7j4ivKhz+RKGR7rBM2atbgRv4Psr7xB6CEFNug5A51GVmQzF
01BLVSO84XfcEsCMuZHoZWisqZXaIpF/DPgrEOaQjCcjcA8haZ1WqXy0zm6WTWKsH7goWm/kxMmp
u3dpECtWnCw9GLAJtIvGNkA7Q6zkyhe9Ta/ZRxeKp8X1aGSPAvk9+PZViTHl40GRsXJAEBaM+q9Q
SP8iXkqeNV73cGs7Ia6/tiUXJgahJQiJMzij35GpJiJ5I/ESMxF6rY6Q0lJLLnmSc5NUtOoFvEPF
tVLc+7q+kWlz9MqclPOMzljy9KrFDTmyJ7600KZwHu65yh/y9MUR7Pv5YKKGg+/3fce+ygrIPJ/E
Fe9EC+KVK6IpxK7NhLZj5SA7JmA299eSD0vQ8aHZWwxAlaz0L1CwvSgGGreihP05ZwwSoGmTmZBK
lKVh02i1mU0gQz/zigvIO3Xi5bDNpIunkWo0tcYbazM1txCt8ydjjlFkMHDjzc1N170vCek+zfPE
7+M2EErC7k3OkBUzbUG9sniVu+9roVbygKyma7do0ryig7iKC3cKE8K9AvmGBC0W/bHIAcE6grC9
ry6GsET5jNuFZH6M1a1F4xZ6AHO63dWLBg78C2ww3G9+aJyASU7hEFB8s7TOVXR1UIXz1FP8hTFU
IP/K4AmBalPyTA3KbSYwcDSHRvN9H8zFXgcc9rJvuRwSwvDu5BGAd5Rav1DmWS9e/jjFikQmySqq
DuW1hV3w5V6qFediQd60Cf7LQMrf0bVv56JcPNsJm7EZJXkkrNE5lhtNgtVGLsPXuwVuU2mJnDOI
L54r0x3zV2gvc2xLE+ndyIuqDQiaAvsRReDmByURFVgxdvoq7SmMA1MFpHUYPYh1YBKFIsIuF7B3
In3xJlXH/sIpwYcP2GDHRaMlrUZZ7bUC3NGTLOl9pdw+hr3JfxO/HG/G9j8gFVxX7Qcp9o0ufXU/
lI3nuns3gk1uhsf9wZ+JVsBExum3ratsbTUNnaKxY9jiev7ca6WLe6b+X7aa60A53sMtgyzxZhJ9
Qr3igaP83O97+QBs3bZY4dhGMzsAjKOMQgdbqKSKNjP7tiGhqRAH8p6aOXE8nM+FC/cPwTVH9j7H
jhSUO8Je39eZf+AjVN36cF6PZK2v1b9ytaXS3TzrPqufCmwceqg1WXpwe7iaYHERqCi+2i9te/jm
IjHyKTb+aqbsf9Xw8EaNPUInxdKX4plycamHXpse59+p6RUOMfa5Au0qJwSBGE1SVcc+iIdCysAk
KSOUVgzdAy+BmwN2n0SJfjtS03XEQvJNZ3Ys0beSUlqewB9EkafpHsOXWs7ouE7PZqFykC+V+hQR
JNsT3cgugBojkH4kSGJm68uzk5blvqwHlFCnPhrhnPEM2oBFEkndq+1llwV3jCQroNxBMH/J9XxE
A+r4ZfsbXrjqe8duDIbpRuoOgmVW0jbYzGB+VWs7GiSjjsLplW1MrmkcgAwm7yO4AO16wFjtc4XI
i8yxLDhfpU1Wa/dbohgMclzk+wdp6J5yWlmt7ELTqwHO/mnL10zMZUFNf66yuMhphN9dnu57GyUi
Gr/RRKch7X4KkTuBRtSTV6OBz4NT/E0q4v1V6Q29HfVmhaOEkgMB8V6gSoFqQMX4KOeJGykN0tMX
BLFKErDlnM2t0UFgXTaz9Q0ymJC66qqRvS5iyJFE1mT4frpNrX38FipTuAKIDBFwl41/CuzNgYeM
ajKGuBmn4GECq4LDSXT/D8n4JgxS79pzSgXqRevUvfZCaKfjknNyAc5GZQaIay8YWLgEQ+hglmTJ
KBITu3EtHfC6BLVbspWHy1RKy2ZEKmNWlliq0V+j1WCUfyQgw/4peX5e3SUYZ5dzNIbstAC2RGu4
oMFbrpwHI+lYKhd9E7hU3TzOOJjMW/YL2G4ZUpcSr/sRDjPiNhJ4Lp0/XMKmezATL+TvLIyEExNG
0Ux3umDEs81c3ZL+aoah+32pfB6cR1Hdg+yWtrUtztlIIKif/Mr7McSc93QYezJ+L4KQ+q8scBei
aViVw55YwRXOI2oXskwWkF0KQs1r2EPsucC6YsaIRMebrSC1nGE6r08atA0SgZoJVbq0DT2SbdJv
UpUREHEdR8UeVRHiPcXq4Ly2xxSJTsabaO/YkCZ5nhbq4ptqm+NOFqPGZzBtowd5TEiHZSJzTnoS
70s8b4Rtbekb4WydhodWOaejbog7BnIVbEBZINC3XJfr7HD4xk+oj7LE2OIQZasxxlDSnyCGtRxM
zuakNdEqmq37qo5bn3vY/z4qyFWCJHcNDlhNqJ2hhEHqzSoG+C4cG78o2TxICdsAyBBM54TL9uwi
H9fLFzUwcu0vfIVimFQhNl5/3+vsyT+SrOUxYHOLtXx0JXkRTxh3WSc4tQYSU2FhCDqTDvqKABX7
ixnhi8G7fDDpOAaeeVySJHMpm4iRfIGuh4sgaChh10EFFHDG0jHdwHe4eBczEDgQGCR+E30KJSlC
uUzmr7izTh31Y6guGoEKMo9bFWkXNCri+K0BUZadbNw4aTHlQaH7udOW4rwldHgHdwJraRMiU5VS
e68X8yiaVlz11s0U9Umr//1LrnmIU2TNxlkrES9cMBtR692cF/KCsZjQU50IDisuDEYrW/nIpGLE
3dKErl7IZp7aEYkkcqnN2SxgbnBPoFK+XiskVqR68OTaQiWkjc1OhK7hSMsr5u/RP49MruZmqhmv
KhKm47zISk3POW+fBkbaAJqrIonyJH2YcvSFjURoJItxhRJ5hE1KJmqBTo6TfuAiEhXCZXgLxUgK
JuS2il3IEXRSLyzfSufhQ5oA3b2a3X7vOY2V8pyCKZTf6p+isceVC3XsPhCELfrndwDZjJCBg4kS
SGvdWZD5kkLwLL07GSkgw53D47b+wqBKXa0jClqfotpTKZ1+qffXPWhD+2JqX1vSbVMwfKlAgJYq
70NfpSmJL4VK800+DmtstA/jdj3kBzq/mTFhwxgryZKSGXw8cwesKDI3ohI0kK6TmT6VZ1cGtWVf
rp3gJ4i/sf+vFV+M9WHeOCPoVeiKh5Hmo6sSNUEmFBJpnltm8WSU0fCJ3dZo4u0jPwtMA+g/aD6T
zDEN18nRgvI1SDFgJnwASwBxrmaO2nou8XSuYsmnsIcayRGMG2GF/5aBD4vFKnhAFnQ6e4upJv3l
s7XVHZZyN8VBX8sKNByRGygX5MncOoAYvJ9++H/s1D3D4kPCdp9wBSVkp11l2iMEUKTSx5vty2uD
/IMX/TxYkhKfsF0qml9PjZg1+oE1nmjEKrJO5vBeJoQfcn/DI+M/kejPikWymHf8uQIbG0XfZGrY
C5ArubscHO56+kzVWauv6G7Q2pZJ8SxUKFOOFfYIgEFykhEnQg2LhjvLqaoPoLPt/tum6nsfkcvT
h93akVq0g3K07JiofaTWOq36w0UZpZ/aSlA55ySbffq3PjxrSjvoHB1b2ErkuKSDQAjvJ/j9Yvim
xTRTxz33E43UpO3vrdG+WQ/mDiSmdxTqyNo6J+HTezwd3CaOuMsOY1jT+rKZZhkFOFOPG8zpQ5pj
pKy6i+Z8j4DZ+nW988h0SYnIBAtWcz/P0G5wd+kA5Ps+sK0wvFJNWcUwBp8cB3pFswWKXhOnOBq9
zthN5uBlPIb98Bbm3HDXC7Ka9VdiTo1IlnmZfGEQtXks9+Bk5YWZ4zPg9+Wu9u/6k8YBUr/4k3Hn
l00Wh79eyq5rPS2BmgTt3x1T/v7IeNbyCEX+pmLCi9YfasjG4//dEoWsiZyG6ecSLtsSRjTUcjgB
Dc2CavcpjQJejncfJOLXn5018NCVlF2V8wkbC9zEMcBs6ux8tl8xpQCSlkKwMxZayk4FjtQ0r1u/
CM1E1jxR2wqir4EqjxvnVw5yNvXkolJZYsXV2p8KzDwc/6+vbH8AHY5p8/a2SU6Q9Gl5V/WPkHOa
2eVc3yurXsvqo/8HBk+gg9qs+Z5Oehv1eoOoDcavSVOY/TFqWHSyBv18zBaJfPkfNQmo4GlNkuR6
QKEJe+6xo1NkoWwpsp4OI4tyl3Y4Gvo5lAzzhfpJiV0xDpWNapc7ZXZCRnFefA+DwwBTbYrj8AOM
OZyYRPx+RKSBIj/obu6Iz3ido04ahZ+MkWshNRQ7Lkj8BW+TDYQKqx088Kd00oytPEVgxXzGSbnP
ntOHP/cgcGFBT9wzXN+ozje8MhloSy35+Qgf2EHNob/Vkm3QW82dWaMZzOoo0W24/p82gG0vHfon
Eml4uS6ZjRJyz1OvJYapuNnSRWet6l9dqlvdEdgwC54bay5GwLOw5P4UDENlEg+kSgtf9Jun5Ss6
yE+gdMUU2YRGrDTPkWAYPDtjCxIJSKnWn71wZPhz3fE6pqwctdRFlq8iaL5YQX/Jz9NTUfuLNdlJ
22BoeLE7Ksg96J7v50sxmC+acOlCjL+HN1H+ZdEofaTC9FN0dJfs8NZ+5dRK3pIhVaXlxyJo0opr
OYE54wPbQEJ8kR7JRKcBSlFpV0m41QtpbCSAcp6a2gJ8c0DUF1NLIXbCRWA4TxYHZR0YAr8j9TJP
0iWIOSB0K5CSV9c8drYXixcSv88cURG02EVMykbQJKmxW0wHQpVa27xorBy9AAliz8wcDcVx2JBD
a+uNGR2Vi6bU6Qx4d7K3YRlPZ0Lic85+3h9jdRtbkJOwFC5bPaAVFFK+2xaKjVZNsKUB0AppPNGi
psKKMIP3zS/YwaNld75qrV81dNOD+06W08bOg7DdC07Y3V7gZmWkIrZVxQaL8qjy32omMsCMx2UJ
L0G3/RqhKz89OLrp/keEG0KRiOGUsKf0wDx+a49+4VXW3XmUxiuZagMNkajPjEgXsXnLwmlQfrj8
kYNuEIz2Ot5oRM3KFhTglP80PTsrniu8KWzLUYaoFwx0OLtauX3ajhW0N7Wl1DXhr92vWoNc/DJY
a0GpiCMXjjEeibdlvItBEo4kAUGlXYY9rYaWzGACEtYa5bg/4UTxNaJj78q9dPjUbaBIDY40GZuK
6/M5OSx+WDtMI8rymkfXHEvEEO8yZY3m+b0L8GwgobO4NNL9iYvuFXEZEcImFqk9BIIBtDAHqSAh
5Fj4rYuX01xAsBtHBQu01K0SFDc1ZvbkwqpRitSdBHunI2H7aXi1Xu/PuXFNxcVqcWfeMx8Szmsx
u5gVkaAQKPJ0aGGsOuninhzABnYvksQeb4JHnJdHAgr0QGz1Fm/ZlQOoSzHEs99RSJEL3hVJnJN3
ULbEpcrgeeeZz+Iz1D7g9H8xlVBrSHT1B7i5vbLW6oXk+0/44fR0PoRcE0a3x5AXiwSW+evK5g76
Px+QR9+se0etUSmU4JPmolRedNDQOcIaS3iVa97FovTxF6K7UJreX784wwkXMqXnf4wNBjvmUK4T
KlrpLWdeCLq1iA9AXuaMoLVmMwa67FG5Jsb2ksrdu65XX8MIgFWu1MAXAJcIOOi5OX7kwFqQ2Uzb
BEnTn7MpnEsLLnDjUNjMswRDO0B4WWWAJAbGR7/1lWL3PAiEsO5m/PlinXhV2NQBbuzbs4sROTds
X4pK5uhATaW95xuSo3Ml0QDDd+wDSggtg7dlvo/MyE1RvJMZn+ADFyA1nmkW4pCWOeVYIcoFrQaM
nUbnDDl/o2+z0KxH+PQmLXQxow7gsyyg1lqKZEMAzylebsdbvpDUQQZiDRtjBrUibFCTTitPXfUy
P/nBfw0MDLL9LuC6BFsiNL01KFK1t0da4yymeSlHY5OgSohaHxwuUxID6sWaVusB2bCcAQFqoXq+
imufPsTQqKbSFWOgE2zKFJuYx0cOgZZEbEnflk82X8nb+rRT6oiakHWR226GDs/r9sxiTHk2y61M
HESMlIlbLnLYiFxHS3ehrsdmzqgCPS1wrd7CT3qCMU6d0OAy5U8j/j6bjhhllVi7RPEjQ71VawVO
ezk6JcOeLawGwJVp3G63cRfU3aACjzE/q+wQyS3ZSrWU44B7d4jtQCQhF3cxx4fkr2emaPYjv1Ui
iWqAUeB3tR1SAOdWGuLnReWRhNTc+94LOiAzWzHUNnbEmw4u1ss+ZkdAXqgLsI8XAAvz8nr0IH7B
brgw757lOXj95CY5HD9NC7xPered1dsVqMkunLQFHfROMUbCbpr8cZtKaM8DFQbVzckQHVE7bHIm
lSLgEOLC0GM0acTuCieL+9Beb+38ZFgglaPZ1Upoo38kmvULJKqMb4ywsttMTjJh9dzD8HtiJG+m
PpDyJNSUQif2bmEgWmrBPZUizLcsNBOHpjPYRROW6sIi5OLpNTetfAYzOMwq7Uzi3s8/uKTx37c2
9TKAP+EHbUVVH2MVrXdtfhtjcSElgzBMV0hPZSNyqfgeYEjPwC/e8hQDOp5uBxEZ0T+LBTJgmvQg
1/VvCjDhw1hGxk5RaajnQjAC318sC+vHeiz56a0BJLYVUzG+eZY9Gy24K9MlBzUPWMkowWvynJ4J
heHvnLGHwNZepBqksfToXRZz99eKRI/kdowZ3zkTKtbrc7fNdSuIhHYTZf0cx52h7qIb1wSEpJd7
U/WHugZl1alBNMeYPEMVvZ4A49BVSG2BEG56zIAlrlC0q2PvAI8ZAXxehW7IRTquoZfEKvHy6nr6
9wEbx9LZdf0sfWb8veXPfl/KCdhI4uQHEdzwowwOzhG7gaSCuPbkHqAJDwcx1faaJ/lGh3uHXMK8
rPO9tYO/R8kniodLcnu5xQ1MbQALiP8sgTJJnoT/Rni/whNZNlOeRz3xBiLOYr5ppqEOh+CtFgqP
NyJ0MOMYLZkWUBNNSS83Bf5WEN/HScMR09kimUeIzGVKL9xK94P5ZizEuKlODkTWvvk3hPq+oEyQ
OgJKdkLqRg/p3/pHRsDli70mnY7zcHwORcN+Rg7ifM6aQ2iLk8xXBbbv/dZZ/+dUT/usRnyLyFms
ePBcE8M5RbTmwvSx9D7UJKbBCHUjYAlGjSJjurNtahM/8QKSbxAl8JVrOtPTv9mTbXYzrdz5QRqx
M+8SjqCcnsP3obnFOsJUSprhcGguQiAn2Fykr5LUX3Bin57RH2J8UAwCR9+HfkNDNqHbBjyiyeoL
uZNeBBlzmY9vVCSOzrKQopIFW4xOcKdkna+Y2cGsRVZMFeCTKnOR3usOFaHe3b4NAdgsPMa3ssp7
q6BDm49XFMbbHLzbL7r7nXj5yLQ/Mr7sH+hMVU5ZWCyiEHgIXgj/aXV2nOEY3OiSuakx+uSdOe4A
LAtPS+dCQxTE3ItUhMwVYbcdzFoE+nHVthMiNKUj9xwfHVC5oC2KKK+EA6VZy14CMTvCY/61vcZK
6qL3XaLS+dgq36jMXrrSsksvpi5GvM74QswdDLa8/DppGKtVbd+pvD2aJR0bCzLkNqzM6u9nUPF9
Bk8UdfAbpw/8UYuiVM9frtOwR+/fC/76B+9EGhnbJiWW81jj1kL84PONO0G5It39uy7CltVYl5is
tjpM9Ma0yM9TpNG0p+V/ssPcXaX02sb+THL9dLXyVz4iRZEhk0dIufCW0dVed6Azo1+gbRKbU72h
FDf8OVpcIVf4VXVUhsXa6mNFo5TXeBDwdDfwePhaIp9FdzKmZU2kxl1nwB7drpsWfABMS99QFp/o
Vq2QMFpF5DC/88DE39RjVWVUicofRjAeIIEEf1V+XvnsIDQW6JI+XLqZ/YukrXv1LnBatYewIdOa
BNAWx52qYMfECnhNzk8lNzcVD3QLDwYMsYUfm4zpDqixNwjTstzosm7AFTVLPQtoyMvv4LPiB60D
Kw2hIdU/6yGyKDsJxSBYqHvI+bQllEmn++fjBjkziU7prLupjTMaGuXkqpUhAmmrF1QYQFUN9vP9
5YctnpkEOn/Z4cabcQ9Paryr2dxF16ySzEM4hwiHF0HSXYuUq9IfJsNzPheLO8qgKzBNpun8Px0+
BKnH8HM30ho2UylkrzeHsTUYrXa8I5+p2PsLD8ZT9SwQcmmxrRh8chjLHFB50bA6Ce2uqwZi/59q
IIojBPaUUU5sQIOAvyAR3zu1wS730h2kA7tFwJSHoR18V18Z1sqVQ1kD22A9SLFFhJn3ydaKw1Ik
TLfSisK+0sREtVpUBETjrpN2flGGAVtiAYnPM0yP0LbKCcwjctmJG44YdAr3ZYDj6+hLKVUfxahV
cj5+t2rD8KMbVvC98Z5FKnISIT8Zwj5ftoRORWoGcKjtb2Hnk+uwbGhXxJOLZym+HMPmF10EMBZL
uEVfrCDMHqbpEMkYflEg9kYb6nuwn8KoQe49wR9anMcFAd1ZypojkWu6KzkYSP7nS7f01r5of32x
GImEPiN4NLqkvz3yaZz3vbxJ966vzs9DdogAT9iGibxPw8UISAhNzBdrN8TcTD/caYf7PtML5AeW
xMSfszy4ESlNT/W49mqI3aTzI5a6Fkhzk/fXMZR87RZ0Nh1uQh5H6+BuMXVtmR/qi5m67PeYN8bA
wLaFw5cZeXGnYBSSiPn9+TU2TkZ+jX55k46pRXk++09d9DjhyfoqHeQ2m7L7VJuNGUNPk3Fe5dOk
APwC9b57freIvM8IlcYAAOy4mKrlC0pg+JwrksXWVoM5uH2Ic3aYHYEZCewpjrFh7ksictdxXnW9
4hRTd4M+Hl+aAWBeDA0aYhSub6MyeRJU1NssWfrsQwO2bKWTcs2U2KOgtvTpPwVva0+YQPrb4LBq
6eOpwyAZLG7AP/mnYxWw6TwkFMlCRWoh1zJXyu4f1OzWTOBCfbGqFDvOz+yiHImdBaEQL6W2Y0p9
fDyXFolw7y2gZkA/nsib3ExpGgVRtycNYJ0HERft5ZN0TIHDFhrUUXeyid4NaR2X0bBXAcDonwGh
NsTLQBFFeKEjCVmq+d2Je6L5Qm/8N/LbQszfBrDUkBVZEIkOQKqXb7KnTKgSUMivDx/kXxswqvN3
DH18cliM0esxYmgjHTA/f/j0NlADNXk0xkCTI6UfJdWW0LqKlQYbFenhQ7YY0ZRCc+ATXcriNePJ
twKIG+30APvoJeWhIrJh9LeejsjASKMjgD1boaBlh8EEzdIok05QXoPkIxm0p8ZK0EUOJEpFY9dE
sk7MV7Hnip4kqCA/W3+A0cHcH5ZT4rn29+JCZ6S2d+92zZaY0vEpNtWgKiLriRop/l3W1Rp/PbPI
S6v31Lyh/+Yq3WCzsd+eT5qAjlCo92t13Kaeh16gqNlkWwvjC8cuapGHeoXWVY+ytR8FOyJwBdCz
lby3DqtBJzJQr6H/ahc8KaguvdbzllFBuJYZ8E66E2mwSfFIM1iqq+YPWKAEi4hAeHfPlK5Wx9YG
OqQEvXRi/6K1g/ggAE8oz1HpSItzScQQSfflFSpAa8HQWjWNk84pwduIJDgShF+YRUFjU8JD3HHI
ipj55dATeoGe+f+MC4iAzTb34EvOlJ9zzml2gKuqJjkjIfvc924S99eT3OhplnCn00M7xmBSkjnL
FVwXS6lZEMnVMt9jDhlXyTrjbds4w4xdPOEDm2E5slZkUZ0ge7rsd7pfoQCInNkm2hVbzO4G2qlF
X9uPGP/q0U/7OjagTfhWSrj15sMKXdBzFKv/wdgQcNjCEpIXYTbLuJ7+2GF+tFSymnbfg+271ZER
FS2r5LzzHnDzjJ064VVHiAc4fLMgDqQpk1IYfitfh1RLAocaLO0a99hGBhCxAYbJxnbWxr8hPAqp
vagdPlnKzPaHMtYf6l8SFPOH8vl7uM2rWvdEOUILQbtx4hXVZd9unSuf8+tNJ3T9uTllaVZkkva7
G4O5vVqOtZyyQzaJcJw0HZDeEBtmR/xmf1ODXtdYcH/PC2CXKPu948anc3qg5AqNWZtJVriSc3rP
xGSZOjgUtfyLc4j3RBj2q3+IRnPPGIAMs1+do5+2WahqcXyNaQjbrJVP+e5QiwtTzsiDA1VlPXz9
RDtKk5398pyx6YTFZX2pu0UrXCRy5RlExCGy52aSc8QZYSujat8mY2cGEl5Txmxl1kLxhHXgTSH6
uML4NfRMN3mYXoMFCdb4vIJDGn4UPqSeQZRr1t2etPJuTnYV6cAnfLRQQZXLdl2yNBjmTRSixXoO
NiIiI97IskDjTKz+KeCZwCsjqqUmtN2bZ54lu2KF3em1dVOMmdWqSmt1t6AJpPblD65lRrRv0w5T
S7sjqkBc2ss2hXy/JnJaGsw92TnDqqhjQDpTy4Saw6DTafBQHzbTrRn1LMfoZ2yZFIWROZSJXq7w
grO5dawNRhRJwC1joM1uesam+pmCMcmMMXNzTFpejdfBp76P+Tv84Zw3+XS8ui5XvWgoAggKABDS
T5vPRc4Nba4dyYlHa3qs+VWi6O/S7PadQJ2aF3eRHxsQU4eKntdraSOq7/lrRL4XqSPnCe/Gd3bo
OcaWCuauiIr2a33s8N3nELlBzxVNyBIwrFIHkk02FFpmwhBT79LqVBLwl8q4vypiAj6RDBTx2KBa
r/IHJlhxenbeMXv3gfIqFeVwKUzGELAnadlzrZcGJehm4FHMNAL3n1WZlck1d1arB9H5U1DLXlWX
gKgICTn6r4zEACAy3am/oVFxSYRLzz4Z5Ci6DygUevQGI98wswhKYEr2XtPuG6YZJF2WdvxnnChC
sfj/rpbr2Xo85xqwinrXIPYPNc3uvFC2Ps76u9+S/KJyz671S4LOZpkxkGK5Azyp1wzMDXwgv87j
KmJme6LXumtJC5SUSLKEEUGlHP58OaGBhR3lE4uY23KEk1RL5UBlU8TrMCRbYrs03G+oVI0oToJE
eVSQXLxizZ0/rnPHbmPis2ylpBtQ18tB89qJiWleJMTboRpb4KG7c+7yyVlMbZwj60VCH6L+UtBW
KFqkDSpauqVURQ77igMfNFw9ZLrLfCnVH5+fvbNJ7fm7Uc457EqUYCIw7DGwaxbBSP8IqyJmrWwU
B21WZxRIjB5gwEX1OPeXwxIa47JyFKTKbI5EwYXrAFOWO6ABQ+4Ya3zd4g5T6h6m5/35wM9l2VX4
eVcgrcyy19uzNr8UfKvKFjcTx9ojmzHAjh47kVrPv0nFYR4wOhpPNr5Os+b0jONZIIl0z8loKuNe
R5PMzef6JZ1qSc06vcjSQi1HUaj6x7Mygg/6FNjwJYsFj4JnP4pt63SnI+4NSOv1AUQz7gKJme0B
tcXfSL7B6K20hAg6G6t7QqfpcAfQWy7D86natjUapGguzFprKQPGJRS9YszF7VJKovMCORkNYz5p
rc+Sz1Q9YyiXiudJXDQom3wYU4esTR/t3PKu8wy9A5i1tHQX1Ylybd7qc1cy8ESfMaRFXEpthPBX
zv0Rcz9SSXyIhfAxU5KHwFzh8zB8rtHfcyYUZQNd5ZP4Amenc/6Bud7ssZVbglDA3Ugbf1Bu1AiO
JmBI5qihU9dYoD0qLNwqHHRWxCOfnyBAV6MkutrGKS9oGqvD83khDlFjA1QpokzFMYstmGNJ+/TH
8M1L4z4QDcleVeBq6wXMntc3J4/qAj5fth3c9MvvwYeN3tJfHwnaeJ4XDJEuL5m6H5rVCHRylUmD
jHX4UMqYNxJgQAe9hwTfjg+t68/Dn3jshxCzO5dgBNEGs7tvktPLDbvgI5ZkiGS7BorA1ltm0OoI
uAhbrbrRz6JPYW7rF1XrSweWd3+sdNDJk0Aaez71rzh/Nu4rM9gUNyyn0CLBohVVEmclyiX3NQys
sljpf1MhVN1WhOjE54T0WoVu+inVLpCHNgNeVzzYeO4NBeUCKrq8HBQHbnfXs7e1VLjjaMeri9Ob
f8oNmPXQrzeCP3utP8yuFP48cXjCrhvV09EGGpQdZXuFGvoTrC8boiSLrd9eGQ3F0G/CAJDU45s5
xyYVEYdt/lr0V8ExLX0nVC9Hkxn40qonfaCoqQW7GdVddgHAFmSk/Pma6CguE76iTCTPIfxQwrD3
FhoMymHRbEje0Ca0VUprLnEWICjtzrF2rtN+lXNC2mgqOICoVjTP6XoWGZ8CQVYTB3eVd3uDQiBU
Y5pa2aL/54YH3+ndCyQIdZilHDPkC6QNwKvScqSvCzJxCUZ2tqiui9bMIEwIU+y0hw83NGxjS4eQ
2EHaFRm3FsK2NY2FjWtquOVsJIy5osXjNx4oniQQqnIf0kadD0m4JLTch5CRJXjrJetEwRtFlgKU
MRPF4jpsra2mKLnUd/RxMROGR5RJTk/zro6y/OexGklLIcCK4uCCWShtL6HJVwvWCDzuhXYWyPvR
cyNjnTS3KymDgOrP0dnN7zNc9VmF57qgFuI4jdCP7Bk3CUQFLvk3pIT3/mz312/9tuSzQY33pDem
4q7sybtOJSOnIK+ptQ5RARQF1o+KJRMKGUAv9+M4oMKSe7Tg2yQjUyOAhrORx/irAY7VISTaGl77
DEWZn2/vLiZYUIlvwe3qoOdQNJFJi7IZgHKDLSWhy0ujR9GKpnEA6bR0GxxLfWQ8RgkjyGcW+m+p
+hrjLCafYfj1hjHodXdgCPcI5vVzaXOWZyzH3Wso0vPUcgOc4L/KAS/s05fny38sjtGJX6c4r20w
a7gfEgyOxRuEec3Ttp1uDk2aOYhJI2hOGYHQ6w5QcAhz7/lFxDq/x21VaZTjepsxS2BgO8P4rweC
6kpTG4MTqBer13TSKF3QBtrR2wQg5da8PLJtRSnHdUXAT3PXUkp1t+ifddu/RyoDW+ZIzYT36bfg
mcxvCbNpglieHqmuRW+xTfvR+7J35CBjAsuyXR0eMgDsx3L/anInXBegZGTlOAW9qlSbDKzCOu1j
WgN9G013nHe5BjXLe16cXydWoJjhM7dlJPv6xfwjg0MDLQBLFZ0SKSlXSbEFlKCg/ufRFDHX57k/
hiqqPYvqDtvkHVU9iDwMmF8er6e4entgqkP6acSjBH1optvB+XMZQHUM+4ajnr7Z5f0tBNYptqPD
ReXWRw8zMoVdD+GV7/y007/vWgt6lJpkz7xjQrmJRX4XdVkdBz5d0eijar8PSMprgU6eqiDB++lD
eB1TfmeZt4DDel0Yv/9IcOKjv+CMsDiPqEEPHLBONhnyGmGMdMLyxcWwaVrULqQnF4vRwX0zXJ73
qRMKcHtAlSxmxECBcsafwhQ0TgTxxeVZ3e5XHPZpiKuEu3KOi2hNc86e8X8Oc4HxkHPSjlKgWZpw
OioEgkJ6B/CZ66hctIx/EUpgWOQlRGaZifV2hYf1rm837oaPJIc/ir4GbDAs4OuHQG/FG5XlKWvU
mSUPAHmgxy2Vwsr8Ns+ctbT4qnGwwWsMjrqCdz+TWq/3HuwzhkD6FS+mL1LdNPP4f5Ev8dkQwwDJ
Ur5RRoc84MIlaJyptdsc/Q5yAM0zvovgoyCaVu9N2x+FHK9gxztHd8AHptsNfRpy6XhzFdtpKo+P
D+uOPakfTptqHyjLlqHuCu4Fx33kLukTqYKZ3U+VN0So3qI9OxAv8MKHSVahNqVF79OU5jxh8+v9
J7SRcrbF0+zOf0yDtVdqXFVxcUZ9arUdPwZuUT8j91ICzeW6eDpHCkCqOpioCPOR1cCUUU3x9U0l
w24KwIRsy0hUMRU62nlYihqjASMEBomAOH8L5lTjgwNB+ylSidT4WQ4mmFOn5GyOXtyLTc3Rs1/c
8kWdOUzJHd5wD5qFulgE6YfWmjhj/n7Bpl2hkEgqzghwqFNt2Te2qbiACGxDjUF3kZDGEhIxzr1R
iGksunNDPbuTxpRmeRs0ZKu+yjRanAhhzltvfDL3BfGyNrAPtFDK8hvI6vxdSS4faBur/u63fTqN
FcOn2WOT4XUJaIBlphIMMN0mWLUL3B2eZmrsw7o0854kxtKW/AGB6LHoHdq3DJHwdtQITBQYZZRa
J/3qa2oYgyJBY3XbWosl22D/P6CheV78bUlYXoYCQy/ue5KBazI3Qx1/bHSnGXPAKQlFpV/EkBiL
qM05A6lt1XbVoOYH8irxQLS2ldDvO+IJeiNK21Sf+4STbB21bRS9gFzFhhTov5p1H9WdrS2K8JDB
ozcVxHF7xUK5sVpBpm36h1SxWfdUTJogXkBC612ovv14FsvJmwTEYxNE31+Ba9Q2ytM9EE3iz7OX
ib+pkKnMttf1An+Le1h1FPDIkr/4abvI9XvC4c1F139vbTvq4A13BVnbfk8Ab3emsLBDFjBJiO01
3n2nGNuzYNwbsrJnYHddPHpW8EEhtyjkZwSyOMF3qa9alciAcCfvxnRMrwCKFyHfpUluJ4v98XNM
pKSsMNrNFo8v7dUHr7+SgwXFm1E0pP3qyJjLt0zOFWMlVVSf6lS3n6+pybr/mAhATBCvANNNLqdW
sM6gjFggS8mwBou2KXf/Pltg+iyE6d09yRGZ19pdK6sUI4+0+pP5GReCp/otnxyB1if5ym6RmSEO
ym7s4+YXS20Z7edC5kXoqFhqpJ8tG8lifXIF8HkVdWs/1m7qPAsX9en7gw0k2+oeBWnWS+q8eTcP
4OG68ZeJjVAV2Tz23J/39LjqSuCi/uE/qRKfSTTgMWtmffo1SKixA+Aq+5vxr6pS8G58UpJYRc3z
NSXtgR09S6LBl61KcXBsCK2WA12zClLDl0abrnwWjw6mCcqJziTk9OmqmWx0xeUYuA1Lse/TRPzD
cJsDqNQhsKsMkUhrv5zVs0aCsSkfQTrSaUGcbG7fLQGFQP7212D0aYCRPzZVRHYYiP7Isk6FUiNa
MWaZ/1nVgukT1mn8QQ4TcZq9mAr1M+AK0M6+1lwPdGNwyKllGCKzm/ER3CXWdaDzD9GyBp4TJ8Ut
TaLqflXp9XlQ+FoArqbOLFgo+kzLbf7gCfyuM8pvQ0fvQEwOkp/eooM3YDiaBpsJCizfIiUfLeNh
Pu29IBJPrY72Htb6qM5CNWgofNy24Dxn2/j5oGuIgWXWU/oCyYMZvEDeDCB+VQFpSRKejzeXPcru
EUSPFdhtKLXvB5RxWmnfJOG1Rg7hEt095qcMCAF50eheivNO+P6DBp/bb/7z+X/h1F8bts1tupEF
5bI+EWdM8xpXoaQEV3gI6KAlr20p6wKx/7KWuO1iijBthDMHwbAlrSxSYQUdaPqBLdIE4YuONZBr
SBsbUXgu7uglQv4BZjJgUn4np+5tCmX8/1GXTY7GFECbR4lcm/PvPM4kZ4XhmD+GxMHphoqlcAfF
Ockq3NadMzVQCpglz3m6JQc5FZuEnd6VTw074jn+kbWftSqCJ6wEQETLIfLvZTPk/lojE9g0VyDq
EO8klRpxyfxf1ujXR1GZZarvazrXAQNzoZ2sCec0YSm5EKLxwTmipxBHKlUFbU64l5aGdG84WOHq
8EvX4LUlIddJjzTktLHv8S8RwJdkPDteTtvVShdlWRCzqyTqQdHK8sPA7RrHQg9I1YXMks0lcf1q
FPS/7/yKCJYpj6CwpoOgWP4SR99pUXOq9DwGMZ5r+quZbrhomafT6ewX/5VEtG0hdB/zwf8EP0Vw
cSOjKXjYA07DfXgrBbOl6nFgejSwEtqkXbX0JrRIsCMWBOO8JhbzGroPPw42LpXshMArVWBrv+Dh
YeBzSHKs3cnVguU/vfcK64vuvyEe1KFJRqr+3h7Wopdmj0mVwyN7i+mn/aAXS+eWKHUmQ7usLuiq
zzSA/N/bm4QveL+O1nDxNh44gpe5kfkydQp7Nqvy6Hpk3Up+RNTS2usgjTqbVvN5dVIjQaH0Z0g8
geq2WRv/Tb90o51EE8IenW6u2/+XMQTlzjMngQYHnMebuPHnkM/YqzUQ1eGWuNZ33cNB8Cxkqf0P
9EqeTcpqglo3QZdvx0FlBM9VR0wPb+KjqbaQbwITyX59v3uTCQfWQ/lqqSX2D086ANkMhfa8AMAC
Pn622gtK9T74KgGNtLdvkTCBMHQ77QpyCaNhlh6w3bY1vjSHvRJFdV7DL2eGOAPrJF2ue8FkTKM4
HjHoVKFkfyzUf2hgOCudVLbngeUcoMZcznS2wkOKGfd5nU8psUZPTKn7vEZShi5iuunKgVgZmMQ7
1N+f/lvtkwsYzxEL0jSbgTboxPt6+R6IoUGrmzgUEh/3x0Ju4CLx4Bto2mK01xI46IPnY1jTuR95
posUQ80bphirCWPuyNvda5KOuVk9pir8zTYFFBjPMv9vonHi+qtWhsRy1RlSlCleQhCO79JL8oz2
dzKKBid5b+YZAJCSoqlgymYoA8NvMBM0rKcM6uN88LorRhuOlloYXQ7AF+10DLkeuPt7mxNbcYFD
f5XiZDYICy38PFEXlotpqSB+hvaPeotqnbjuGP345NiZzOmbPpMQPpC9pXrEPvBfguYV5WrrU6aT
B3k6hDsivPwUY1AowYYgswmpAxuMeDQft6GFV7sIYfXWDYLv0jOCctaGBFUOh/C4fA/s0R9WAbp+
Nqp2OyYyi9/L6U4gzF/PgF3JFTLZOuIMUulfb4mOPnITEKw76A9PMOsDU+ANpRIIhxhe3Y0H4U5u
fRd+vb/Kx1Yk5bYn1npFH56QgMwxR96XRMCGRm6+zCQUjlUazof1ISDIY5i1PUFg/VwCk8L3vtIg
kvfwXG0bsTmI2scfYXPrcU/+D38+2byuH7oh1QjM4vo23U6ApDWBjUwIC1PQ2b/BfrimHSecHhT5
5RldOe8XNnL8VMG9EY64HoaYE+xy/803Nnbm8h+X7i/PDRclPtvtF1WpdZQzrs4VM8UVtBnV32XB
92CX8aObMDJ6mvC4pqe1NM6yYO8Yj3TcUfpsPoJNqo0GXrsOJsc5IbKu5A1Ev7YABaxWvk2Gw6BP
cYrsiVACAFd06eYgU8uQShu8dBUuaUBdy79uGbrgd1Il1xij/cyJ05kV4a2iOqhKdJ6omJnvGaAx
1aJff5E3g5yk6mvPzbspKWXUWqd6A5jav2MYCJKPS7W6Bdfx9MbgstquG++RT2mqnmM5p7foNwx2
r5BKPS6lSwXfBzSEas+KhtAMang9hd/3PU50CgShn7B6LnHqPfiIfocWr6q5GyrCIskqnuHgfHZt
sygEYnc3SM7vmkSvfQBRM3wyPqiH20Tdq8rkTmN+H7m7gdIlJyHjA5n4bntHKC+/nm0HhUpL1NtP
6qM5zRisyHkuY9HEkOSFLsJ3qX8Nz1syDn5RatU7x52zF1bwEv2Ltc38U35jjVVusUKkmi0mT4W+
Qxlu0rCj9XYAOH2IphXt1dLM2b9ImVHoOn7owNmlgAqVzrtPHS4pjZ8yBItgCgJs10owQ7HTV2nJ
DPMt9hEp2HXWGKhyuOpMVz8sLjxya2d8saakqMvNtcHpFEpfjMtoqkYaG4B8P3mMjNVJeU9l7s00
F5B5QY5OigVy0OCcU/5UOqt0QmRkfayu2NupPBSzii/PpnXCjZPuP3gIqU6upwx4hWNVDy0ebTHx
BvLYoCVgHpy8ItgO87X8yiX53GMRKRsb61b5d1gp5XV5MQjMtjmHtJaqnrrQtMEuCv1KnvD8pjV8
2nl7Bfttaf8Q7CzY2LGS4ulyrIbtHhAPuiV+LJT+3FAP0Vc8x5Mx4ToXw2p8ZELFHhvMwkdSLIe9
nuMQZNTlz+qjZ4/yWZOxpiCmmF2601Tdt3dLPow5M2RY/SmJoOormqCvOS9+C964tLsYzbvPlXr1
t2ZBiugnEcBwJVIvynQZFauOaN8ul3eCmmIIUVZ+CCwpdIGAFUwFIj9YTpk9dx4E+S2QEPq43NlH
t4JgX2icFweFCRPKw1TiZwLup3M2jCgFYIgg6BpvvI+yIKcihiQHDRdPJKLCm7oHknbVY/+vO+WT
AWCPVc0EAMfAO7r4iipt/Q4szAbZRFjJc86o0tB9JjM/8UnG13tLopA9woimwENRY9kwODjd7YoB
HpcUd6fzf8dnhMWTHhmV++ReAIEpkGSFgIYgrq3canS0uC6KVQDLvolN7LxJ7icc3+FI57xgxYSL
iqVEOyb2rBXcf/IZ2riUVPAqb7ecOjjagSe7Q3MxH4kqIcRdsTg8uZyqn2xqV/GSq42LfBcQExPS
JYFOAaTJ5TYsQmzJlfgdtUlC8JXH8TteqXrGq5xZ2jXeI9xBAAw26lMSIjv7H6AA4+TZ2aVmVaSs
PQyRSNK2fPcYZLpwFUxL9FvNp81j2p6LXLYeVUFJVkZyGJS5E2mF+6saMGDIBvsTF8wRswn6EAVT
NUYlZqw883Kim8v7LjhttkrbTGvle+g0LO8zxjggtLiNc3vTkXNb7yfJkx6vLua89NNWXgluZQHr
3tqOmnq4N8VjPPHXB3nWRZa9Y8oWb5Szi9RbcaRNwlXOU/US7axlh1ggAHwNI7EntC7QYEFe9Js8
6k9obCLD6nUCZS+xYLxMVMhGSI6DlfS1h0TR9vzB2Aa0QYswH/xpVASG7kAtCTmRukFKeNn+/qcH
nnvqO71dMCJEqJnjV7LGKB0Lm2Qu/m0joL5moWTDtRw9mnL8yFv5SNcEWtH/0mVZ5y363TrH3WUS
8uza403LDlfzpH3SiIwClTx4tVfpyH7h75KUlonWLVndPm0b5EJvyUVynG06yts7k2ivYWz5RYPx
hwGEUho+LwFpXoc/OLlzXj6rOm5DN503c0b7thSBqnRrqYb0DFSxFlTNEBfXMDgu/BNvHWEFNowW
7evD8p1xoDsZ6icx6lhfiJjFCS/v+/t9SP9g3o4S7vJS7+I4Y67Xp5eaC5TC7WspmglK3xTlB77I
efdqwe4YCJjOVM/6bve08qDGPPGgOiKGDRMUWfJcVlP94zvvuWAGzywZFlb4dgNVv+ZLt6nW98Wt
Q7Widwjpfgnloyw73WELoOT/Tsb0vb4rF4uqQ9mY3HtdHiX1B1omV/+i1FmTSSykNkztYi0rABAM
bZwPfx2YE+VBV4R8ypZ8Kz8rpljW4EIi+dzbyW0FMwfCxo3ifDwtW28DCxEsHUnzrQNiiwaItWqY
raDatkXOCqiaTCLYy3ieu84BUBnQWUnN3F5cfSoaMlFqnFOGaAOzW1LuCu3yPl27cyg/9zy6TLta
s59+Wrw2BwEbzD8JzIk2xVYO8oDXOMOf08IpDtwrkeWZr3sh7qEFejwWSqTgge6KA1ZlcMwtbgFn
pE8voG8krqpsyHFcslQ1LuhIhKeHkFiv8BFhMdXeNtneFzO5h30Lleag1FmL4XOT2WjVBW/NE3aw
D1ydI4dVPFki7Jk9wpJ7F4y7ExJ4+3L5kcxXJJNm+tRTxHV4/I5YfjA8YI6Sb5/Y4qTixWt5Du7Y
+IgyOMRAQODWVtV/3ML7XS43fr2PJP+czHqFXkW4gAbhzWwz4mrbj7AMRkVJsLmXI4337pD/25EQ
t8TRgCA/2ihxWfpxO1EEuaPjiwBXKGILQENEl/4lIHw6uHzXIbhWV0raN+LWsIIYaUo+DshAHXvh
9gj1wVzJeSUJNznwseVPSiedUV/mnAfGbJS1CoY2Xv5G6M+ARB4aNalamsmsA4tk+r52My0AC5Mm
Ll6eY1fIdyrc1N/2XSod/A+l88OG5eg/MEVg54nUT4VnGunaffwXKEDYjWXVkTVAlbK13vJDEgQ7
wg55Gk2TyNAwKzMgerwD7V5skKdgThiEZkMnaNLspnmFu+h8Z5qkxILnKisOhD6tYAzX+JmUvlqI
o0/1FOXkol9OxiiX04o3DpkIsN7BJFKzk+VuH7W1I55yKyESc5TVMdt4oKH2B98YSEyOdmTNPTev
hX1wMvxpmXlDW4pE5KBkVzm9laxYB2MtXbUF68RkA/vkCM0oWaJ4gsHwAanr+ueEoPfLjO1eD00/
FvkgAeXy3u6SQmUQpdiW4yx26Xe3dIyy/8qVyyTDHKAdYh4Y+S1v+Wlgg85LnuNiY37PBpYdM3PY
R9nOm7hAvHBTgmLcmkz2wFBVHeWLEHkrE8SsnF9vrJJv83GROJlFhRd1FMQ4bxmdgKjPhdX1Du5l
GNwQebWkf0g6xXlkJhCNz4rXVid2FueUUarOfao3VHMkaBj0d6MtPQ2HKN8xtabLJ+lNG5Ij03QK
ZqyolkCMACSZhG+u79H2ZBABjUirLean2O6/FUNkMCeJt5nyMDUHVq+5224VRk7ZPtgjpfXFfB3m
Ez3z8m4hJwmiGxD3L5zbXCmGw0CbOLnwKFD55TSU1BHwbmo+EzFs1hlyrytxhSa9kYIfCy6DPYuo
uw34N7jEHA/Ipxu8DYwKKkFihjinH0c6Z4c9suvlVeFBhMk4GKvVBc4EgF+cq8GOWLPmK1XvxyD3
7nKzP70xKY1F2Pt2aTk746im8wsuWamXUv8BOuKYTsN1NURPbIYXfdI2AHjXe2AnhOBjcIzIaw6u
D7JkLNcYtNgLTWfQKXIkWOcyB1bRP+3xb6v2kqKjhDCYOFhXXK6sH+Okq2OVVDO2+KbKPLHLUp7C
rFXn8/99fhjFJEtvVhSpLjI1ZeKDRpXOGgt1bqi1dPIA4nlfsm2fLvjCIYJQaTsuHbCakGgPORd/
ehd5lmQbUmUZhcBcXC6A+GqQ5JumWkC82afNrhQNuQrJTld7HI9Y1ZgxjRMu7e1zIjpnLaxpT/I7
h6ej6LJVNaNHNQvP/g1PM5GX7DHGCgp5PoAiToX663hK2uCW1SXCLpX1lyheianLxoyUuql2TsNi
X2wdld20loH7Za5yFhIKNwT10xQKUgdhWZQqGyevXjdV019b+KC6BR6XpsXno6jLEzH2uCPiI7u2
hR/KBWUF+Fago7HWepMlh2muGSu7dl/zVIRzZUb9VoJnexC4jJxmKU0jIlBsE4bewEG2sguZeA6H
Fru9ML6sUldpxiu+0MRJ9wMVcSxBDQ8DS9GN1Jzta8Gmndoh1aomhCMFoMeCiym/LCQo2uV8d2Tk
Oawv4Z68P3E320b73nUq5/zbIm//UYDAomOP9/e327cgeDDoEoHWLltYpTKHfAObD+fmzhcRTDi2
CvqOf+DOPrbxqg/rdQFLepL4Bn8U1bvzPNOxbHimV58AkdFjDVEEr8yuLnRWFVyoVWEJEbxg4QXG
odqmI+159i/xQ/Fey5VWis0lcngw66S52AVI1XEgHIdMNZmbDsTHtXb/49v/2ZmgClCVShzf3xQP
i/WvPP3YmV+1u+L7pG481Oz3g1tyW55O5yH3d2DKeVcqTWPMh52zBaEUNv9FU3YAN66eOJ+2oDXh
rLskriuLATY5tuzhQF17EKeWX8c/K+eTYsklb6/4HSKn32ITv1ZF2QK9xb6YKiNLWHcbgLySlz24
bX6c6tgIdcYJeJrm4UHQD3wY3bTADqKZouCHYKEx/9lVMq9s+ykEvgYyLScZ4/A33uCVHughGlIR
GzEJTLQkHgeddKtg6AYfLVHMGoe8OSSzqnyy60Rw3c+4NZg0pxG5ieUS4lzYftFVgLK9HhlNbozm
+Car9zIAmZVnSWIUCVoLa+wWT6YvSr9EG1hdFJZteeKVC/+BbUYBr8+rKraqqaYWYWCn6+qHQKOm
rssrqY0Vu6RjGCf5d1ZAvFzuYFPjjyX2k9Oe5YvNXkxzTRdUKLNIHj5/1O0rgvQ3jMUZXIBqLMa1
+DRcHMF+wcrHyCksGeNhbkADZQjOIDjB4B4f8p/wWjhkq2+/l9U+eWfbra6mPdvFVZUfF9mv+Y3r
u9Z9UYzoYcdJ2ct24xqZIem7V4ihhtjEzPqr5sipXGlPhS2HlAaFBeYCIPsV6B7rH8fh9IHzfpiQ
u93L8Xj6EgALY1V0vozXrU/TASl1lsMfMe+xSGtxbQ8viEsiHL+NP8apQT2Hiddzsr3bsVSw0c9/
U1ox2Lf7GfDuF+StU7yQB02MOFF/xH1XxD/LNkpYjiNNE/fj3jOPz4bw6kQx6gEICIczxCSj45Jb
uenRxMtP/NQA9Lx10t+xHct9gZSFjGe5cLIjUw5wkZDT8R8gnE0QRyskrMTORci2XIJ2qBMuZYEv
HqznxIWNAdGOGjiUFUdGEa6YGAU5f1Cv6WR603FZx0UWBpJXgWZ2LF3m5tCfMB9ZKHQMh1Pztz5s
9XfpP/iHXsTRKYldeznmRDCSWW+lditQ9Krebff8Vwsf7LAULl42NwT8N1r1oyGXoNqdVmz4DtcP
/EdHLaPthslCXwbe7g1Gd6GdrzJXbA2/KiCuueWgJYssYVZc7ipQ+0lQ35F1eusbhHXtIMlO3FlX
DIljJDufLjM2KxtuCS9wK82ij2P37Exhn5t7Cp7hcWNPGns/zm4p8dGTsBGhCkCu63mNON0jAEYb
LzT9IuIF04DOn9Ecl1fXv+NwT3fPt4Jj2wCkGw1P6bQe2UYob3DRO18ee7c9R4ATRN8i4lnp12xx
v+zuGaG066nQgwhcTnzDFzg4sDS1PVINHXXoPCJTjy2IOgim1RYTbIkTbk/MKodCkbJNBhoiUzab
Yfr7vDeJZBWSpz9sCgppio3sfdVw5vlJ6ZqDN2t9l6R3Qkevmw7n2SMn2B1j9uPSliH+lDzkkzsH
HTFB0hYfssXk4N31GOB8AFPmPnsD4fJiYzYxM6fm+QxSE1tvmC+PJ3fKrS03KWo4jD2O7h7DnNqk
it0uF7OA/TfC4yiMDZT8ncHxbQU0vvVGOsh1P+qOTh2DUho5F0kxtddoUXnaeFBHrfTMpRd57pR3
tzWCPe5w8UjwUEEjoJ4KcBNV13mrPnibmzusTQR8xK78dFeg9MvHIXbMfR3t7lZooVAahu935g3O
kiiotUa2X98IIi6MkT3TeIuzh4wv4sdKJZjrgpsxh1zjBBDL67G5lfOMRc2I6kpS2sz3Du0GUMAM
0Y6WcuhKWecuddcPyB5vlqQpWzMRqqxOkGNMqFXnT2RW5+CaFk8nOuN7KPQu+LrojhSxRNiWodJK
7DgMklVqkfjTKEQMMFOjnvWyYnnOElVE2ESX4pNG3yVeKW95omh16bgtRs06UAXxsN+ei4X3NuOO
UFIuqF+Ynfcx5yzg0SE44J6gCIjai4L5nalQQW9aQTohynRjK3386+pU3chS4JTyhH3PwqWFEqUW
+UvoMKbV6TDIyN0g8E06NLgq3qYVkM26yMWvQQQbOYMw31gRbkxWJIdY3x2eqHFHCHYqEVqa/KVB
OPeo64m30FY8lIJqrd9dAY5xDKvPPnjp5ZvA8PSVZyEd6p6Dts/MBVZv65/wFuP05lKiIhsnt9fO
JeTifGYzJ5X4mlNYQEHzu5I8e6kL5QnUUOtbBIT7fBgwF4p0TaLSgORuwe59+m0TMZOLE15wwpve
QpPBa3NtBNbmTd5EUkfPUHEzUGz6JXqSAavVRCtDVGfwT8l09VWRPp8E1oJPJ5mhI6DrIHbe1Crm
JlMDVN9+Ysnl3jpUM9Rti2nHhWPkGViGRwCOvOOgOkWWvCT2jQUtHQqnqCw9FJx7Ibo9YnuRNdPw
TWAVv0Lg0gaewrVp9JscswQIr5zZcOFpiNAK150uX5vHecmICz+c0dogrKbD4LH7fEE7sz1iAQox
arsjnYzUVaVQTr4Gycrt8mcm3X44sAw65HF6x41W/Y0HQTNnBhBRMrnfE8qPXGypk3tW8hxxgK/7
CSFVg8oHzeyfM/FqM2saT9oBH8lQ36cgAxzEgiTvniUt0Ho3I505jFg96NwXceSrLD9wUGYQk2aT
TTMa8SVxMw1W/UacMHa2C7tkfuqHiQkurSzD6CTuIJfC77jD+KsKRXQ6ZvF42TNvUYXpQWGe5MGE
KXd07/ogLdnh330hoOrFDzxqune71yeTObAuuCD28EL5qFkB7mr2b/af0VWSsA1pYtGqC4AuMuA1
eCVwmZNDTueg/IQIm5OURvZVZN8TiGw5H/rb4fmU052b4hvGNTaYPhVZJGHhSZGAuGsOF6ynWz9M
3nVbPrTd+/W+jAQ10D35ZStsImKmVN58LTo40p7xOeacBPzIHJoScm2CjcgJil5b4UMFelC7Pn5M
ilMnZGkz4AZqSLET9+m4Ws+4qU+Z30nGbgXV/Zb/obGs/4oolIP/AYs6eeE2O9e1IYD1zfXkWbDb
uiSca7Pudj/WLzrfGxWlhRnn9HqHUGqNQxVPrHQCFfQOKHlyM2HzWcAhONAj7Uf0VfI0Rfu/1e+P
kXSykFern8eiZJ2GtG+VyG1B/qP2tFFAcUtfqumD+Tk7TPD3YZAzXZ0pNGsn3v5a0qgC6PtVwc17
L/nug0LhT6r6Vley5KyGiAQZVQVvGJNaUSFR5oapiaxgWhLGuYj/+Ifm17Akw2/4Gv4nmwoQlHis
8SKNnn57Z/DvPFc2XVRAMK5TJBj2ZzT+Eyzp4o9k5jsu+e3d2GpAG32X3PeAvlkX7VuD9yd6CNr7
6NUiFrrppFdecN3WE1DQOznbjm7blwz8g8omdQ3KlnZ9gVPz3Nb4LSyA6YEU/0yJx6ycWMoi0iPZ
AQXIUPNt3PF5aRMhWcBeaM7qbUUUdvynI41UfHZ/+zf1COkAy5mNWfFdip0wUPHePt1OCJOR7t/e
msnDGps9ODBqjLuCa8Kditc9X/G9AebnAMtyc+EqhY/OeBIYNDFIQQ2XLKejO2IRdVuBBr5LtcgU
5GQi1WihVnap9t7A5odon0yuG8nG/SEZWm3GPQrzyYPKb3/oNcNtvq/Q69DZ8WYojUpWiUHnvWeE
Wt3M11Zcaq3ND3WhlI5UMcsBJ5uudMSu6DUTv9XTDLLJDlFYLTi7EzW+TKRs366dmsFLrb+wDNoY
kfm2ycblcc6nZjY94bEKEibOQlHY+CrnhCGrvWD+BJtdTMiPWTowcq4jpuns4JwktXcTA7vrpyx9
LWqfwGwFZg7MlN+aOJ1zGz50s0K9EdEWUlOqrPgI85DihfMlkUQ8QlU8JhUqAQH+qxaFrRkfd5yu
wVzdLAoyqNEqbGPsd/G3fz5cXUHOoM4uxtMxhMU1RyuAf6+j9NXck0yBmobZkkU8Gl+j+KSHMCvN
pcoPNUffkqSXFNJ/8MLnQx1AWqT+Kqv1pYMAKvmVosJCFv3p0gFQLT8lgVWRL7LgKPH1bgROBqFf
48PBfqwi4pW8SDCzddAGyQTY6RgnkSVKx2hlA9pAWSZpAfjh8s3DVl3W1qob/eqXz6a82pVeoYfe
xf/LORzSTNyzoYfgqkVheVUfosYjPu7y+1ayNTnA8+zoh+k8O9KG8mI93G4elPvYWVL8U2HqHEki
2huMga0wKU9M1/1yPp2pOa0hWp7LiIq0F2jPkPUi3mBT7V8IdlcC8Pak+UI6INpAtPFrqlYXa5kR
G8bIw7QBAYTdneKjTtSGXuAwE8/GBiIwEEJcALyxG58nu3k6n2iaVvaJyuG1F4Q5aBKvVcPi+FGZ
EzvnwyD/73pv81OBx1GQXoxxgysPLJwmCJyVhQog56drBTOHg/hYZcDPXq9+FcQYGBupij7sHUMf
Rv9Wofwca7SemLr85SsE10QKdHL+cNs4SwHOULBOZL7x92Ohz5oP0HzpbKcy7XUi5NZRmS7LLCpJ
AjOE+2qIjr1Vp2xfeb0dJLD+3N4Gy+XhKR/617Ml/AIc8CNAnIOc0S+E9lPIsrRD2VTbmiVkAnRU
EhKbv8SaXHIuzA+hfWvSUj5kdTM+8WFmwmBUg+3qP4BFi3v3xx2WXNNhWF8LYMHUHfyFUmlVuWWR
aelFjMIKyMYo/Ru6m4zNrRPkL+QNRsyLY/nhtOSCNRH/2xxrrpqC4zpkOad+f9GdcCfcWC02SqYw
7R4FZhEjfqoXh7MTIVnj8f8xDmkWmmLzDHbY4UDcBzj6Gwx4Nke8qOqqcWNGXa0xH7m96L5t3oEe
ltXwUq8WR0BCNBVVjIttMy3GYLYthAcXZzHBTac7WyXRawraWJY4Exzk5Cz/Fib81If+O7rfTcSr
jiXxRpXR+GWhLjHB2IvsUR3OvDEgoMXTZCM9PhPojsoJJqqXePj0k+o8AUa1aIDyYPOsg9XmMHUK
f9TgSL8JxG5P4di/XJ9RyEAYC6cluyVzO+kkoE0/8jDNLWfJoX+UZtplZkUGYpB4Pbuhtqw8UA86
J6DB2ihoB05gnA9M/MWa8bJdd8fJGYyAKWPRMSuYA+z+2viL1JcEfGuar61ONJ8mVnm6i8/jNCNL
4spX6Id6F3avC3ySMgOwAQ8itbvPTIH6IrNjUeEHk4NH7XF6ydAswgoNRAClwvqe88ii7zXQGrJZ
V7sexWuOwc5GQUDCMAMAGowAnMrZKoFBse5t+/trx98z5yOBqD6HAcLX0ao4MbDf63BE55RvWMBg
wxH3Am1qAg4YrLKraPSLIobmXgCEY3xRTcZW0ubTIZPoMfNVSWYSQF4gEKmpeGKqG8clBUDoBJUi
IxRr4MhmV0faM+RFRaVA6pUvYWAhgdTwPuXLD8SOw+Hc/6wHd5L7P0QagZqyvj+GDoDU7CBDZMzg
4CAMAH7/el7ihuyV4BPDfjF+ERbagkHab0zS1KKl9cHUO9Xj74n64ZIDiL3AjH9z3pnKT5w2Ct/m
tZbHYPQ1255c2fBaIhqWe3yHegTYEM2TVrLfznvh+qlv8aypU4GhZmM4uY8V2jGbiKgutdzeJ+4N
5oqcbLGGduc3gSNduZ9kBYmjkDVn2H1inFhZc7axmPqhRk+yiBYpotdxhNSyqTmJqhdbNJ3zrdWy
3bIO1JEeqRtfW1jqGKJX31hHOJpMTF9vGywmuFuu/yr+D5DmVC+7P9i3KZHmcfiOVkO2st4PQtGv
QPiajiQm3p7N8JnN8o3P1LYYWAlGSO/RD8Y7NaMgEHi/SZSPwEwz+t3GAnYuMN9RGIis0sqqh2r8
YJ4t6bCQwz1GHjQqBa6J14+tBOK59Y+T4/pER3EVfHnt/8BGoBXyM3+eOvyjv+3KU3RceeONuYyM
OSjmd/TZRqnoUwXHf1SVlgMFmnx4m0G94Fl6jKQp0O/06SDIerKEpiNhmVFCMaTa6zyagUoREqpH
Qedx2yu6GeCmI5hcjBzIr7i/DJbzOQusSKlCSA0MDLcnOjpfJxlonj2DM+fjRPNGKSrLDpr6bqs9
n6M9H0Qh0tm7VSS/DzHpnelu49w2NKYWIwa4U+hSKJ96iV1Ffz9mYfMgO6rYQqxXKHxHgpsXIAu3
XM8PfKcitOXzCC0iNWezrFFh67LcjNQg1VEST8nJB5bNtPrNYABQeXEQv/zwcqLDA7dG3tCRIleu
579An07rxN1cWzMy+MMzTv7tq5QHLJuiTCC0xX0+UvLSExFY700LTvuaGT4PNgW1ALAMJYA+m/P9
AROLhohK6EMrCuJB+e/JH9ZGwJb09w9t0L3pfsDeMyCMUg4v4tgPGkxBpSmCJDz/dsUXlzPrtXo7
1PtLbDI9kQUKpAQcdtDZRWmJ8/2pil3Zk97ZWK72z6SQMpLcNOvShKUFvm8qrfPT4ZayqiG1vodH
4kTsp4CCkK/7SvYXykHxL/ppZBvhWse+kX9k2wnuQyPukbX+d8NkmjBBRocjeqKgovdGYCqaKeOz
bRwQckmO4qaCqThxJSwEKgki1vQLsicj4DoAkBfnZwXdxweYtyu20r7lsD4iOSDO/ckxr1yNEsMV
+tSwFcf4SoEcC9H0WDNp3Edqb7h18BHGdA7VWV9eaHuwbWow5WxKXgzLr70/egC4AFCCWI9RTIFn
zzsuiNFap5S5un5mcN4Hnj1NQW436OUmG9V7KDh2jnBrT6C6sZBRMTpv7imzhkNyWbjgwJKthRyn
JZ3GPGfkbafYcecXauMDHGY1CMnJHEv06ohmzLLn0eCrFyn8dhSj9Io8L+0MKSsFv3AuyOJqdeYG
c19N0m8so48Hv/NGqN1VXZLpKwzlxvZ7z5ETlqVsjOsDp4lRt9CdOde0rocNT8YG3xhYFt0HL5kh
bXdpetbJGcJI5TwUFQZHfXMKzKHpCxJmeKCk/890+JEml/hNGg49U1LmPvQDwaMRcr1xEwEZPzn0
TI8OMdRvoNbGpAO4M4tJEBwsjdzr44iyhLAyh5AIKUnvMvlAzYZSJApFSPY4PyJt/pO95SKjY5SP
rgYnDyue5EO8uc+wTHpjA8laEBUVszN3F+K73KAhiL1mX5SXCspYlQoKuTfKUhjsGGdouZd+nZdB
XRGD9+PQvj6tpOyb1gofGl2/lwOvNyis2fCoUeMhb3Icy+cGHGF5lAI4F+vAin5xIEuEBvNWN7Bj
GBzyNuUsKlnG5lZR4OXIC9Zq4Psl3f8/64o9LHVyVz/cIKVXXy7sWW1evvTlQiHMy5XoZp2qd5NE
uwRT89FhgQyNsvj+AngRmCBmJqgAFWd3P8AhuutYiymK3WkF2anYbKhEI3sSWknV75xTySreqnXc
r9asTR8WQHErrO86USUKRaBGqEtgL+FxtUrC5RkyJHAIaY0BjNHxppntdWPN9msUq0qkS2W8FuDg
YHPINsGeeA3N/Mnf3q5t2+r4HZu8NdeGcAq8IKvsDlbsM9ROwcycqe5y0wT7QgyaTWDPatTj1qmI
GOE97tiBNlIrFP80TrruVkTkkpv71BOpSt0ZUi1KGhpBPQB3ZyqC+z3u/zXDt0NkovxLfvwsoDa6
QqGl1teBrGeF+GqpmOT5Ndmm382LGyqXaTCaR10QmuTGmThv39pGMwjBi2CZUESjj8elPb7tUGVN
IyyVwYd1h4whlr2EfOjOcm47Swtj/bs+C+FW98zkF7XJR6b6SKpafYF99PIoMtxoTmmgPO+5kDK4
WCdY/jO9hNxdyNf0r6uw9bK+8859t8BjePWgC9WrKN1OEHgzA6Q/7AkSIudbK/1krDUTHTBhMxsF
pItiT25U+Zodlb2FWU3GOLIXQ/2twD8hiWfdALFZXl3f/GKMvZ/K/y8rsn61X4xc+Gcho8Rdhb43
LlmkBKROaskOScIlTxIYtNAn0DtK6IMn7o+dl0u5u4+vQbvEHypypY+eKmNBQwrwz46mmjBm5Wn/
WNKr42wDS7oEnnfl45KST4lQah6lkxUuQYzVJJH/+TQEo7lXaZ47vgVhvgaX9LsGW8JEcYlM6hIg
VqcXF5RdXe0vA8IZWW72VoToa9R7iSSwf00o7uQSiJmFtgV+a3eLLmFtgUuiSWNOO/aZkjZxw4iE
y+/dhYjl6QK0YdrMirj3avQ/k2pwkd1FTuji7v2xnvgb6Am1IUS6VUAbHJrZTyjQi5cST+yh8ox8
gEcrB5pg/djbuByafuKkljynwlMUthbHJYSXFQHKVAg6Mp6XEBgp2s4xEmgQSdlwWpaiSfZlYS4a
R4mdgPmCBrfixL4C/A+sr4fMc4rw8cpiKbGXQz/GWAHHZ2T1dk90ypYIjdw8RXlLJQ087PHETo0C
YV45Sunwr+vXXIc/c+UzjxPczaiOcpDbBtU3affy3QoSeYYfbwE1//4UaOwKJcguy7gCyr8972Ta
vxTVWtPJtP5IGVhYrLCUCmui9NR+WNDl0ITmQwDdOSpl5Uubq5lHrYApn/GFW+ZseJ4WRHlaRINo
ma5CZ0j/O38xm7uDTXRJPxeNZjdC3jQKPVr+0C8YTcNa0lqkSb/5fM6WvGs+9ay5nyKGxEd5qa5l
bOWGLMTVWvJP+TigrFXo1wCw0Fz0LXPzQimJ6tuyqVpnXzRFUpnyuJ0b7LqHRsizGVs1o5helhCF
sUt8bj7+YEigTOfKXosrE0j3iADzNxqaI2F+N7hdryoRionL90tb6i8TLMdAKU8WiQ6/yhux7wcT
hDOjdrtKDEauG6RGBVN9q72CrCmEaB17jXUsfnzkB+Ts7FH/ZcZQzn9Ams/XxIyJwBmi64zBviZZ
UUexfwuUxtOk+fZVpS1S7Z06mPm/iIc8Hen2tBBAxnDW0susQvutBRxbnxifk0OUR7GFGF3Qyrl+
jK55ANn4pIn89CmaqMti0jKee8CPVkufG628o0JjDlqZxFuyffUYHREaixuw+IcoJL7S09Ec8doj
XYmtfEZbjLKp9P8tNv7k0jQZ2kEFU8XxjjOIXZH91Zg6lKrUxgxXVcrxOZCt2MJn9tWvYC/IZJEo
R/HBBPy7rFcVcJRkmp6MyYqrIL/d/PmqdLAzI601CXJyoPwuBCc2csOtVv9H7K/xZG+LA0otIm89
nEOI+OHt+624CFWUcVX6/V1jsAZM4mWhfEFkCXZSPTMe3iX1wdQl0eVjmhsAKKxAwiQkB3hQ4tGM
NH7Fh9kODoCKU492A7KoTevR3fO5paSKhIJQWp4hj/qh9Hed4VsqVRKjlDcGKNaPNkwMo8xzRvFR
ThdMnGxNU8P7wIF4MzVg7Yik1jCYhJnb8iNd6ctvzy2A1GVhy/RnAuQ6HgcwNeNboxh2cnRx5oev
AxKsYDrQJAlv8XfRXvYIPetU3KlHMf9I1dLvCLL6/VyShvaFS3TDF+CvdIuCROmHd52LTdVXm+Xj
Phw1yHlt++r3vdFb1Xz3m7R3Zy/rNRyW6rZZjqQXDVlCdlG1buWaoG/mLD5MFpgufUur+VpObs1s
aZjByZjpvL6OCFZAyJiwtwsnImzG6Rg6MUYcy45egez18KWbZVWzI/aZBOP721D3ihYlCLxVcYEL
dcQ5TUxQZV4iaoGCy1sHWkZrKFKsFJ33bnxfGHBZjzwPnxiXDwxveri6Re7u+ru5gnI0jNuNOHSc
V0rldRz+eAMZ8v8/A4qmxI5clZ11ZgHqs4G9blwX4h7IFFIQ6Bo6LBi2akGOJBStuC2wcf0nwIFA
5K0OcvzxJ3BXZz1jN9hXJ3VMgVXdkfAsGr0IZSGEuCqXRi286on9aY0uHhn+Xm86QuS6NuytIuH1
fZyVD6PKtQfHMfWNqSiAATiVMPzGBc+LbW51HXooXVIulaOrFVlkcOD75huF8b6tRXltpsvhGhri
uNLbBY1EeeSDVvQTZFmSJeAe9ICyvpTQ1Oa3qqKv2fM406y66NRVAaqMRjeOOZ+gLDoeRiJvafKg
aSfr71vuAkc92NOnU13qykedSbTDbsIti4uHCxo//aR96N7RA1P/7ULhDp/DHv6iCNFrgXw8rt2e
b3wXEuh0oc34bYSReBH9uKOBRvtIZzV8qQcJS5J6jDfvOShsJleg69pUVqFjycn5suUVInIJrSTY
CnM4QC/ZPvDHgSHu3y00tVBToXLmCZDfCuCzNWlog2DQgxgUg1erJTELhnC/i72t/74Qzn+EcyKq
LBpYbUcv5iZX+vJWcFmU4kFgRPz6BBv2xeEfqpYbuPhLOIZxu2pJMCchgmSRuWtLZeKosFGBC5cD
0pJRsN1C7KF3cQtJbP/wZcwNFdKbxudv4ATpjNnxv18pDpUhosw4paEL+SvTEl/bq++Sbl+H8kMG
lyLyIra6Iq3RAsVXC9+7QSNlGHIroNf2M5BvMZewlrnD/6kBAfwiswZL/o8rX7r7TTYNLvsJH9M0
eowRvlhTk9DFexBd6P6/Te9a5k/tmwlVluhoGPSquut7q4xRpnA6KsfePOJ0qZG7aK3YIWPTniaN
dnXemskp18+UFW3WwlnH/cNyUMGJ/o0O8LMU+tYzRVEpzjtes68EUwCKDT7DxpZ/xEnFV8X36Rpm
bXqcmP1GX6BSZEOVzc86J2Lott9Dw2uauxsbD4RdjHv/Pie3d/X3LA9+kXFLsBFnw9Zi7td7qxMq
JNdX5FDvmfQTS3kugQaKEpX9Lqge0K1lxuG8O3XNbR9LseOFgobiUDWMvv2OfkW9s+P5FmDMWeP6
npDMpFugOKBqu91wrE4sHh45wB0r638XXmdkw6Ux/LVafHcHEtAelwWn9f/v2Ls9uqqyuDLVUPDI
pnFkMwDhZUKCrfwc9mCMRT3jLfgrDZDyQraFUpo+IKYifjcQYymvsClpf0KEmXvS8Cw98ymvPesT
lf1Um6QQ/eH8fzVqsGrHdNg4qF2OCV7gDk0LpKaa9o513qD4FN3+krTa592784Qr0p4jzr2g80xP
l4CSqh2QORpbuR4JE1u0CEHzpzmCbW6XcekPl1McEWE9S19W7MbxYRAJv5Bkwy2KesM2MFDG2jgQ
ovLQW9MV3pOkHC3Cbr8v9Zer8yvTo0yjdt2ckbUWZkIx9pb4LfYIBDJWIrbaRu6FJg5Ib/qJWohM
x6EN9oV5QsbbXDL3QEgQ4221dtRXFhRSc1SXBiRSWNIO/zIuNl+fjB/M5m9n+rQEzEVA6XRSAC+4
ZnCtjyElyDl46dFWQVlT84z3dxHZ0LOaipwHDFeVSmeHwzwCVWFYo96EoEyaHnzwFPXWi40Kopie
uktCnnnmqFbh7g3gQa2KAjPPVrh+kQp0el07y0ibyzdfudzeJuS+GaYL8MWhZ0Og5D79ayhya1HD
WA4YnJkr7VSC4wBcJS4ZYp25OUbrxl55Ojj21tP2xJqP3bWzmMHtXRQgPpistr7dBYUol2MBOOa1
fUBtgv5Z4EUhtGW2p7LtWDw91by21eZOiOwo7xSAFLQvTme0vGEUvL5YRDr80ggjz+V/20NsabXQ
DIP8UeQGa6JobdnihkxObxfwm7GTW4HOxDWwt2qbbKcT9Bpz5vuqF4VkWhgT0zcSWzC5oxqiaLyj
hGuYPQhROimwyYTMrSXuUDNlfeiA1zWDshTsg9G7G4zmlE11YhXqynQ44RMyQjbW8rEPDLKgdu98
qg57gb1rpl3etujvNoYIkeEdah8c+rsMrdd4DjB57wIc+OG6BDK395ulmqGdlQ0+WE+EjTo9KzT/
zE8mKzJ2FpZ27eq7c4w5CcVX2OZUDuLkQmbPbt1saOF/DcfSgQ+QZnw1dH7dajFe32grhlPWOd+5
9ATdTrmpLaOfCHpgC4BOhCLdUC3xzhqwXfuB0Aei/yGQYNJPX30XaBD0ON70ueuyQ3647tH1tR22
ud54cnLtra1rNZ5uMT3UGPS6h2YWn+1+YKwdQ1zPC1vP0K8lm+z+RUZWaM8xEiyJIROIwj+L0Y4Z
iYhrTk7/bOseeUOZjcg24Z+bBqETpbDil5DtPXcnVgcUpNOSX/PQ+nkzq92i9MwmRl9Ze/94/QB4
5orfCRHuLlUgKq3+zkB1efiMh7AE8o3E0uVTuQwwtN6KgdJOEJ3GWohy+UbgDjGObv2n47PbPOkp
SaWgBfUlrf/Vu1E5VgJzMdNzV9lZCKh8dROG7f05KV2zFnmTDJ+/B1/kWlsGx064Ju8urge/b75d
lBI58NV3FB7A8E35/3d2rrO+Sdk+LPfoPh2fYn+ZWLGRgc1D7E3V493F6sck5v6+JeWUkeSag+Ld
zADnD/e5ig/gstcTKW+z8fRPsHWFA2nqUGuFb5iHR/Hq1ALcmxc5lkHnPk+Zg/3WjZqY0XakvKws
9jNmH4NECv/kW38TgH38Rr1/2tU7vcuM+B6TAfD7slHNNQQ7XeN0Uu3g4GapWTFmtibLTU0UeD4K
JbqsVqxY3TSTB1IGTvew7v5S/9I3ingVfppP7v2KG88rFV4oFDmRq0W1u4srSa/rh0Io7ndp8NL7
LrpxcizA1dstGwchprmFmPOqh1DSA5GFwYfroCBlP4aQAlHBGMWQ2I94JF9N/fXgDT1vYJUxME60
7omVzTHbMAGB1GSaNPIQr0Ho0IDayZV6cRMtGVbEvqeczq+3MeKJQJ04V7iETxJesDarf44qIHX1
WFU10VqCn/XK1DxwQU0WEtGky82gGfE89hS3NApzjog4xwaiNXks9vRARFg/HuOGuGOiqda3xn4N
RDnNSNBnkTJfjc09EHoOnNMsoidpE8VPcxAisaIRiRzavV0E3axrJ8g+jiEAuj9xHmGcmmM6ROcv
P7pxRDTfs+krsKy7qDNCs32OUN59NP+YnuCrqvbSrU9joqpsFKY7dLUgmAWtt1dI6+G02fN+zB87
U3Rpc4d1owov01g52u2aCJiVEOH6P8SVb9Xjiww2tNjY7xsJhh16iLPm5OYmrvOimieIcSXjoK1U
MW+WhvPnI41FypHj/tV8tGej160DBc3lYuNZ8ZrF0kV9pc9wJDCMBRYybqD7JU3tcThjvMoj5atJ
DeMoULhwil9tkfZlQrV4XTk35PUK1R3BO8KnOymLwZhoU0Lugsu/fScn1bQvsXRfPLXVc+iGbJRZ
DgWZI4X1YjDd8L7uocpuu2KTaiHL0ewnOvhHCeCWckHQEPPR1a2O9izqUBj2vtT/zOFYpnDQQgVQ
ZA0y0DCOOCFlaLWSbrFloTp5jHsb+PoChM6+Nj3T3icN9pB5Ddy9QM3UYWs3M7USk+dSSZgi5EVf
pJ2AyeWyzQGgcZd9lkH9RrwQEToJxPwXO8qnrNQV8+t4GIYEsWAdlK0ccwea3C4j9wJuGjouH+7A
fnAvx9mJV+g8xqVMR66WxzkY45TYKm0XgbvmbemCtGyRKnAJo6iq+y/3SDYtUJxRiR/x+t3VML+g
cBPY4wJ47tpuDYYM+FMrfcEoTIH9KGtWBp1zJVa8LTwDsi3u0qAjxD3qYPL8vgx5knJVSZS001JU
at7wvignDZdV/IgwfLxOL10Q52P1Ns1QZ9GvY3AOVUQp7s3Fmrh1t6Zr8en0Lctu0C+cKeZYQGPy
syfkxFkIW1Z8adcYKh8XZsftllNUTS05J02BYoLXgVaMK7XgV63aCAXATMNEDfqiYKlr5TtQ9MPe
H2cF2AYS2gTC1EhIsJ0HIxPAvFYNTwHF+25LUXKgClvXEA6kYDJ04j9Ebhq/J/+VXTw1BzrNgBDU
lBc15mdHxWjDcnVBciFS/M+5I9T3mt2ReiZVLg7T6EDT80pc7AZHxfERS69/zaYHozb3yW6vyv6C
SA/gA+Pk83HqgfLd9jqCTSWaZb4UFM5pJMFgzy+9N96pgGl9ovIc1E+VgQGe52EYn3bS/GxUDz7o
olT0tN/lR5VHHGgXozFsk/w7ycOxJJk68AN6OviOPkztSHBdvJbneqGegC4eGqr5+7UZd1LeU5LE
QLbWCl/oQWhkTpUT766Iufph/PJqOpFjzmdWIvXjktcLOX3I5+8XIOUHB35fVACzCYF28zDGOiGq
JOi10az/MV3Kt+PbL+EUiDAQdG9HNtUR40RRXRJRkupKMNqF4j6bLx6outG9++z5naJP4QKi6cW0
nPkx0Erko4cm4+8BNYI6+XCpsr7uaDWFsnmZDFkpm2KH5h1AB+EiBDjtWJUxH2W6iWFss1xgDPAU
d+bkPFZV39+nbNMNjNDbln9X7cYTw9vC1L7dvoqVRZTr2m0EY/oE7CiIPp6B9zDFF2fcWxlCqn6u
RWcpgQFO5PPgEFxcYpMCvSWGg5+fJwcwqJ8R694Ddn5WvgOwFyv0dn/WF1cmUUGTRsrCx1HkD0HG
2MvlcctUb9RwUP6V6EUjtcQW3sxt7Q5ejiTZyN1ZZc3M+cCN9HDR62HRljeEDa+erEHIjaG7n23G
WvK/LMFhdhrWlXIWYxCS+Wi83Fp3yuRsXZf1Gd8aPwFXmjSGJHINoQ/9L9mzQCXhue+MxiKxMKsJ
3heW60gCDudayNBpk492Jg5T7ZGJ12h043kXsXx9hwm0vx3v7R6PmezgFRJqgCiI36g44IKPde8/
fShuLAVOMvQiv1HvnMYqxMEAiloygnIzrCm+jaDgpBxV6rqbeCAR+ucTRSoJCBt3JK6Zfs0JnLQ+
ZJFJM3fKxw8orTpS0N8qg8zLIbP2yqDIoJpfMzjSp87+ci07pRDoofkIoJmKM0FkzuIb49Tjk45N
KcGt6+zqUQkbMnIMkjuCLmPQOXtgECVz9hXHDUQoErMz0WRN1PijsWDqnSHQSHwhAhs+50X40Xw8
RVjTDNNF9MJBeYXAJvPjAxjAUsXm/yWESpHzMnsb4UO+UA7UTPW2aqbtf210YDezxc11ptm8H7Zw
hPCwlR0PR1+QetMv2LNmA/71X2CtLmLQ+NdWcA7IMqgovhE13BBjxvMdBKzwNtW68Uw+05oSFvJW
9cmYQJORN0ps2tqTjU948hhiuCECRz0qSNypKM4C9zOgUTAxOtentme64RdUnl6JUElmp4iBO20n
2nWVDd/7teBKGR9t6xvPxOCd2Y9gjIEIPnWfIBciOHuKmKfRCuzeYEdQmNDtCvVr6Pw1TvH+dGKO
Se7kQd+uN2v8eyHCMoO+vpWRxs05o4yKsdwfokMIsChqcQNMY0XXWaaDO+9UL+fmmgCTaMZpn8qk
pZMlE6yJhh3olhTzXNIdjBmd09nTs0L/DNAhaBEV1QYUtZrJ3vjqn1E9YVy+wOytsmM1uy3s6ee6
3NKTYkUtopL9fHOWg7q62c0Cph0vFUfIzDkcbutONCC//ox5ksv4AmNkr/h4rLIJvxUMm3eY8Yiv
5RO7OmRYopsnSXFdK54pQdR+j3/bPsyi9dGfufpn6Y8DotfgJzt+aOtXutasUa+g/2+/EcZ1cWvw
9LRikFtb2FKKfz4uKY4D3ghY/WWZ2dflVFMSGizss7lF62GnpACjn9+0Ba+l1lKEPbT9+nxlzByM
oxo7yRDwFdG1dclc/FPKttHs/wDuFzIdO5IRfFfEG9JDq2tzjd04kfEwpQgP/Y0KhOgCVWOraSQN
+iL0kD3nRS8U22leBjRRJIQwuy43EIuvoQTGvkgN9ESl69VvxjOXq9Fm+zDemYUlbvJBYzjYnxHE
VmG7LiywAZj+L4M5lteT+6SzA8BGS1zV/9Vd6nk48AkUDNa+BYOUMLFbn+3g6ugjJgHL4Tsm2Ihx
M9U56Vuq/C+3uyCdJm24XaeEZvG9IBDEIDMgMKV70Xdz7tdFYsK72VdmHz9KUykvdy3D1FdKzhMb
TLdLYVCE15Rhf0/fGHj9WXTFuNbmYUMzTaJaHikDGOa0rDVh1sr94B0sphi9KTCpdfFpaNMEkst7
Dz/9upKupaZ02jd2ocduy8puxU9YsEPE4l30FXAYh4sH1V2MKrR96Rzn7ogL3QZSJ9wjJgu/hNpa
DxZB09ERufBS6nwm8/n8EDa9MrzCUkDpsjHZDr2NooY50y5RNlB/qvcmt/7WRfXMPz0l6wLN7KTm
hdVBCsjCM5XQnnKUuPrgaD7qE6mpi+dy13NH8HH90Y8Oarv7pEZl5TvpjOraesfli/33BlA87JsO
P87Hzfh0QYeX/xVP3AdnvQw+iPgCSNt66MDi0PvcIyaciAkTFEBEhNIp4AiEOE62oPaL/Rkh7dlU
RBfWhvrKHS5YR61wdnwB3+IEbKNHLieu6IygP/tZ2xvUPn/UfDnROG89WeXdNYrrL9v8sv6Ubvvq
MVpTbV83ZzE8Qcku3wwEkp+D/qEyyILHcwIEpPO5fsLLKKWd0ZRbU+k8n/15v1pY7S8vE0w63kDD
Mc5SsOoRWTlTzZ4nsj+3jmoP6/wAukEpTRyORRWPExt5O0RJfnYaOJwINpTdrPQzDMVwWlh7jivb
KFwN8lhqEkvqn3h0USExbEKf0elHhpA7iyKLV2LnS/6GotYlONAVQhYxO4b4Nro4KjFmnvTw+0a4
e8mRxrKQfH+tl3cMHMRIIz1PMt6rqmlp0aKN4XRTqX07CT8yXf4MLGh5W8HTRIV+3YijzjBQZRHo
6xVJMCcaxbJUR5/OVhrFoEFMZVBNqsLhLT0A2TWg6LOKxPlLxWeBF54BQ1+LnYj1culVXzViXsgy
hhwbDTC6He238ObYAM3EzQolPYmKzUQzpcUGSYL6rANKSEYe6HYG98pZNPVuc1IS7A7rj7EV52fG
Yrc/0x13wCnDYjqlb2bTko40mOUGJJ4UP+OcTW226VitCiT+6GkQLw7tLQRo6jyc2FgD8aCqEDnB
hufvIKZkYMDshMUMjQnNfvoCwF7mirTORmRQfv2F7nrlL9J1XvYdPjw9SSiEUp3AptcqBndIegGl
L5w7PnGwqXTNLUW9vi3hwLpN32lJWZqBkpNNJTOBGnkn2LuRSSqKMHID3Kme4r1ux6vQcw/2G+nx
ZOiQ1kl20NVWyPHAjw7jlq+TEAerofLim53H9VreQAQ4HRnj0POehNns14QgyKNzXrhCBzBq0PAN
+bxNBYG4MP6R4/fVTLJk4tAYnyf+Y6jU0IIyBEpyf9yZn2N2DMUGjR/7nf7apJF1dbDpMjdJbazN
ZAabOZxNH/28+7073SxPF36Nw++MU86tJ6W5VdsuJPayMPmCPYZ/yhwrmppfEc0BoWeup8PkCOuV
swA0bE7rjJzByrZBvk2tzsUzq30u8puY9dgH9NGG9ETZuVrTB9f82WnDsyp/lgMyCgUwg2d90WVc
aH44MIeTfHEa/ihtnu3Ncl2RCzKgqFl89IpkdibpMzdOHCbQUjbWrctb7qxnifHKdftIdPJtdtJk
ixoVf6CFXDt2mU5loxsfBXcIB8QSeVQ+GoKVu3VMy/7Z582essnNanJBXJVTIDJf5JobiQSIMbNC
U5TJbJsXlXSTXaJT/DOohIFkTBBd9GA1ZwzQ83B5jk/CtQgZfAo8VEBAwQNj0m9J8RlhqNtkRS7J
EY9YPYdc02HreKBEVamm6Kv9CS4PxFa3jFZDAfNP4RoGDAkyfRXhSQjd9lQtq3vagqee3tT9ztns
fylHYykiDjAOY8fq7iyLEX7U1MMY7gFE3c3n8o5Ffiz4Yc3Q59v/nrFRsQM7F/K4uLO3iY/y8mzz
BE2seg3xzb//G1WDyVk/mbJSmPvLgAzywzQ9/qrAAFXOIrqBV2YehjeF6/ejJFRoN8FPBtbQXeKb
K/swsKP2ez1IEng9l183pCPQotbMQNFYVwb7EMvpzxdIDenSclnLPqXXwbyp9jgtagSZg1edtejg
c6jkxt9e9nRl6MCPNk4LjJJKxnSHsyhIfnG94nLnaxWCP1Kc/06Fqzvlr1SystMIToqthWcBOWyh
XIDcy7ZpyJiimAhwkeJTfixOA+VNiLdoJAyVinF6p6Rp3iA1RUgULZk32dJc1gBika8ajWT1w67B
qPxpMJN/PezumR2wSMloyQmJtkYv14g3I/MsKa9435MLCg1pPw8Py2yMY7A70S7Ozg/kutJe13S2
9Alk/4kX7T+RbIV6Yr67GwjUYvEh/gHhpdm/XkebchOYkEctfpIdedo+8c8LWxtKhZR84Kin+94T
h5Ji3Hy6OYUts6ssh6oN9ocGBHeyVLiVMSaV6gPGN6bp4wM47x2RVTG/4e2m84Kb0q2zk6/nYCwO
JttG78c+mpdGSW2ilZD0OFS7xrlK4x87EdxYPe1JQza+2U6e4FefQzhYIw0q0pmxlSjy4cjlcJsv
CrtCkKIAaue+ltvAc+JaYPwQtJrkAgOBpX4wC3V49vqunFCIwKGccSHWh2yk8V3CBBGT/3+ccGdV
LSlTirinz9bHVDDA/vA2smIlTG+/sJlru5mj3QXOkLRKLuWCCejCq9yrW+PRXPSE6zjM9vc6STKG
NcSoSvhloBpYPl00MiXcZZuHIoeyHN8UlSKTpvMnccGu92vfPoSbwM0teMtBu0xZXKmkoGJeUIIm
WqRb01dMnsLXN9RHjts/K3ZvEQzxng75jvV9ISU8tczopsRpCtygXQLZg+XatTU/GwcsexlTayNq
/mq+heX4VisdkOPQs47RdBEcilQZke0cXfqg4qCC8kpBS37/tZ+6KUN4oaQehEDJQjLKAWekHcsH
M8vGth9UkX9JJax8kkK6dMPDyeEbHtoDSXfU5sbk0+OIhbLU/kIspcrYf1TlxHiXHbOKCs2PJ8JH
Y/MlUM+sm+LiCcYdzxuJXwxBQhnH4FKsxeNDTyxvadBrERnyDuKCjwEL0pZGVmITR+Va00G6JfRE
XXD9Ep6l5l9R/Qy1FLF1MjmPICZl7QmQ9k8Mn3RuEFTNF5ggyHS+wx2NNDy5nDt9Qbv06tlPJOB1
QiLKKTz7KOE36G255pn0vmuP1VHkpCw7EX+v/fYr/8ksc5bqebKU6cX/DhfWvZaTbE9LFb/iyPy9
DVTqoBaqY44cQEr0VctsHwFUMZPkotDxe9QvdukR5jQpYc3IjjDdHeqnWUy1nTxgA/ZuFEw9sPe6
SEbXrzP/dLdemAqY1+/mnBLCviR7FUaHEMauEvYP/jUpBOkHYu1VloBYrlY/WQvivr1JU80tXNy8
urDP1liSdThYxmGTKz9tro81Xiy7TeXG/NesGgohe3bn7GXAw1+ZaI7p9D2u2EoSwH2BvyhQN82C
sV+ktwCi3b+p1bVWdxhBX55WEmC11EAHIJoOES+EWlbIer2NzfXU8UsEZxywHKx86L8RM9CwtBYm
xmPq2PaeORGhTeaHLZ4FBxnrtATIV97zbzFIoEJ2pC3GF9GeWKLEQLCFBiBlUKDA+ZdG1j7+hSJ2
k5U19nS3UyfbZzzdRHtbtmkmSYNLVPJPyTSv6mknXOSGXqM9O61CaAEg0lLeyEc+22wlXcUgIOyY
gk48lUuD+LdJgHdtzWkI7h4UddT3nhpZ9N5z3P+gIzaTuIycuUPjka4YcaADP0Wo6wDSnJnm8eaf
YGQfmUU6wSqHjc2rmRWjm1L6TVUpgpton1eMhlOst5oJ9/6LOlPOr/jlhKZ8DRhH8+mrSPbSp93A
dVq8BIGTORn74rZYXFbY6+iRPSwMJvNop7FajzpBke9zpwmnV/eAzOY9kmZNn/G48kr6qAfzKQlS
1qvlO/7RcvrS56cHgNJn0IkEMuzeayGi2Nz+X6U3mr766D0bx2NEMEMxRWH4u9/0tAWT0aA9gHwH
Cv2QP69V49PzQIzNOxCJOmLvcvW77uW2JkqwKL8UeoLjr5mxEHhhzZzfXgMZPX//wTG3W66cHGps
o21BWpoGrn8p/p9JjeiqOVh4gI/H518Ovv6Qu+j+qWzLcSDnkbFZz2Zxcpp4utqrQySpm6YxBUJ/
71V4BH3b2C9vh7wXazt9OIJ6aVd56NbLyKw3mzB+du7M50FypXUKkmQlUU39X4CW71z5BDiIkmIH
MHvzfCUZMEKf0vUtMJqzuFro4MoR7UKaj5vugBtqdXq6ts52UlVNo1PpGeATA6jjxZmJSSe/xRnb
JTU8q3a7oIlDTDPDMs4kR992PuJoNR3AuatzBXoQpwJsclfqHJWO6FAYqGhAz4sB5bcULPafk9Gy
vrx4zC85BZzqemcy0wc0MyZ4lDDXsWedZIif87T4/JRz75/38IsBbDSU4OeoHu4wH37wlOuxqwQk
13Uf/LtYtOcF3Nlva0RckH/6tgtY+WSUEDApS9nmnMVN8Y+F43c4SI8yxcXbEQUNpYAp9BICPeKK
rO4aGAEDAThvO/AQs/YsI+79avVRnkoWtdzoRg97UDvxNPSXKvULRM8bVagz37oOJfBeWMiDRu/t
1T1f9HzrcSpEHy2rPoYPxFgjwXD2AcEwx7TizBjmXpEmBCeo9DPYWsdibbsFvcTR+nUofSKdT8NY
udxL1W9MiBoDFIs6FvP5hVxh3RYp49RFoufN0UHOMnSXtliPTgxC1dPoS5XL27ECUKMgOZkOg+db
hne2SbxGehdrWrNbsQOFSKeCUiiTqBrbj1fuB+6XJDMHPYN8IM5TrGA9yHzN1l/0g128Z3FIdJ05
4cp7fyO6j7iX7igx/W8eW51DIbXGj8ugEFh2vPQ55+RRE8g1yyxx7OzlWIwtK7MrP7cfOSeE5Wbk
CLl46ErMrO4NRCX2Pkd203k8xeETGdkh1jRsuGC5mYZYYWukKU2KmmuNcZLg3mpsaB9MRqasnrd5
c0/xk0s3O3GXn5AUQSNtq6/uq29HQ/oqtPQENSd+qvOj9fnsZw9Cvtl3yNFAip29NMl0mxrEs64V
J3AO7mGEBrWwah416Owzx6zXcQY9rF1rUcd+OJ4IeFvysexr4ttE34uZTJEIDcUnbm2+CCzVAxCJ
djDsomzM6006IaF8BE4pZeIN2u/C9V997tk5eN0EvlKlVS0H4SbWZAFg3xZ5inFUYYyUqTA+e/1j
N+fBpx51KyMq9lTyhC/DQYMRBWxqwK08iVhn22OgQfl1Ue9D4U/O9yEBatFVi8asioZhfv1Km8go
Jt1RqwZsBlId5Uv5aDZxM/rdJ1ldyyzfNt8oisrn+YxspkEtrdBu9dNwcF1f0a5UZLA+7vZt3Tte
+A/b7N5cO+qOID2fCBZt6JZu0BfFP9RWsZ5jbQyHTu508Ir44fftux4u/bYI5rldwCnqYqlm3HB9
QH3lWFA7kd03JZj+1OWmzWJWcZGlk72P8b4JF4nBadn9DeTMvxUBRDNTNSWMom4cKMQUz3G1i/Po
ToLt5o8982RInnvv1E1Nzq0PkMmk1dj8sWzZdEKmYEjxYNWYHbNhhkNQxQMP9Xb4nYe8gMCpdp1p
rYn+KO44gCx+pSfRvHVd/IKMDr/1/hqb+e8YJvI5pxfZvsaXtzkIqGC1s7QkZr7Tl9p4so/BOzMk
DY1J02Nt2xs6SU3mEObB1v6nph8eyVi6eOxpn8iwqSkg8olaVu3QKy9Jnk8Sa1InUhBoElGI0fzv
deAnp/v7FWsOb3qygfgLdAxfyhz1LS1ppbEM5csUce9tyiGWI98PO2XtnMkK1NsVwojmt9A8xDGt
4/rJ5/zLQH8kXSYgWprZW23OrMa1hLQTjwaivhvPfUgCa6GsBmc/VzFQ2P/7mvn6166uRsn6lvfD
sC6BJLvrBpssRjC8/mlfQK4sHVg+Gq0BQck0qKRynznE68pyTYlpC9ZuWei9ONB3cWMxyqa0tQbg
p+LPEAT18dkq42MH9279JhpnbWK0XX5rPQGptGtH2sTgsT5ozk+f+D2pFsEgiiXKRYjLtx6uylhH
YjDyPl/LVUA1bnQBR1Xi6UCKNcVJ/Q8pmG8wedD5qkYUD+t70/lWGF2svCV22Lgxu6b47WLWww1T
ethXCCM5mfAnOT0S8LfpCsO9HuI35J4DNPUIh/dVw10YszP6ECzgICMSrutB5UCMoR6YGu6qG28K
Ygec8tg+lAQXQZ+gkEQu58s08ilhnCs8LFSwfN2vojOvuaC9NWMJ33PwKT2jn3pXtyp+iPTqjNmH
IpJINV3WqxAZgwZgTUTKdvlFCb1+SOAIGirQfCKMLQ7wnnlxU1jOCt8JGa0WTA4YgfBzSBSWNqU6
g+xf9I+3v8C7I5Svu19O4pvd3GoscdBjbEUoalFa3dH1T3dPspXxppPVg2+jhoWgQ2XAifPXsrC0
wRc/irh7M5DlyW6h0riVD8y1gAVAgjk4HI/+qBzFN+/iumRe3Zq2e9xR98V8TUG+2GPrRChkLBF4
PcCh8rMOhvbUqlCZHJAFkN6ly4OIrzPf4AswUtwCCWDDHvQwXWdHN/dGG2xUBzQlNvozbXERxac2
N0ix+41e1rGDwo/ZbEz3H9E02SEOdcX8gUWNbl8gk8JsjafN1vmA9u5pjXttGLVZk18HcG6pFgKS
CkDX7f0iRwbg3ACSKvUjel3ofQDSxAZRNGVwOqqFSmBzAgaa5oYfFzZ1aXfnaW75mEhppDmWK/XN
9fNsZAmTJUqR8W5NgBTHslyXeKwHKsYZFWThQS26pWRcGkld21lMODJI0OotVZBXCKDUC/16g5lM
MK8ECX1JHlwY5k3+CAZHwLaInJqBzOCpkXCMEfRlPlCYqIMoH8yIv30F/jPEk8yhXuhDqjnMFvmB
WhuYrrzkJTFqWkO06sZuPznoeLcZR1Y7ApzHRhEf+GHBwO4wrce3o2n5ZDhvvy1tAOL5bKmXPtrL
K6G7eIFXjcT1WFxhWMwJrZmbmbS4KCvUDn43R8TmPlwzUcl8Wgu/9+c99t1YMd0DKk9xLNlku1mG
OQbGGbd+8wvJpOtrWWlbwhQljcEjyoINxkh60F+JeVjEyqC5m0BietgauDv8lhZWjcOrplPpyaaU
4CBiB8o4LbwYxCqOnkJD/7I9jLunRLQhuZG2IaDu4LJklrTCA1oGh06Rdsn76HQT4kKkzgkDW2YQ
rgP0PxWUKyc7e21tlWMS7jaw3p3UD3gS4JlyYCt0U004fyrctuFREdlVuMCu6qoBgREpnUnlpEcH
y97Lg/BkEwYYupN1ynWsWGExDC1rxrIMzl6a7xmQMmxMWEsOrxOHuJu42x+3dt9PwPZ+gykfCjM8
Nc7BPajOFUyqNZosRR8p3DEVohuNiqzzqgfVB5nMlCFS7mf+Zp7pkmsvh0aV5X27jrWRUd0uvU/v
2NXqAogeGOsHxU8d09/YMJzb9XqFJrVJIt7jiGus2Pm7Tb5Mv1rrZvEE2LPTcREki3TDEaoiIeEH
e++24qdc4pnSudW0yv/XSHdMEq/D3d9EtRWLc/jMoWXELAnzdmvFJU/48ynDK0ABvIQ3ZBNvfwF3
/Hkuy9VSTvP8bcKS3Ruw3oKSOIq7PX/Xd1h0ThsfQOHTLBz4GLRWDhrKflSVc01GOPmPg92mIeGG
L/6Wpo/5tJGWkVyIXTJbfpGkyaCEsHRFbAyKa2vLjHgFzh2ndTRApe5ZGaBx3wEqw2+jdCDAG+Yl
1IzL/ySYKhLFIH+8qW2i7oj7HDncVK0hllwYOqb8kOyRzUsI3/014+acfhsgCriEDu5/5jJFBpCi
LXyg0sTzTqFsIGcQN/omlJtfYvF7renfv53uKEbmJNlmI3eqbEzJiuc8KbcGBM6YLfcDDVxDwAaO
CtIT+QQf/H0fbl09L9YE3CUFPdZxg10TxD14VXdjpZcPCdUuKixaz/vL4ZRZrJ32Aaujq4d8jrHK
jid+hUhDh+iYsqx8A9iwZ6IGb0wHGAT1Cdb5xjYFFJ6094sqME0lF72VR/hcD4/PCVC1pRw8z5y1
k0gi98J1d1LxfD9p+5lrPu96V/ErAepEJYO/6a26NR/bEv6XCy/HSNNI59eXwUpZZiZNN0PtSrnL
r5yiiacJuSL3ihQkzY8nR3+V++qgM3YfBkjHTD0DLhv3LNdZytHztf7JpkBJiuTs9QNniYT3CBV6
FbIHuJuKMWjBRGWUs3YRlcdHi2Wlg8sMvWrTMekKqnFywOtukrSZHox4YmzRRstViwzJI/Bau5i2
5nXylDA345Sf0h9xz6xXc0Ic7Bpb5Z+5ybiGnP9oPekxAmOOAVjAFl64aQKeUohSbZp8smgC55ji
szeBNi/7A93iLsRcumhFr78VX49spntJ9Xk17Ax/k/RH4V6A7BurKKj7beMpYlG5owsIEIk+gS2H
EB3xWJyEUjl2VVYg+7LPlsZ45akmp982y10PLHKp8h568lPUUcMs+JGwtZHVSpl4FWVzD6SWleVy
YGhL1IcJyW5IMwqJdpEfd/2F6hJZrZ0644xFg2N9z72GbZ/+3xYGhAkvu3JgFpNkvImX5iPfBWJy
+nfqBR4S4EZ66YqCu3I862LO5TAjUUA4E9WJMNyW89EztBHbHGrb5Jn5U09wy98wGHpbB/bCdHZQ
+EQ8K6lR/ykFHLzWz6i7MR4q1nAgWr3fWlR5wCeiNoCHhUFxQOeX1o/2eIEqM+V7dA5Q10O7RRuW
AWPS2utQ7FkLjYtJ5UP8tIyBAuJAkabjS/ur//55qTCZSmFPlx+ExQg9+PBSozhsfNP92irUIj0A
8vuS36otJF6ElDt2Vdu6jw4wwgKZNiAyyW17frHrA0kaAXLHd9FsliHg45iZEmHtCLc79FQ/98Ha
Can7RBY9XfPxqlHNn/4+bthfeT64y1suWRaiodzeLs+ThaVzExjmC5uNd02q93lDdkWc8O2PbHJT
9ndpcMXxp36muwaT+YgYgHsEkz3eLPNEaknORpL27wKK2cgmKwsyL+oCqmeb7LTHQPs7iEa1S+2A
TeIwe9gVohzOqickkm4iEJpYtp4ECzee/DO+tyLuVRjaagEKMdUuGnC2IPQhYv1M+rfIYdwEm5iJ
XWMLu6Clsm9eQ1MjfrWgdzvaWNP/gPj/yEup4A/I60wVNaxszmLXV5fIyFkptmtAAc6pdsWt9umR
kObsFECfdZ/FUPgO2QoqY6VrVZ700GFTYTjIPIhs3yJTHg3078HP5kKwgA4fToURlrgphPf++7DI
8PZa7TXXrqi1FD7sZkpwiJ0zOb3qNcXQ3G4toTCM2sPApaM8GMJJifTbsIk6mgqHnM8TO0r0t04g
QLN1R14yLwmIZg0rF+3NBx3Z+GTfmce4hqBcDLhUkFs4zU/GCFP8HJ+lGb0P5ZIq3AZxB73gYPLu
zko9UZujyu0XXNHkLvgqOYWWYn17F4r6WZQAdVCEFygXaEVxL3LYm4/TuayJ3W3r1rV+m/gdmTcT
jKRB1PZzmFzwYr0kpNsva32A6Fy1yg/MW7iT3lPbx3P6OVAMp51PHzb5jTnfVux6R357nFN71yrX
bHmP4oUDQcMS5ILVYUTllRqCjoayoO3Jd1JwVBriVPhDa4FlvpQWX0vnYIRJbNWR3+ssjdtDB33J
UEPhwMHF19X8kbtNVB8sGEMCbD2E2VWxOdSHWz3HwgaKHmUKCBfwRMHdUrN0ZX+J8aTz8WrxipER
XO2euTiR5dEk8XC1pzC0Eyuim2Ayhp7W1stndbD39a5fp0Pt75VZB1HC5bJWazPwbYY8h0shyTsF
+EWnAFOyhuJLmSqbFx8EIlyGGcPHUxhi3gZgfEc6nvzgF1mYtbXBIQJCz2ug5SQ+9HKiYuq0v3hw
1ptP/7o5YM2omLvuCNbsEvtNBKZUMe5S0hgEwrJpcsUiU9O9FjzLLdJQgXkvpf+XocVsHPPJ3Kx+
0YkwfrHfclCZ4oesF1tfZ+6Ff72H0OYng01t+Qb6j0xq+NCT2PebSJU8BBi4/2DGgrjWZf6Swazu
E2U+cGQJosOBtbfB0xIWaF84wG/mOt9DgGujk1I6+DQ7w78+9yBhQJqF/MDfuo9C6WDahMaklEMV
ZoPaBZykmB78Hxuc27kybFdaTz3uQ4NduVyZRpnWbxvWGvASrH4/S2ifPYZ63BgxQ9w1bsCIvLTt
KPtz07JT68oI3f/FWI8MxKk0jXStvNCuJHZ5GSw9l0PhiTtmpEXSw3BSguq0TmgpMRm2p2Z/J8NE
E9ixJTP8A31wyz0V7zvOqCFheh+SBby+MR33H9xqVybufU3+LI0KPKAIaUXdOUtW+QRuJdfg19By
VvqTTTkrdCS1glbpTU+jsRlmunnWIGTKQhOhdQomn2qMsPiTp/rJ1AgY/h7w1vFwTEr2q7GGHJgO
iFLwQr58fAETX2jHlQmxl5He67knlEqrW/NmcC/tj0/Gf1OSFoBzIiAMKRRqctPs/2WKJKTag4mL
h91DD6kOM/makm8wpGagqxntIxm/7rQASNLZq0OE62Asx72F+ely9JGkjkXLLzlkYtd2KbCanhrj
ijZ/E4RJJd0MVOF/ZDOU+yIa9iLSpzWIt9NLGWWZZOisUq7KDYcHnUgJMNkT/9w+8fKyb65Sl5ve
R80OTDprBHXGCUg+h/YtpVxS33db+03N+WbyfW4ZGf2GxivdoEZtVRIl59j59f62MhV7cSA5d13+
ZAZt5SQ4q4VCnJZM/pgbFbDWG4MrQL2TDZEkSicUpOFK6AVfCpXOlbaz0OACnXv6A12YueBMdzcn
Tv6jrsyl2eWkuT85BQ8vyP/h27ObJ42dzpfcK0RLObIpBY1nT80bkh/GwRQ71EpmD6serzCSuCmb
47x9SfaZS60j/ZpaeJFJACYZHBlC56Vqz7e0KCG5HhZ3UgzlncxxGYF/NHF2ht9ThdVGCpPG7Awq
oFAT8JJpJ/LShe3lWul9NCTJpr6RFr7bKgyUskfvWZgpOWCCnwaOGCKzYDKjEekwzlPjiPPN20yw
We4WbVtxjQEQaCR7QtNsGA940XKISBohNAM/XVZgwCPsQ1E58aIbUHH6kWeVvXJqzGjqR8pH5ovR
FKyJ7sn8jF1DzQlzeriB0MzS1PKARLkf9r9ikgRkaUmX5u7riicUUBNZOuA1OU//1FrORJUkH12x
nzjcDDa/vbvgVeOpI53Yv10dj8WqVt7rLAhPWFNd4v3lzABnJF6xkgoQBTP1spkwsxtn6uzJBIrc
RnROjArsB07EhzA/3X0E5Xgt5eq+dvq6gtp2KdSx88P0ZpAUPq/rCra6EBcfFGznmkLy1DUzXtQh
CfyQ4rZrAzz6h/JuU5c+YHr64MQfVcrWQcG+Gc1qUaCkbyfeBgzzddvy2SyCezynCNRUqGBFzxz6
J22ioWtd1m/mEdRr/388546XFLSIDGgsqsp0owlNaLX4ks4k7P+enz0VYsN9lJiB6/pPGpFGwdB5
UpFdfen8beXcEEXszxsLxzeH+FkRwyU521koe8/JFM6OKlbZA+KTCGggQlo3QAZ1JU2j/XWwATf2
FRwutm9SvuNr4T4mAxW9amziHn+V2PdzllHb+RFrs+yCUXv+xljI3wMOg8e0Q1Y2BBbYLaKS4w2d
cjsUclYxmH8KoAxLmy4hBmc2RxrDhFL2U9FBxUqKfmRmQ3ld1xiVx2XTrFeF8x24vUtvQ0I6VHdI
Z3A4cBUM04AvQTpFsCmouGFs0/WxEBKrtwX886ozzq7AAjqBgYtyCvmJjXHzABhIyIVzztXSBld7
4KT42gF2hxf4xMGNb+U1RDVwZZELb7T5h89hZurCExHFAPMiWL9D0CWXmTbkAR2Dhktx+80GCpV1
WHVey8xD1heoexSfKGF/Omp5yPzbTBJi+vYRmI+OoliDLBQ7h9bY5Ua7v5N4XVcu9yHWv/Pkzh5P
L2/d38Pvmv+N1TT9v8Ru+muAxqXh85yEhu+lOg5TD6C1zIq/yqMbLXidg2+/bejA+VTHGZcouleD
Pws8Ipls9oXrLByXDFQ6X4as1wnP1J8plecwmMObZEtP+h3mTyzp9qbjO5yqur+SHU1kZA0wtpX+
jfTMFN/9KW6CP22SJOwBNpulrgJFd00MXSF35lq+G0JOCzY1VvMUo33rpe1A2BlbyJUJJN8Dx6ZB
sbfAd51mtyRLugKLU5Bl0NoEN7FHFOVCd0rNWlDpLOuPU0+lvvwge9IxYgCWqxBIltMtLMenYKtL
kOdK0g6HUKOYqzeMB976IUrmbroOUIBHEl5e4XJ/nCWBb8q7zvhFPgFs5syrGCY53acPQzkrVwzw
nCXY43Art17mUTv3fuoiLmkh3ijl+bkL+16T98Szf3S6iQ/GFceg5UHig7Z4uxlOtfryNh/UQq4a
jDeOhf9oPR100+8wyAStvpmO3VcZb0DTa4CIsxjRcKh1XjKb2r4cWC7AiqcLH6lDuKg4m0Xgd+1M
KWg1OeP+PPY+Z2dmBg2/gAxaV9b4w3OpBzk+EitlKvcDcyMbYEhxWrqH03IdW6VykFip0zyJzM/r
TwLI6JYWMKqcosrpuQ4GCI+dgnHi/6qAkTByZXpeJwy5/aoYMfpejqnX8zDW+vN6wJ5UJvzgDEK0
j+lnNJrdFyhJJEFui01OoVSdlmVNXZkuIoSFRHmsNbg0BOkaaHVukm1YPWbhHMnCx5wNKjpT/PVe
Fe3c5vDBOejd11OoB2wLah+fk5iqgX7SEKCQe4AuDBNsH0AjAQfwvDJjpnlSmOh9vILXFzcq/K2e
09GGmlodqS6zq6vwfWJtT+UngpM5hj7uobwLyJn9wKj2gYQmVCDFBWOL+BhcZqbOdfTPPi10GGBj
N1bVzGpOipY1WpjP4x5pY7IU71lZyPxZAUuj1bKewztVYVpD3syqssCLVceqtD4Ayl6HHqamcL8z
7ZkSQnKQFqdcqCNtpIVNr5RO98SjDo2hgk7lPb8RheZQcfdSzQOK+E6LJWH4SfF9HgOxx5C82ESI
AePuMllyCcbMRSVjtH/GnbLsqeZzuIY8t8opQwVG3gk0sX6InzPgW7iBTE/VEe+5ozIknsDIJoE/
IVdhl4FF6pkwAAdB70pNu7ORebL43WgjzRAzsmubpaIMK3N8c1xE7Li8ZQ1lcXecYoTC3Ezeoh+j
IsckxB9Ib2pAisuBFT2d/F+C9dypYkH8xg3la1GD31eLKKUMmBxPk95C4rayuODHY1yi8vSsNENB
pAjyAKKpyOW0qk2NQ3Hv+Pk3nNt/qx2RdUM5zjO/sSu+vVjx5yrw2sQ7DaH1BVhUG3cu/ADEn/ZD
L73q3qvDf6jGWsRyjuIh8Pf+NBgXd0ItdQd+aUpo+n9HceqbSr4doy5fVPdQxFd2WBvW03l4dizL
IQP3m0PuVyXIIWeuleGXaZopfaNPVKajkxnG9JqfiDxck3bk6gBqX+rXDHXlYptFVKaHuTl3k6sc
RXnKey28bMe7QdcW4JpWZ8p4cjgtLeXQ8BJez0nglbtyk9anhLIQZl5ukYo26reokdD2ziUBlT/M
TK4IKe6ss07eRN2uo5U5vlsns5kll1dOKEp7ek5K0GC6WsrPvWJksz2eb+TeWUJrNZk/JoAQhgoQ
w7TGy8HPX6bI2fcZZiiHkCr1K8iEgn5M52Nkp7In0fJQqv5Rem+vwVLY34QsqCAgcfdt1mlHKSAM
3CT/dP7Ggq10rtfVMO/0/K7wI3mkrGqXZgvKqhmKEecGysJBHyMsS8MLqN/mbOMZfCYiah9oKBBq
pp/1HtJCx3uYy0FtvvG+R2Y3sV7ckQdjI+TVt2kp8msyRi/l0Pv9zNYvJu0+mJtd30HbWF9j+02h
JJbRpwrmsi1ZEwoq9xaC/FRE+W1uTNWp7Eis2W0JgFyoJcahA0QOZG3OnLKCNisvCiqJaMJ2TgFQ
kW0yBNZBcDpWLTxW2s9bFHWQbZVXu1ucCFA85lBYNEimw76BEZ+r0W/kMpdy4gvBcU8LcTP06Qpi
5mtEcEVuJysGgOoorc7yaYGr0NS5I+39uYylYvcFBlKAL1AjEWT+k1TeHJCpRzEPz+hPsouTjaIG
NDsyQ8vGkoYqW4MJ2+WC+bQqPppOHwVkrqAYJdnyk6oVmLqT9AXhaLKtgZJIjJbdxNkVvIYlzbBf
lgq1ziWiQCcnET7QvsZvFIfdcsJYJLRDDD55UNiQO9G5ldaiFB4Oz2Ockn3vQrFSS3yxAtlgwmim
CaFPy6oUDcl6Xc2wcQwhX662Jec9r/aAASUEZPxeq8F48TcKjrgK0Pv6mJD3fNlQTdoMJoHKDp5N
TH76TgAR2jFZt+M1phsVpNreUT0cLX5gQrqtX9MMWXcAFPVIip+82LxvONRI9eYiB1RI9eIMBza3
Gk+KXI3lGClzGaPbiSj7gIaaLkFeQopDDosCvIVRAL//CsgOGXBRE89RhdjvRierHh96HwG18yek
wVMubjU15dqHjArQ87E+dyzxn9mbKDtklmRTsTQDdDBKqNXFt4hYaTXOB0akcKaQGsMZHdmr5qv0
uUTk5eu92ncNM4PUGVX0peCEaMw2xAzlgVDzwgFESzeP0hT7k82J0Gp9K/FG4e9AIdHtH4K/yVj+
FDoz10e7ta3VSadD+OmsW1RMWUAZLqJ+velqaqOd5MgZPdfK2Kg+6zhmjHGy6hqZ/dHbHNz3ZK6W
4nF3/OB0oERBiC22yXSdl2gieI7F4tU8wUMeRVyibXQbJbOo6PxXYi1ylQHWqwb1z/XTk9m6zo3z
tTwrvX9Ab1dMVCi2bzBEadNZWiT+9f5wTHkO4VubzQDsHQPboZDBuiME5mGQ+bi4AhVAM7H3gUiY
h1l3doRzgj5LKkSWnbRioaRHiD67BsHjzVYlhPoUmYbliI2b1hpBlwKei/DDc/mbsYJfo/E8lHed
lPrNUkCy6MKO4AtAP/paGdyo+hR5vapvOhJEsK2fkDcHIPCeTl2gGFbIK/hYk13++kMPN5ezxrVo
pXLYs6rWK7+kZo6ucorUYRM6GW+zKFeCtX9rkzpHHzVUUSZr8S1lkVRbzoUaJ4iICKCpgc5qjb7A
q+FGsazCCCAWQ3FAM0fD/WunP/2MnfswSgh/8ekZWh7ONIryIsr1jJ476qPHDzOZfNr1x+q3zt1V
LVp+/PGWGBqFV7oOnIlj+jZuNy57j5BCLAKEXtpXYD1K0aO+gtNr+P+9Sp+ka/Hm+H9Kxlg5LLh3
zcOMogFf+Cw15A/hAPGXyngQ8k2F1Ihx8jlBjLbnUbqqimgBYROWjX53RRu8XPVS7zA2Kmy9Y95g
krfFf7zalmoN6dumIofDs/9sZDLuoyVO1OD4PlMpCxbsmRp/frrGhnQMrBzaHmGQgswVqxh19pFV
QLt7UFms+CI+Xrho/22mUvVCJC1fqEfWiqjFJsK1XZiKslARpcthG0wzr9Nk07Fn6zVh12CpNqS9
oHEJwyGHHL3L1qCarMxzmlafzBQgx6fIezsqtv9No1ZJqUFvEzabDFnpfgcft6kt0VuU124qaxZF
T5s0gwR040SBUXJUE+Tmn3UNfqOZOQcC5oiCEhC1AQORrv/h5MS49V3w0azoMATQ8BX7ts3lEAdg
ROwDwWyIHhdoXGrdbjKAEuy+YlWAW91svC7PEfws1vQo3CaN4R7lhTT2W3TlcyiCtUGEe8v30KQl
CZa+PH7lugBD81zkc55eZ8bRVKpJKlCO/SIt6jSXctN3s+aSt5BLQljWEgryJcEaHeUy/mV8KPDH
kmxnU1Db+s/b4vQ8mXusILDWEp8WDIIaT5EAs3OeSCfLa61/jOQE4Xwy9Um/EBecseE09Q+F1XmO
dY+YAp4THaZJ4m10JJqMI618InP8S4RdvpB8KEn0SjO1j/sy2iM5sy1jlSBsfw5dPOmrKnYrKIfb
2JAMZtFcx2pwR5C7s2SNh4syyXLQnqzgmDEkOhT+XYpiPDPLeiLejSs7bbJPTgEtwV/nymZIHeeY
k0QseLZxA9aRJt0puuAnTSbR1CBR/neL1TDfvKdtv0kpFARuZ8/JZRff8BXIRKbHtNP0q5053vtn
mYLYGuDGzFmZXTiVYpLQ1ITHih1l1sJIYqFehmCXkuaJp+goPwypbaiCipr9sUwpAKNofTJpXTvX
w40mXHWjhx2Gu10jIy2csgmtvouLlLevdniztd2gFTzQ2EemNIjIebQD5WjLWpWga7Y5paPW+YB7
dUHP06BitxrXbhqxFyz6jqiky3Jmjz8zyoDrr1wyoik7ubXh3pNIvnp3E3+y/+ln1j0/wQpYVpdb
dSuJrNCTy2/3VfI2bRRlNKluA0t7K+lvL5+l7YBPVE3gYdq2Teo/K+TbIVLPgdrm/V29+6nCPjBG
uGSanyvTFaXk+ZRKe74LpPl/8KiomC6UD5eknX778prjTlmhfPmr7jDuPcGLr1Sfkp4cf54jXAjS
kz53bxMKWbJRrkXTKOJuonlfTwa3me0VG3j/oiS0GfVQn5cZca3JeRYmAbQXmVnixazy1ZcFAyUf
3uQLbk2wiqIbxWqgIykQgKz77WwOIU45rNn5jJAPpdmTUKZco9ClWSiSGvlW/sajwhsWXNWRQVSy
+ZCSBbqrpcg+dZAmvoNbjRKKnnWk2dZHDweg+iI7571EETjFVGIaBczQS/1vrOzgZYQm0avt6aT2
ylYKAQeD+55q29c2dJxAu5m/O4le1KurHpNm4rSCWp/UP5fMZQXedyu+CSqgU8Q0oTS/XhOj+wKt
2ZY5QFClZ9WVn98RGsF6kTkbm7R+N+k3roxDUgesK9T8Rh2BVAy2SI83iJmFQJFO/dJmQL6iRkaU
WaJN68QyalmZ0hc5vPcfbfJ0HAwYqO6IPJSosc92yv7SBwCtY16nd95ELjqnGdh/nPbv1Z2/KT5V
pRPWd0Fkqdc3zyaPEC1kRQmDZsAaRCbZ6zUjOANiGQ1ZL4IZi0CQS199YG4YwNPg4EgLEcSbhr07
DUTvGRsnkXKPnS5x4erJEO2W1Aim+X8VR3Yl1FeLKXEZlHvhvG0y184QpDebnCjS6ALx4zCFJtsT
rYRBzR0q6299J3v09Hm1qLqJ2FqlAk/wkNa3IbGmNprMPsHle9rMbgC3xuXOGj3ZaWQ6VpeCFro6
rdt1GIqnUk876TidG1Hw9DRtpcKVhdVWA47iyf+YcVakHN0AE1vDviN5Q/M7WZjwj9SG8gJCYqkI
ToDgjinV1s7IPrK5qtSIvOG5NFCubHwaRVy/XUxOjFeDR580vDIq1Ht8+2EReX+LYfk7UQpJSJlj
mit4cdIDzt+X9idvsdbdYdDMHZTiZlm0FunCAzGtq0Fb43W/M86+tGYDwfKDU6imOaXL2bNvsXFf
w0cXNTRtFjdd3jyey3uegJW9/AyN44JgeV7FimMsYMHvM2H+YtwPNrXDv9hkK3lkY3EvArutZWsg
dm6OYokpQl9lmrPPPU2/SGc0DIZY574T9rkWJ7HS3I0ly1Cm+ZSxMy21wNT21E9FF0vBBBBSapiu
cUCG269ENRvMyK8AS/WHLFw/SSiayw92m1HH8bW12nQcypeFlgcHqjSuvPcgcwp3qhJuTeTFPEOE
j1r/tOgv4tQnj81oTAlCrnsvE/Rh9scgd25023T/v8a+BAU5OEXoneQpuK8gol7EdJ/nqQHTZktE
TPztZU8fz4IHfxliRB4l867ogwxG75ByzQt0JvlQC/HUhCIRF/jzc36c/zuX5fQbN14h4Vwinx91
Z3NImTPWKOvH2cJtw9Ax2/BHX8DR0XzCLTtUuPgzDgufJQi1hXwHNZ+94CV33Q0Vtv6Ocxvk71fS
p1nbxOacW58M60ZZvwXPsPBBpmOG9WwDryHm3pO8kmsWlgU/68JlAal48f60sUJopXzXmVeVBxlJ
6NaqdLSye514biXdQohlUeYNpPQzZJvWWpPXbYyJeI8txYT+wgQmW+P70n3BsxdBsQQQdvtUPYji
h2PsiwI8SSDC+H0x5BN1qtpg37540pHmcWB+1hbQmyBi8PLOzpX2n5ZpeARxgb5XPTdbrSpMjSXp
fzpZ+pnKcUR5gmL94SWTrOf8Z6g7k52qgPrdUUObg7EzGFPfIHP1g+Bok6q1j/YidANV6w0gbi/l
O8OdqcfpHVhdr26zSkOB+LKrLS+uwgj4qQssU3dxm8XKgIYEm0STKiUIKVuehiVrj+fTM9jXEjAm
eJTYtBfZ9BCTB24Xb0SRrpuBBIFUcPuQYlE505kcqnbNV3kNpI6O/LbD0WFL1oMq4sanjf7Ir0W2
VSXXWbadLbNOmY/8Tx+Dnl/yH1FSjkf7fXzHw+GiYoPyRpdM4XluQV/b3aSj2d2/lwDz0aS0vCR4
DIiDwsJWayNOc3xWgJ+q9KrBO5sTzeznTKfrydNA0ElYQ9EG3S9BxtMhFFGlL/ccJJXuoZBslueT
nrlp8U+fCV3eyl1oj8yS+UZgcjG78V/A2Q6sKppOxuHCv+myGvYTCwEIJP/Y9wfVseap5Uy8RXVs
CnCAd9Or4KLLPHk/7YkkTbKtD59OvDsPE1/dE06eyjmOT4BYkT4wdYmmgAmztb+EhfwcQJVtGirB
U8itm3qQVh8MCSVNCZOKmry08EL0fo16iYux1tjgvCg4spCI4v3f8wBxgMZTznSEdOb37BPYLsdQ
talav9Vy6VF6bvWXrTU3/Qt4H852Ypy/+t9VP31hdEUAwZzJdTmmdlpF/BdIlwMg2rZmDLA7tPkL
XKcblT2KWwirhSKllwxs+OMV755xabNytBWHKjcoZaEf5abeWQ7QtPjzD184O5j8t/99yHsdqW7R
lj9nOLhkpRuWgYcGAkugcCuqwRxCplQpNu2lFZEyaC85ZoC4+qbW5zt1YKudUYbsASpmhqANXRMI
xNE1oU9SsRQgF/cOGHiU2gun9mWyug5W7p/UptMKzRTJ5dpeI1jvMZgm0yvCZNFAgCYE1/ZCudno
Lsyw974vl6Mqoo2QOqTJB4bKZdWt9aLUEOzfHEvs4DQ/2NGZ5J07RDMo7dxOLUUy365OPy1p/VKU
irNS7dfnzsa9voMGGN6fu2t5O7p/iqprFAjnzbJIxNT1QWCXZ9r2RqWR6xS7Js7cd0NdJaagzu1M
6ts4VrpDbMsCgNpMw86i/cnAGUAvDi2wPoVZ1TPA7y9hDtc42E5D8+5tNDFszIlIbwbzT5NGXUSf
rg8TI9VVNlI00dqG0n1CKStBA84V6M7bA0h/3hcCqg+6Vn2UnFb+alxT85Whr9yfJ82Y0Lc8oZRa
9b4KiMDtcdxe2fBwUYswAmpxaYnfSMxDlLZ6jrBvnxD7xRzgCe2SHidGav5dfQ5izvgdJp6k4IHj
JDbvscdtELtZ05u3/nvg+2z0UF6rPg/kJYXgGD0mCeAdR0IqVF9lsxI31XoxDuwnHgWoDwareHce
UD61QM3imd14HpFghvgvBmYWj6gD9mwhtMEWmh9r9jglPiMWslVWP9zsbQgHikViS97+JdLk8xAY
M3glyltky7s30n0ZfQbJ0RCHobxnlhIPuit8cOooU+tt52LSPB5FCFkBvHXf8Atj0vGKEMm1hED1
90q/f87MzuotA8i18L+RCEPM1pSV0oAHqpzoqDMIJMvtrLfa/UN68QFMAUhhRHvLhqoKeYd3cdQg
fsXEZRh1QxaupwEN3ePvA+stDiWtz4MzndnTDNDyl6rNFBXVhd7b/SqxO31enETbyMghJkKUudY8
n03HRhCAMZLfb5+7dn7Bkcq/UtbsXL1vrYz83eO4osy4u7wtig/DNM2J+ZHrV5sBlc2jle1bApIX
uxnGmcEY4c6J7DO98t3aF7uiRXDqBuVqpJHbDgq8/UwLanAZcls/mHNZL+4Q2u6Qtd6pxwUjK9pU
ES/3XRiGe4CY6/irkVkYxL/gNDlFtRYpF3RBtF3kjtDAakd4q3ktXx0Lto/mZQakFvcqRcaV93k/
63kepuolnv7Lb0qCKUj6sLPgVqkNCFJH/T0HHh7RpI6pwFJe8bXjXnyT4TprrMtRaaWJkQchgpgM
HTaDLbsnWwRTqURDc/6eZnTKIH4S0cHYc7rdCH3HrbXsXl8KSjEaLnVuCrGqmMCBlCxtjLw0ktlb
/IgHx7ypUh0GLDdDw+Vn65Do6jPRYBkDl4FV8Jxpe8EtTmO3sVyrm4xhzFssW+e6vxowCux3A17n
FRKoikse58Nai+XY2j004ci9MMvtt9n375E8s2gL8g6F24YlP+4Vh20j0lkKtxfCJO6EXnml9PYe
beEPgy14HJNalKfOra5pcT2vFZozWOomkg2UrgOKqLkigLM6cR9uxCTuSN15LGEnoac9VQyuWM63
lVNwFCeHvSnCAnya63kuC0jHGKNtDEYZvzE/K1J8eSYlzxWWxryWM3Y36dodXxYXJ9kt5SATCwus
U4pdEdSYqrfMjFweRWjQX2j/x0TAfIJIf5V9ramgWxI/BZ5WqilJ4THdYEz13fmcIBdwGSZbB765
dFBqusNB65c1Ma7ACB//Mxt57fStSsVnD12YvmvSEznfrqycWhRlvu2/AYWZpM7XFNr9HA1JmoVI
OkJAy7LQbd8hLOZllypuht6BtAjgUcrQRPtrJ1NjDWu0Ob5ijmxNURBHtV00ElVOUsHy/W5cDY6Z
X4rOmPpyllxuW6/F450X1DwHoV5ipnp9pH7tDUHwosQ5yt5GBvbaYPWZPfJ5uXXLRwzTHLPo1+B0
vXjG0dmDEFh7ruaWdzKlMyM27KqUoB7fyCj7upTh4vmiCAfJkqpMhD8Fdwn+W87K7yUzkcmS4epe
ghRWvo/s+wsylEUXDeGkOWc4dhzrnTx6bDgSPBT7ub+DopZpqYLCriWM4eFDM2qrxCAcRZBBB5Tg
FpwXVxZ4zjkaNmGYjHl4lCCgychLgZ4qS9pryRAE71UQR6OSP+PWCOG6HIdEXzQyzaPQFIXzwNyQ
BYj0F66rN+HiYA/x5SBoFzsWzNoCasf+hu2zbDEbW2+AWC1+HmXMcoTk39M/DyO+tLSflvD1+YWy
jUtMM0JMCwuMj0QoKRDCytagkPC3VC/lSh3FSjvKU60EAPtmEFzOc7btKPRxx2TbSFMwKrwmOUo6
Cn88fERIAzhxq1q9zMVv65BVtFeoOMCHU2G2pVHZesfPwwbz0RrFK+xgcJ0An9N0HOtyHj0GedyQ
r1pGlbjJbmK6RxkKDbkWfZksAiM71Jba88G0EM/IbeTpsnuQLS+01xfFVgprGxHgDL3RxW5S5coH
848CI6iTjZE6MLcgvlHh/2hlbYWP8oTB8eBaJpjYxBm0WVAxjMgM10Dm594UYj0zWuM5yWE+l/VO
i0cMxpTu42Kw6XyjYpIDgjvmUG2ucHsc3GY01uw16MFvxN1fXKxJdk+1K+7BevBX5f9QoyOK31pW
1cO/Smh8UJE4ZxzyIo3Hx0fIJ/J5MvlZAeAFeOgcjCNnYHSe5TD45Es1UIzZg1lHZQwsZYgbje9y
n4F9gEQw/PcgeE6OSAO1ayQZpHVBPe0mOLqNG1x1wU1axGSHAOviOM6yBHzkkKQCsjuuHzs8G4QV
AtmegVhOuEaduZfgPSxF19oQTFJM432ci5BkooyYFyZ00TKJHSbn0tD/eDpIjS9zUZxASNcpbOiK
NrHJbrGa1WNGtUKOemxzRNq51Q2Cc39t8ZP47/5hUcujR82f1JSDiY7jON4czQW6ghbe0K6clT/b
rLZv4tePjWunqKbqC59Ov/0hU/73s04pktUXTUyFcLLStpOgnYp0nNGRWR9eDTtZXmmjzw8XM6Io
mbjSVwbJd7XCij81QdQ8QNe702c8ygpjJ1sa1jaAKupQKJHFpPLD2oyKNR/n7Wr1OYVbaVlkDp9P
mF4NmhUYiUUlrLGoaPhsDKeTUl9y9v+MrCmloDsT8EHpv6emY9j3UJmAmabkBrZqIYWkxwEAtiet
luk3w9mzPGEGW38aeqX6v75n7G+laKmLl+/r5YPU0AC/nMLHYSBP/F8je3u+c/zMptZCfSQC0aw7
Wuhr9ZWR4e6hgysuicL/ZK2qiGR3JprTQHVUIctuafgrpc9WybwOhTMOzTxQaQ/rEijLHd/+6xyV
PtoqRRTfE7QO4/XkPQqU+QTjKeNPp81JH4g/K8QGYz4xSDKfmGBF+YJFrjdILZjnKulv47DsBVD2
0gIrvxSdfk7C6s0Rl6ia5cuf5Gb+arQzxBtTHYpZllds3MMW7IqrfgHD32zP9vZge4guodgKE6T9
yVFYCtJ77qARH+dX/X0AEixZXZ9Mwa7ZGZJm57rnKcyoruRq4PHY/qxPNl4NXyqRILUEu55f3db5
pagNQRkEPvuuqIqeP4Ajv/Pty2aUk9fi4fNpgd8NiiEXi+hBXsUTeGs9MaNo6910xA/jMmzLSGAu
Mh4eQAfaBGu13+/uo/vInNA9O+qFVBHOmMGdzjWVolrDjxaZHJ0BV6C7Tv6pbdy6Z6B0SHX4nGMq
rDlffsydssuLtDm2Hdzn/08ml4J9glo3liASfrOzLyiQTnh6aOhjZqOBx93a+yNpCCZRnJB9+xJN
yhsygrg0Gaytvovgk6YMPL8laAjRPZdTVSa3palCO4xy+Grd86PRYnrbVGzUIEjHKwPrrq1dJGXK
arC329wYk4WbIyjbu5RCN6vADNqQsvovT3WzWnkDKZ6wR3W3IBvbk6wNDthN9kE1u0cGxM6R2AHJ
ylHyZUstz+7bvaqv+muPYKWgoRpLw2jbXREBSJ0IRR7ur0ldnPcc0ynQK+FRThjB1qfHYQKPp6rp
urI7Fg9eAelcDiuSZB3SrvZxh3kHrwHp4bEdbXIuzu1zDIq4mGxHjqnkhZeRkax5KHBiYhzzdw6d
HYgG8vlGyV3Ipk6PTxfEGPQ5DGBIRenhA92d+8DY8pLmMA06D11WVBkyzbkDZ0b7Vn31nE7Lnwfs
CS8ze1+Oir1ekPjt0g5nutp41LYIdl/iU9qAYGYRQ7YKRF6XgLPi5///GrtW0335Nqpv++mGW5Fn
hfXf2XYI+ICn7TPFFI/YF0wQEPwD4txGA+K9PD4CFJKTJ9qW6CUlBcQzam1V8K6fY+uLKBVVG2r5
/PGsvizEKTB0ljY+N0hvebCHjrI2Jx69CCnY4UfQAvkCseLC+8V0R5zdgRjJ/BRw5XhYXM+01Eek
A6OUtPXMSi3qtBHGvm4wqEVT8359GEeAvMEeAISmXJ0qx7IgecPqOIq2/gALiHKd6sS6c9t/G2+q
XAHvJgpgI413y24I2Y7hCsqXIq8GpeOTDHCK/vcFxYxMI8u/Zuv/mMLbeLYT2NnUGVfoQgjinfzN
0LcnTtwhHyZWWum68JdHUKJEyU6z6q42H5jzm4V4r3Zra+BAYL1KI7xWmlCIM1l3dyFdbhNAsJ+1
qPBvZNEC+DDCHRsA/Vjup/+Hs3iEjyi8GdB3c6aseswod3uv9HqFKdW3gEdfkcncr4J5rlPIKmOq
Zxn1+ZkyGVjUUykbdSKjt3SHW7RYzOPEEiEddBenXhj0szbXRMMkLl2EEhwJ8el30kZuYWXlyC0V
y/geFjMx13WHW6Qofw14IefDfI/JA19YFxpXcKxdAE1ZoBRZd1ipjt/9u18lnZPQ208axM5lbV99
Q2PW6u5wE/7rircBbcZrXS71sCP5aMuIFXZqXF/5bXChSg0gOImCP02mdIFcgUfDE1b5nyz9QO3g
59hqPuteXDLE9hMEhIUbWnl3b8fLWfFQbWJV+5dryPt/8WOR6cqqmmHnMMmZFaRFdQAB9F5d8HGx
XgrDjMEZ7sP2VViD6Zb0lihWYFhMs9eMVsntBkFtYTXv+MtqHVT4MRp3suBFhtr/epwC+edVzqE5
pQVOUHhPyRbjCiPc08+P60uF3BXD9iw6XF3ZGy3jj6uB6hlR4HGScdWjE+7y0K3nlFIJTQZV7QRh
q0eSty6Diqa0p1SCqKg3Zqo34ullVG1c68f4JjitAOkZV3UWV/aGHfcB0Y6jOVuveS693g0JhCGI
U8scMmP24f/0pzmfNUOhJVyOUCpMTIEs0l+zAMmsokp+9jTEz1g6pmz+qZFHelw8lRgJbw8HnvGd
XGFsZaNF2uBmS0kO5itsA2lP4dgaFgqaZmmCItFQe/r+qwYHXbhB5MCf4XRGv/djM0dt9QsW7M00
CHcw53rR0NeXwF6eGxUj2ztByibd8AdU3IB4Zk9Rdo1iuQa9RaHrtVFPTWji6YnwlszrDy8ghmsN
Xpri0k8dmPAID6q+Nw91bIOxF6oiah62q8xTo/qtbV79Hzt1njlKRU6au8fvS44yzkFEwKGqk7io
h+nMgErkSBKKIVttUtbg5dJMQuAciKmm+dV3RTm3qT2ecWsVf3wJLJ0OQu5x+TJdUME0nv0mwlo4
JgbvyBeGTuUXEMN9hSQttiN+8fwf2v1VXG00CUdApEwk950bSfBv6CtZHgjMTnZICfA7BIhLFg7j
dfzInHpEuXFHmQknc/HJ/Mt7L64BPlq3uCDOpC5cnn/skEKmfZyWdGL2iEwLnmWp2fYDzG3/hNwb
A7V2pWxVp1jbA6bLnfByntxUJXZ5MB84P9iXEbfv2stkVR6fZCioNfTZYU9WPS8+8cA8mgPMEZux
NEnzY2BCtLi3+tXyf5d1P91j/3wRk82n77LErD/mCP5lwnicYbvsxm/YIAb3pyNWsmyPuKlDg3d3
jc9/NPFz/gDP/yxL00GBQXMZmzRJirsah+GbmBs/vJ3u6KDF8nkSSAcwL5BhmexhiMmaOXTKp31e
ttEmuo6abiY8Fk/hurZgiXOrkHPbLEwpTpjf8vnXcvYa/JKPZNySGXWOxsn7E2+3BWDQciAzzudr
6yuB0lhMJaUsniZxJZjmxk7S+DmeausUIJU5IldVggKcu541Jt3AWx3Dt7GEQjsqAgDf6p2nBU3E
UpAL7yqRXk1oaLSbfZsmlEjj7O173v1pmBZtz0MlK92GgragmeJpWffBio9PYoERxaojE8ssBFN0
ial4xqGbPo2O+C3AzRlhMo+qrm89zkyih2EGWPf2r7pcmgTnWPEFPH7IaqQxmctuhg+Rtaf1jucd
HFvEB2bNetRIlwJLMWgPvrZ7YbeOlnN+YBLyHnkBvCB6kTKl3E50+jFENWci7jvy+eypWbrohaPz
RlSGbsK/is4NiaflY2D+ONmisd7+lP4AyV6kluB6DtSMjh0NW5/3CTusGWfWv/r8wk+fL7FZA6oL
X7zMbhGx+Wl1USzrxzjnUQ9ZjDYgwaYGqZ0sPhhmGq69me8t4ZQdjT44Ow7/Iwk5bi3fAhgv8lF7
bnvJOl2UBsfXGhHDb18SBgls8HvMMcHOKt9wJRlDbeu3q3/kqRIxJduRnwjRR+FchYToM06I+q0C
qDxUBzJMF3VjuhhR3gAGv0+BwZzvX0Qs2vyB9hOOr67KnvfIFJBB07RaamJryigrltRbQ3myYrzH
5qRe8jkqWYK2jcGRDO2M5ABY8Z3ZwoxwMxGDSrgxY8LnlSmud3PGjOpK3OgMNaXFQvwDBL0h3QXG
rMrkNQOqt+TMOtF+sxoqtbQkNBhb0ZZgUOcWyr8+TOOH8CRBgP4iKQ/doMrVWRmzPy19bEw4D/ps
PrgZ7meiYoXRCv6vkYOPQ521+3WZ2/9xs29DCg06x2Osxca69VTLJvBbKJO5TYTv0hFjkl4vc9Vt
QNoH7dJX+8ETZjTsm1gDxYfeTvrvqU5BW5/sBP2GupwAQoa0K4YTGKVFNunK+36e6hrzeM+WHhVV
DM8IxbsKCihetVtoZe4ssXZkGDOGm9qupHGyU3tHin9zT/WHH/I6CVyomWnzDlG0DfTxUB1kZTvB
oiSrLvXLL6gXE6dOmVSxwqWD4M8V0j0LeLIk5MzW37F5OU9kV25ozP8nfq/lYr5QAHxFYUglyX98
e7PC63ZmL3kUVBKbMy3nKGzvX7K6tWE20NmQQ8elOgZV7uCnO1oisGJRTozA7eTooVX0hV6Lu7wX
EBqOvMrcV7yWH9+MO8vDlru4h1Y272E89OG33UuM9+AK80CG6G3JU0cVsm6qTvnfoe9eJKZaaAiM
UMZuM1dbsbrMDBlLj56s2kY9QQVipKGCydW5ZugBMkiSXf5kmixyXhpNvN9d4ySmR6RB6EXZgdmi
TrQ8N0yvnq3iQfK7Cv7Yi/vgnAF9HwwLv+nAfEGGA5+lonL0D/VQnWIAZnT1EJBy+bGupeGnygfY
Umeis0KoeZzwSExCuVGcpk4zCaJk65JP3k8uIUj4rPHau8ohxBFRTSfdB+13af44TkQTM5bWSIwc
7UlhYXwBEG/5BXga2OErH1YzIEkacoSSGFXSt8Ov7vbyAEbH0FKS+QGOtQlB3ADeap9NSgk8RLqb
gdHJax2LPqt4uPAAFRJCYRzQ0P598axL1EEPxzxP1JD8JHniLYQVvn0bxEjMTt8HaH2C3RaFPMyX
s2lD1cLcl3w/2jXwzH4MnDOTAIAUf2MTnI9v7RrqRBugVovMSWah4sS/yFPR5021dOvOgr90SHB1
oxTjnenWeGhnI/FxwsC3Vuk62aJMCGjk3IEaaMikAIls1TmBG5lludOsHYoYcIstZeEDby8k3Ldj
x0dBcezj+6H4ET+bAUUXHGKCiCP8N90sY2PGwkl2gmAwF7PIEfkbHSsIhEo0MpBP44v8jkDyjtX9
UOzospN1IWDjggyxGq0wlqTDo7kYEkM6mljTQ+OKwtwm6m1P3yds9gCzQ3Mz3l6mGqxiyVuTxlWn
wZIpgiw8guzRPTWcPHEPQEy75m0hrz/16U+9oB/VSK6OxLHfFtd7UYy97sWW31OJ03KrqkTZfI4/
HG+XKQpWAqJQnMGhSmXhjG0dG8OCJYRtSUhEIdopo0Bn440PZv1aJchFpY/BJl3pDBMu6+03KFpY
duzjv9YzTloE0dmO11ilJh66854DjDf+LYs2lmnMn7kxC+1aUq37LIISdB24KdsBKU1aZNpm6EHE
DZS1wsCpZDZxOcEtwSxMuHcgM8O9LlIUnvLVL7ZEjgCNQC/Acof4DpYn0iYO1gcNRMJHBIcgMGBC
dc4v8kUTHL/MpakB6M3ZERieXUV8y8QapLqauH5K2NwC7KLYtLK5F4OkWmdsfy/8hxd8eUg9yQ1r
Ili8I2RaYne9UovMpAHTdDnKbfnC4Kv200jDU5OB+XqWY3DLIVO6vMz/frZB0cZAgciIuUPlAt9x
TwcIjOZ85NSQ49c2IzYlELO83+MOewRGjTEma2GVn+dEGEdBGVUCEqmkP4uvyLzYh2Iq53AEyPYT
+QGmoUIsuIMUF/PtylVISJ0kuz27zHvneY5at1Nj92VEhGVyJM0kfXAb9Emjo7MpK8+5AmkGfuuT
qojyx0qKjyB79fpikDB0jj3hPxhvYt+OHaSks8TlbK/NDKbFiPtZdzM/k203XygnhTQrX5erwJC3
RRT00qChhPOd/mFAha8xmEEBL44tKU9MaD+HpvZMUHPu7qX7rx7LtxWTdh8rNurxhXCI1QHIwa/W
xOO0lHVCEbk/9PerhTzcwCgsxPY3rMAf3B3dJuE2NuKjeKE6Yb7CQWTNxglpJf8cTjVch92hAsrA
4TEoQ9CmGeWerWVmt0nR6cOycwI1icOqQMYHQL53IwY/cYBdETx/pbUsVT/hbB03az4rGuqfBVTF
IL02VeH4HtQ6U2ibgPuRTJfBrv45F/87Ybj6Ro6Fkc4MmuUk0qUeh+QUsc3ZxdvyWuwdt1RDBwXr
VA/DyDicJSQz62dQBiKFKt/BJ63IQk0R0713PxdIH/WDJeidvO0EoEL+/OTP0sU7kRXylsPsAYEj
WW8j2GQ/URNh3mL+B4KG7RPWmQ5BvQv38wMVA4HTw7AlGx+VSCSpAP1K6wcedqduL+ZYEO0VfhLe
L+vIS0pS2PpMf/B0G5r1oeiui8qrc7CyCuaf3bRxd34l4BL6dRQJpscxemOtg4xK8IGVa+CCfhGT
xww2CxECF2YJ+8jELPqpj6GiDJ9pH8zqou9ryInR/D707cR28Mi3q4Y27q2g0TyXqeYy+OAsl3IS
zcy7QZJ8qWE6Hd44MzzbhLV+kWXajKR1PkbiuxA+SziJJy4s1m/67y/97X64vCFY6b5Lc2lMsqFQ
UMOA5jIKPOCdhoLrf7y/zknEXLjDnsyz39zzXprygVSH/oYjaAsHNxuL4oPwYrQ/2OICmiZc2WsX
pCamyTgMXMdpGj5i1Mj1pEMTDVEsfNEN1zf8pQPVyqPvPe8rR7SvmTtWCHB/5JOEUPNvUFqnI9Qe
78DZnH0qV0Gml8nL4xn7NkZnaRfJBhq+x/WozO/U0xyft4A6lNqlLM4MnNfdnuvjfIeSYiBN6I3/
hVJPqulV8mmpVKd0GvtMUA/jd7GHOXlEjSTpTjMYx+cO4bFZRT+GP1Fb2qCpFrtAhfKLGovV7vYg
CLj6ntTWwdt52NLIOTfmH6KZckeVEBVjUpqsFvvXUSGH8GczD+3E81K5a6dBOvNLrfU2AbhZpczr
jaFNlfITURGiVg5x2/7cJqmoNW+XirPPxeBOiQnt6wzf8lrgOILHcCRHLUk0ENx51ReDufrcgIXR
tMz8JwVgqViWjJAk/3g6f67KOj6cLkJbhnUDexelIf/bMZ/2DiiX12RncpVdFFjd2qet+ReewjJ7
yjPFhuJU/yYJt6tHPedRzFHWnzTrkk2qefqXiHQEK+Zp37V3RwiEQJL1AtbYvC3lZnmqrT9BDf5a
ms9PDI8OZ/U2yEO40XhwYgAVpyKqdpPgpsOOJ25eP/uses7J6C1dxoa45ScBIBOscea5VRWaX2iR
URwsW9YbaAhIMLQGsmDOp7aKWGVwhJ0G4JNzgoteleUva3b3lBgavaGM0vKYtNON31h+3Rt3TXBa
Za5w86wQOc86OANC8AFJQG9r7ofSzkWMLJrhojpsFyTRJLo9/WOu4DtisOzqfrlJgpazW8yIa9RM
+6get6Q7SRADlN9lAH41Sh6pWlSi0TqZvy7xfp1WogSTu3Er0IYRkho85lA1WpaTV8ajsCs0WN5U
1lRAzgrxz8vnzcB+eolQOyr6QP2uejUXwFe9gC6r6UY5GATDhCuL8KmFPY/RVfqHAFrntjUHZlvM
xYxNyazpZJ0CJqCCH9KmdqrmXdrL5fZPQeNQBbKsBTfcXbysLRp8V8NQG33xIrwDUw1dusGPr8Y+
lp7xJ0jfB9rQ4pz6rroWd9b41NjV9JOQ5jvoApsk8ok7gZ9ZEXAR5HZheLRxblz1o/9/pJaNEi9m
Te8T0EH3uIkuR4uXr53t07Fp5SKG9tF+0WrhgsGMq1+VDy6CG0ojJlQkG2lH/jvWB/7PaB/leUfm
CUACrWbAjh9UK8QhTmRYh+lQXJ51ekRUf1J/fLvLRm8kkhqLuek7RuCIQAlezaxrPq6N7uK5XcWq
KxH8KB0hajvl3htRNGSFa4FOtW4GFst222ZS7fI/TQ5t9b211kTGgj44AftBwXXf+eJRRta5ZiiZ
nTi/5mskyVZ9dbDDNVZC3L55OatiZF1kuvgdsperYNX9O1lKnQB8+q7fIozIqnbR4cpSv/llSHeZ
EOjczOINnGk+y2LthYA9/W/REnyy5U9i32wsZQwVI4ZJjDtsjau2XvAlfZlHl0dgGb7lZonKaBaL
QpgynrqtAlE4PBH0hygqyGSNoKbeFY6dJDKWg0HQcJasvHopRGCFn7BBN1JwGn++XaxIbjOR9Ta1
H4mhl/nquEnr33VH+zCqYDOJsIRSdkafLA/8g8gXu6veY34p1qYhR2sARXDRe6OYsDWpEnK+vp2c
2OIxPnVwoLuGauH1xF95XW2VChdrCEiIb5BIJkSKZQ3WWUSX/ZzUx9Zc1fEoIhxX4dw9oxhDn7Nw
xHWa2LKjpTCaKNBU8ggYTssrky9ZGFx16pTvJzSSMB18B379e6doq0ELr87qu8K9FoTzMSzipy6G
pEZc8V1G4Nz/2M1dPKb2uLSnfobnBbfOHEi1HkVY2knZATjsaTJFsptFJmaJyyISNTe+72fS7kyY
bZRWnwj2Cz3c8SYC6k8BsZ+Srx+YgrUwjRjNryv/8DNuGIbAY87XNgXl/aPLVU+a5pqcvjsqGvAi
DTjOkTU0FylyvCZiJrekrs7lzqKj1gZp0+BizxWEMeDjtrC7dcIj9tLvYbObZHFaWp3Zmrh9pnSV
sX2I3VLTOoYuWYesXMPFUC7khwEkW+ctYQ7CMDZOi4+QKgaIze7/D8n/+zfg0WRfogDQYQ5dtftA
Qp43H32ZHb+W3jLfuksfSmVgHUSq66PnC3gw652g+OFFwslvx08dShyV8Kbe/QZ4ocKZjl/39DaT
QvLIsU8bVbl1Qb7LWmRQ5Y/3IZE/kzMGmIA4YTEO0KPa6DpGQZfxBLWGRy9UbA8L5is7QH7/WUtD
FSHorWnDPOd6a2FsG7PYzwWRjH9Vl8sVOzbD2iRxqy/xy0nOvoYzAhPI03pKqtW6HqFUwDidsYMi
NJk6eL8OLeUgD1n35mJDpzkfNhN0EKPMb/Sm+MHDIoR83KMR+dclDswL1+cujOc78stDN4I1zuJI
DzLJrgJg/eBrCcjQ8Hj8/KGTBejAz72ShUd+E+A2e4dMdzVUM56MW6MrxFJkPCTyjZ5PkYx1pewV
sfDX+xhmItrNn2Z20vIxEhIk1jugZ5zcBJU0mpScOkaIdtq7/IP5D/vhKVFnJ91QaEiRR9hbUHox
7TPWSTF2CblHJyoeS/gGtcedUGONGn9UlM05lv82HpIcQY1El9HXwJzRWO1QkMGlIs/PVZbnIh45
OL03oc+bKO8IkYV0L7ONRmbpaC1DEIDeh18SzjMLwnwjFxs9dPogU07USdg289DOmpxjqj87V2Cu
4Iu03i9lV/POfUirTUN6SLgKPgZjy35+dwYOUBtIQBosIrs/gA88FENIwRj12p/V3Nr97VJM25XS
I6xT7+EB/I33M/OzZzvVrBxbC/9vU7G2P8e7F3LTo020FLWwrh+tF82IiLhpMh/tkKBMRwBij8pd
altvxBysvCCeRDOGb0vjUxBE+/WLwLlC92IIt6/b8jG9gLRwtnqgge7goticzAHUlu0ROp+euKlW
X0kQdqLri9HeEfgesWqxFgUHFqh62WNGGTlVie7/1DNO8iDxR66KPfcsu4J0drV2BA68gLk9J2/3
YFlBuwXBA4jl8AZ6++qF+EV2wOHkG4pwS0dRLdv01otbLwE7aIkRr3E5T77qoOdhuuWcFfX6K/EA
m9ek8//BNrJMrd4z7T6kqTM/oIAy8Jonv2DSbTgfR8M3q3/1KgEGZHz2SlVnrCydAHVHfELYaAq2
Ova13sfJIYArgS+UjP8EkZxiJTu5sbtY9V4gBVOGuE4FgEV1IMKQARm+QmLSWhPZN68TAVvW3wi7
YzQbrqI9oeQUcx4bdLrqiftO/8t876NDOXAxQmiEvWmLsV5ofpO3WFcpXGDk1zLKsIJ5BLN67tjv
0ACmyn4H3+aAKdzgAGL8Zr8VOc/oDROmd6uDHWHjvJf+Kd1DZYYQgiNwn1qgLc+kd5puA0MsLhZQ
68NmNKrc2uVKnu1yCfqnoP/TAVqULOB0rO2plXlcnyHom8kwFoxW7hy3dOWN2VX8A46WYC1MsI2j
Gx2Y5SfbqrH346+g6swEldxY/XS1HRIJ807hLUBa4rpJ0GhWrCyiBylOVQHQcKiV8q9zcCqaDg7s
ySCVg0RB9Ouz4Fq4XYloh0egIA7is4GdmHbCudnrGiouE8l1d7xxCpz3XfciLwXoWssLjgP4JM2Q
3Jl4xWN0Ur++dkVO0xQRziGGTAKYf0QB0zX7hYSo3ZDPYUTKFolqW+NWS0+aaez8usKdghoxjXdH
fT470zWidXMeHuKyrqMhRrwtJKKmxwRmS0s1OGbdIpI1oORcm6PXwewIeW2JYDsjznN78Xui0LLk
/iayp9WosvfS4/UMnviagavRA85dSDvNhhScDCXJi8cDhqD6K+IA2bBnhNLzKEBtY4rTunshHzVK
xh81bgOAwjsjAc3cmSIfvFk/vaoaMpP3Yli+XvPCSySaH9ldUv8hhiP6i/p1XhnM3ywGwhlYM3Nl
ZWtBWv3DrUsrdbj9YxCeWcBdLA/AdVpv6pbILza/ha0/3tVhOBJd22Woa2tezOnFLw2kLNuftg6L
TmcmcD2d0JzSUg0Taoga5S/GZuSwbTmAIxrFujKHGNDVvpS2Gl0pGAraMNfxCS96okwmqHss0XJo
uhywhECUw9kZH8IzdmH4bJ38fzJE9fbyezy0FC6aILRgvOf2JxriI6+vtldm9eZovY4cxMRLVWXs
aSGwaq6CZQFgkbb2lTahDqCdDeXpv+nRPzIGbTwng97ZOUy7dcNvFYldXSb3svpzgfr3pJdiOFkF
qjfuokwwjorEWPFMLEvdfN5m81kFN+xDP1tIOq7ChmZIwUuhNwSQVWGcKYDhlsfsBHt5IFlmssbQ
74T0OQk9K1YshOj758oTcEuEpMiQpLOPYsaoVwRqSV4Tq52lrmUerhZUC2SakEmsogeDPH+GGOj2
P0bCG1iX7MobhHR+gCMnpenY+g5xlTXYImxIyb8g71Ptee4TOKFGYzWjEDtwX4aunZ6l4fIGrAOp
9xI33X21tJYDKQ2U7mzjaKveqtoMgP5BnvLSKlbSjkZXpUWIbCnmWe13PD0Ru7+UfhAwcRMtLwkI
2HCCPyFzhNmay36COIyQFwczHfJvDaZwJrazEw20YxMCdi9KNs1m/1d1CB+7QleqTMWe7AhSoB7u
9ETRa0bxq9OjzbPFqY/lqzztqvoZKS1pUIfQG11opsD4RTOWAkAcAezZZFseHKpf0GOPY/HgZzht
S3MMNwsEzVl71KGwaWhoY7BOuiGVBaGeaF+O+f5U31bGc55v1hop4sALs55iFvcDD9DXiid2FXaS
Ok6NI3lv7B9+rAEalXpM/ueAfEeFGOJC9JQT2X7o9PQjIQF6WSpLicggU6Ew9S5SqU4wk9+v0ie4
pR58eyZwCeRXkGHwfQyFlYciwn8G2bgbAyt4lDfXe6E/TTgzBYQIURV+KjxqkqNEP7HMyxmG7Tj5
JdNdWUpA04bHHs35X+IeViMy1ylZa9zJxlsnv9hwVSAwT4yKJVI8YJ8T78UrLKk/BmG2Ti8K1wg0
ATDgE+vwbxGImWyf7Dm2Fkbdr+sLr6xD0EAVWyUQg11cHIjNEZpxI2OZfoCSKpA7W66mXfwlhEsO
9z+l80BAzSeEE7ASGfL+CZ5NOGSLqyX62HOgTaP+5+8JOb82x00h5mrUpiub6tRjdrtn/37jp7Ha
g6nbR/q7fZlXmeopwaSCseDDXM30H9ihwT+W3t9Bt40W2wB2Eu7mQA7HsQigzUUp/KBUxyv8CMU8
qkNjbOudeEa7hHj5asC7FBF1hL3AemWS2tKSgTHiUzUkp6G4hT290WSaeP4UlCFvAYIRMCj7u8PP
rSim68+SQFw42HtaXYIf26gJbzo3Zn+8irTpfT9Ugrysw4yXU3n8D1nW/8p+6ozgT53ysgr8JQJ3
hp3ACcXm+hMO6rSR7SCHFfGto+XYxx7iyJvG2QH1bfb9Eu+3FGx+bsR6ISSHLDfveFWkq8ZTtlLM
Ht1TAREJbVFrCEjEOb0mdnEFQJyJmtQLdurQYz1w2i4b/skYcq+ipEsr4oFzlDt5rJWih7S5Aqya
UJyUqZ3zJTvdVcVRGHV+lyN5N4lGPl2Vl0wfa//Z9nMgvfH5pO4Zwv+eK4lK8aVTM5QZE1KHgDww
TvUwLFy0O9gzSEtNH9DEgVGe4R02hE8j9vg20oQ117lv2dPjx7P9uM4CNKxXtrvN9W/FETxPoKFw
ul/z3r5pO/bxDNg5P3b6EQin0khxWOoHLG2Z8b8RDNZrzxc+CuzyLKnYl0pkgaXHfh4Gj6GUxGdD
nrlhVUG6XmQPlFxq+dh28pJDL7Qt6YjhQbEk70bq4dATEBzHsWAM2D49A+AmDrkcnnNoQhUO2IcU
M9S8dTNOSdV2bIf5eCuaGtx+osXq0s5i1wMAyO7xU66PHoEs6FSCWkuonaab21aNeMUBvgihk7JC
SqKv8fI7epzgTJU5JEcfJc+ETIii3XWo+UYrbuXsIGfp2gr/6KHf9hxzxIOCSL26bTovlXN88RAZ
yort10ituy9roJRjKLuKuBQoeApjBDkzrRILWplEMHFT+Ndf2VR0z7k3CnH4Wh/13TD4D/FDsUJA
7l4OMVDC+XC9WtLMbDBi34VgClhnO4fJr4qpN5HqTZyLGSOPbolsSKHvqbH6hsw0DcAeD+YerjrL
yO2BX72LdC71+GALOe/wMmBMV3WVAwB4lrhyUYwgnJYrCHtYIb0Dv7pQEUz4m8StK5zjwLcXJGbv
YtkQTriMahPt0KjSpc1/sa4YhuEo04BGZOjbBeSir/sB+4n4wmOAtX2YboEk3CIX0zcSTDWizgKl
EqdEhOgodWYTii7FzhCIqb0tVQntPyvoO/UOt353AE9DlT0jjb+Rqi1eyKXaYzK24LTjd9yeGHI9
V97Sas3PPS+KvgDYRVA0jLRzYwotb/dXLhE+tK+fr/8PRxU1aYVV3oE12u/UGlrGRHA0Vchycfwg
Kc+J1XLZ4kLrcAeupbLiM8ChUKEe8/PXTB69KsQPsg9etTb6l6V9OksDfKHedRNzBf1Nz6IyvsWj
I5878Ld9Ohyp14ym/AVy4rNpNTKpgTtweDeWUXpqk9FMAW5NWJeIbRDnfsu1HaFc2hvPmtdjQH+g
aZwdkBmua43FCov8rZhggR+mRnbIp2fmzMJC1MpM9EFXbYRpauHG01OQyCMjgJTeiyf6Um0biRgj
K7QJm9YmJFGFtkvh8+H3SHliksYsLSRMW2mX+TBd8ykIo4LXNlCqKuTx+fqz+mpT6Ir46L3hQQt8
5Jf7UlWjF7WD2t428qE/HZSMrsBHEqG/ezz22udE1jauJMjBBpz+OvEkqCuFuX2syPuN97cMrZXM
OBNgiDQrniLRIxPow5+YY/KwxzCBqdBVc5kpUYGVshIpi6XRUyffHF6+2sALOlV0QobPofh3BXiM
FwW2rdQXNyTKe075GFMWrD1xe3lAJNX331STuwKrLL+8R1XGTKfA92ri2mzNjilkY2d/nbnx7GBD
QsQDu/ycdEAhKzEpqrIvmAMBFK/75dstAxwiwSWvgPPrpPRYXT+fAcoiECV05Kal7bkMP1lvmQEa
mcBjAtBDEI1JjvRPcFpI1wqyH4pN43gZRnR4WNhQ2inDlBsR3A75W+wzgIH3I+LMIuoYps8SDp9r
/CnF772ZDhIDfADqkxU7OQ8qFhn9NVnUOIEYX/dugfHz8R2Z33PYmTy/uVE1Y6Zv4e+36KqXpUWB
u6xtDfJiPOLdxhXN+VarQsLXXwG64zHsMRdyC2tyXPGFlLimt9a5ngkbPGjMGABZnyfhqLsvVtPh
HBI92JXP8b1cOAy7Jovxd+LCMY/bVxhHS9nyP20gAIKD6TvYj7spkt5OKSIJEIHNsUUR9dBMz+C8
yN3dgXM4/Z2PUhICz7SpT0hOmNIBr088GWv6z32Y1683opLqLqVQEnYlMlV9uQzn9GFblRE0Kf6r
NsI1fTMtapYsZd7TYp+G67qCblf4zPTHJ8kQUH1nogu0s7kKKYiqGY7/GDn1zIODKjAYcoKK+sAE
zG3xPLN+p5dIVQgwyZeACnkIx6YXyefyEp3q74TG6+sX7q3bajKSbkWDG0XLmy780BV+a/CS+KcT
CpTdlUOBNrOncC9jmR49YUS6vRWZFkMVTVYpoaN8Hbl8JPImq6r4Zum8F7WNvwQG+6rtoQJewQ0D
sf6hZXoaqFIAtjiHpPzUKHyZCLjvGQF65qYywujgxJ1YyD/jZcu+9Ztpw30sATSYysP4z1aiX1sp
+7ZQdnOFPzg3axjknZGqHaXgGKcT25iBn8MwypAYxkCgYwPWVqnlHF2ac+1sZdy0XcCpF6AlfUs9
Ket8l+utFXEu0OHrNBiRlWyen0bfP8/Te1gejM7d+48rXCbJAya1LT+GcXhBg5Feo684wgm+q5H0
w/Al1gdtxDAA+pWqKWNZCxu7gx5XmxVzfe2hdBG9S8lHlrjHZuziMXzaeKyUyYEsyFFqJgg+AOG2
Y1zsHcs5qiWtxm1YzrDGAcWJWhv35PbW7CEU3ny/rpfz+mA6jxILHigvhADwktT6tPzZpS4oWT2k
qSgrC9AQ2okTF3kSCgKecypk5xymskoroVuLst4FRT91wWVKSozVg7H0r6WNLrn1zj2TthqpwrM7
asWGx/Q2Eo6dmu96GVF7Juvxfafs317K+AFhkBI8T897kUX3EWosulOJPeY01W6JVLhasWmHHat9
0+RxwR6eqKZdhhkKdYNWboITwKBwQZDqfAFy909AniFzo0DVv8UlF449e8S8xdi+phlpdjGUrhvj
8Uzuc86O/96KSrAsk3Ue7XGuD3KxvKMwTsqRDbl7rsoYhoi5Go2rRJcb6GaUpnoJhzc9ZitEyf7X
bALlo9AlkisXtmW0gRsS6IQz+2/3Nwj7gqhEPeX1FekI5wwUQ/ld6S2ChctXWLbDs6erc3l99IGJ
MP7Nov9SBjhjC1yJEy8W622GshiYgywkR1+htSpECPqC4tllPHh+pZdF5AaDLwqTTK93e2KUok3F
qh/EY1E+30t1ZHqcpU+aIKWvDbxZaPC0f0gzVHmYbLXlMsym/xPiwA8xn10fguZ5SFOoGp8nOz71
13ql8IVbfkoGbWW+wiRzcFm2ClShi/xNdi4abPLT49O/nVjXdMDFUHCsHfwuWjJYLYUa4ulWyHUT
q+GCFuXJA9ZlZOd9d1KEW1/0q4kiknZNsm7geytZA37slnExfXBpjVRA7XlxCOZpG6/QQJT/RBIq
K6M214N76pqNx/QGz2CWry5cpsMFWJS3fUwsJ1cuaPt58vHtYV6aLKTqFYsudc57QV2dj15ft9/e
27gsXvzB3VQ2MUQFhqIciORNmoLbEVh0PnZz6WaxY4GAOVwRhYrLYDAq4V14X8KC2F1RnpFdVmA0
V2TQI/tg6pupj5AF3TKZI0y3gL7dLGNp7fcH6utMtf1fBJRp1iMBb/s08Y09xiKc863ddVn+vpAy
tPszhVlQMzZOxKaHB8wyh8tPzLypXsyJO5yU3c1Ez7T1GSr56gNyDhKcdecuqf27nI5oRdqCnuCW
25CxIU8Rj+aumqjiN8O8vg3+ML3ewxXHJeUHA/3Xfk/ix72qI4GA8pBs7zKKFKiZuhcD0xMCND9R
Dy+1I9eHQacfCzSEUxahnKsbU372Xn1lsa/K48hq80G1Up+eutSdKVnh606CQ6hC5EvcRFfwsNh4
N+ThNqQXoOK3lNGceRL/F1IMn0WyBlBGJwZ5sDAa/zVPq1jPJn1plbCfNHmJ7qIs2/RvhxKU8tgP
8fsptVILO7PN5GJCz8QyssT74vppqi7XWXMKrM6P+tf5hw8U/eRr6Lf7loG7FjcahCiA9t+XVtgD
+yUQOH0Tg/ydUIH8wOXPMMgxnPNdSY/hRT2Ydj+aEugdgfxmgFUlwZj6FtNLsFUXedtgGyqOOm1p
JwinZpKoVyugeCUH6bEeFjnURoZZZEGA48I+zBzt3EjihpPUL9OqUI3f5JENc/i1eqBSX5z6uREV
UuV1cY5nhAgzwRnVZbVw8Q/GTHZdGKr5Hgm5x10EvsONfLSRqCmJqrFewUTUVblLfrrps1GiDPQE
5OJLz68bhK1QG38UUo9BAIKlhPmLedkvJcdOIXLycpMqPefeE3RRv2yy8D7hqzYug7N1uKk2cAJF
uPkXucWEp9okqnVcOwUbNFTj+BaEHJTHwiEmV85xiiTftQAN2sycHaK2TCANrpjD7wVKbT7e9Lqf
t2XUJGirQeu4YhEnZlTzDlcYcTaTJxW61fDyR5OWVn+o443l9iciEF4nWJgaE4UDyNA9qooLo3ux
LPUrnKZS/T54YtAg7ErP8SsThmgokGMefxn9xPU5O3dgNxyrJ4/KEJA2xO4K10dXq6QEnrxlTfO5
3QHM9TgPiRuXS4NWU22ZNh0ee7gC+JN+U0XuROJ2dJTFgU/stwjXVVcq7Tqtn2REb3/Wv1r57SlQ
628c+Gr10akpK2CrTlJcBCwOvZNjrUEvaPCSScc9gyEg5ysboEuOOI4ePA8bcEqpoWk1vkR15zff
gX8HTAu/0hliOxNDuX41avpi9FsnFmniJwNVju05W+NeIEjp7Z/Tz5PgmCIU34DW/M6S/GGRn+Zp
Fd9g4uQ2c0jpCX8yMok8MGGIkqsuBbqJSWvmc3+kxyZYeUTAMWT+LCL33fqBcUsOtVagWHBhyALO
+1FGHCiRh7KdVNvgupO2RNQCpU31vGc0abSXXIJa+Kdp4nllH1wxQBBhOGkDu3xBsejCcH2mVf9u
HwQEwIz1IoIJqWXJ9y8UGIqe45DS9C1/1HADInbFIWMPjN8kOXdOAh321Kg9l5Q/WoNgRaA82wus
A88Iw2KlKlSQvtm4p60mN//sPTYeLZQD4u/7OohqUQK1IyNn8iYAkmPt78nZa4jJC9ekGZoooc6/
IqkP5llHX7hMOUCp8PXAstYOsXelK6AlCUwRpdJeGCUGRoAzMiVJBC37OJTRJZicmM16lo5OdGh/
RwaKNNsbbU4qRRwfYJKo1E9RAXGnlTYQ70mLs4SX6bqeyIdSyPhN3xC2c7WajA/mBhERCOd3GIVG
5QhueMpVLwib+n3Ncn9QiTFz4lmpnsM7JSeFmwvlf6imtqLR4kR1jacHwhP/mc/H4MKFoPKG2XGq
kCie0MEdqxg5MbGu64w/ZhTa4LGHbaYF0eWsRYNVlkxw8KFVJh+vcCaSN7I8BHGt6s65NidmKF/2
Es0oxb3ANo0SfGcJwhXorQdErjPsYnA2awSn9SyY/a7NPHgeFCX21HLoxjiU499z7WZTK7bnbxMI
bUm1Rso14PcwTch4z2RpvIi2jtiXdq0zdHJfJK/b3sYd2H84kNiCRu/70hy1pG1mqHktnVhBkXbK
eXg3ksisKlnZdVTq3Ww2BkswUcWi08dSwG9PdWbP2nmVChTxpPvyq21oH0CXzW7cD56EV/XjMwEo
/Y9gmBFphHufJzis0duW24Nz3846pYW60PLcAIgYAWUbQ/N+JaEercWgtdEXC5O25Fqm7BXtT21S
Im6JNsXabWJwLYxnEdIoYq+lKAVtFUfUK784yZPXBry3qUe14oKWLCau3rzEhCyylx6ELBP7XwS7
0j6jlKUnw5MBb2D5maRIxh4jDUbpFUSUNVi2KtII5gjoMcxoYwAlyZbLJ9cn5SSJQRW8I4as9miM
3P7hLDqhYS0wuWW4kXv129ecDqWjOm1Grf44t2w02bdULbNPjREHiOEr8I9bghzTsTxKRxc41uZL
CmxHV8r4OEPwch2vMiVom8QssYPVKZ1cX59RIMcR81MbjuBjYH5Mt0ywP/o5sKrc930ZLA0P8LeN
YEM1Xd63oVKvLogu+/Oa/HPDfOdtytZPFvuLRtihVAp/uZfzNzNbU62EntZmwn67we8ooX03T4QB
ZIlo4QHC8zXMDw/1uGYg9x6LUwQf9E+2YFqyCrNiqJqhqcBfBaJRUKierP+P0RAfAdpPaQqw6opx
2WRKMlUSufZ3Ys27NikdXBJ7xy3WEGGA+d8g7e8OKo7cxglxPMHFVEI+hAw2z9U/zj+Qg8REDxQ2
vClTVWHs8xHgyfK7l7s3MG/dIFCs2Gnc5W2Z1H8+kZkBz/EVxOiwanCaO0M9obmoIjYrUFhd4THi
2ZzrNfuBAscj2/w3pyamxwATkPyyStoQ4iJYHJziEhye3gSPHNgMnTR0QwuCmlPE+jkHwfNDVjvq
HJPkxgz+psxFv3izSucnbJmrU2XPrvQlQeQ8k95ALZ2K7uB+mBmlOJ2+Kb3k2cej4/OI/QLQHJ5a
skcAo2lvFt+/OGMB/027EsdiY71WK6/OZ85blFU/z6qwoSsj/6sMbtUtTZimq/rQD8kwA2naJn59
vUbHGpQcjEM12ejDQDDZjnyCQaBvEFfSCiROHfZGhbnYvuIBKgSfHgo+XLhpU0rfcecFVA1DqyHu
uBRdm+dSHJNzHeHyvCn1z85SKgr5B6m0tDh4JuaUiENfxr1DEbF5ZFJtS7Chaj86Dx/c/z3ET0Z9
uYhJIud3qa7tCZn7Tgr2wOl/mtEYXXNZic0iDjV+EBqPlz8eSL0JojVPWZBAkAsjUoY+EDhPPbV6
GdNt5vXvVBOSM/+KUwGMmYDkYD0a0AthwJHG3BmnSvOxAvV3Kc2Uqnjz/VkTXt8XaJ/MQP0Z8O6P
9hBnNk1ugEtDjGOWMZE4OnO5C/MY1P8/jX0pJyk3ZcqHVLO0zQJX7Z0995cgoYZkMJfIFScu/9Er
DQiFZR22rRarf498MqQOu40xhpMraDmYcSGOF8vuoc4rLz7f/RamARBL5IcbpUfl/wJuQ2id8QMJ
/Gy0v8+twZi1M53RA/do6RqOLLUVlDAj98pZpS+1Zz6J9aJzK2QUKYYi01I73JLT6EzsT84zJ1fJ
6ZjdwGfdRXMBZhzyI5RwaomtD4yUpHIMwZA80gP/vhTLCscQ/N6YvUXIXm+eDFArfFldZVI8FRAE
/jZr2HSgznyBW7Tbz/hZhIR+ZTAJUnF82VdB044iePV5WDU6tgSN6hVC1mk4uOqNPM4CJrJa4Xu8
DgtElSRnmHR8DobkFzU7UeYcLVax2NumAJfuqPWSxxytuyzZXN36s3Qp0Ae/amCxtHPDqwUcbrwQ
h2QLyf1P5Ac2XzlYk5oRgXaLNqR+LJ079U62Y6PwX4KrStVsZgaaAbyKwvkxFkJQOIeeEhLFswKt
EBd9yb85401cSXxpsprKUwVVbmOEjP/pWBb4LHgGs9M1mV06BbCap87EbaY1uaFjjzJgWEjCcNb5
VYrERdZaufLSHzhpgVZunZwi7qV/l1ruZj6HYgrXhMVGqp5AxHYvflBwtGSnKd/kZMpiowaMWX3d
NhsA8/NwMJAWayG53PzchUMbzlX40zPku/QRiC9IpyxuwElRAX8u4aFvyRYc1gEIblH9mIdQNsXQ
bDzqL19Uis6PWNFg8TkvlVcReRC3BYxZZZpLgbYZcIb9moFVo+I9aETC6LfSMTHegk/6xJgVgzsa
qp/3ZDwxkeQN79t7W1qG8FwA9x2tZ6xaHTZrpekL1qxzOWfNVEvc88pAQjZXX7LO9rBfjWhNuI04
ieDEr+HVfgu4D2eMMh081lH+WLNMf5MKisU+is0gYEOIoAh7YkF1mFcfo49F3mJ0MwihKdXc9TDE
W44Yjts+5FLzOa0mUn6X/r5o+aLuBgK5OprDwjfL+aWoBByEov+dI/awAfVfYoOuGifF3E1i8h0w
JaXp60ysK5SQk67X+QhCpeqynoy91GUSjZNDXB1OzNEd3PQTbL2vXwW1mvDnqmFVJJkZbsHkwSA0
UWw6iMbbJM2Nym+cgtP7mwDQMwcQKgNgdVvf+13wrXdkjQWjcx9vPx9E5eApEEcHBImN5JZA1xe9
qOKUOJvU69fqBw/e7kZ5INuZF6cPIh87kwovjx/trJZ/MDjubyKSsNZIByK+CFAGUMA8YXUURsp2
1l3QEBmkVEIN4tIWlKHC/jmmXzP/BdqvUN8nkPp7f8JXJ9PsjV3myRLvM/AxjaKqn8hOELd0O1W1
ZFbUwdCk9Z/g4WHbwQrry+rhxV+aNtvAIf5sS8d6s5PoOe+wxN9Q24lhb1MVsGFgQ7KxJWzPigUa
dKbFRKatAzJyaNeswbs+udrEPTwT1A31H2MUrDP5SLE5VFqg2/tHnkGXgl8u7qbDSp3/TaqMSMIM
heqa1EYa1+QfTAw9AkfLIse/6IT6DWy/UsNXVS3I+mSVqGVAfrS+18+EdMIBjnTiKgbIb2svGkUw
rNJWb7BoTnYgz3eMmJixZrabnRDJFkWMCDxnElt9AGC5Ms+yR55SDH/ftbkhBlVj519CJf+Yqp2d
wKUnu9lUytpIL727cCB/YLP2G/CZ3jqHxo/JpKLHz54O3WW+3Pg8ldz3GioVhLqg8LuZy6BGqaqL
keNeGRYGGZmHAfB0AtHwq0SvvIkw+d2bazHod6EI1ysUGeXKKanRZFgFKe5+Y9/KfN9D/s0GmDr/
aLc/+G4LUc4AIBJYT1PizNNS4cSwJm23iWFzhnDjDUn6vH4NE9QImOo8khgxTKWPkgFv9x1y4z+6
aUG1PNZSRCyeFa1n10f0RTt2FpEk34z5h/em0GciOqoNvmXTv+VFxPg4Xxx7RFSs7HWN8+NHIXek
OJ/It8nYOt/S2G4tKbG5M+AIOuUgZOfe7g6dC0z9sp86k027LaQNTvee5NvBXtqxQ0Bh3wbryBH8
pExW4028xHk4f5DSEcqM1m5eQetZ5imXWVVtG18f/kM38kqkMBbu8s2gL/D7NaXRG1KWU7mpipYo
2Fb9GheY7OHRLtG8KoXpQPm94HAQYImrUu0LZcDtc6NP6FmVeoy5VVtgj4u/RJjLL7/nKsJ8zPaY
7I9vqavZR5hRIWyLw/C3cUAxGC7ziPKlP1GMD6kO3W0jIpu3H/5tDh42AyHfUnNrlZVHodfyXOZP
PT79LnnVl1FOlcqBv9mlsQDhujtS7Pv+w06fh527OYiqZvWnaf0Krjw+V3jNqiOPBHDIgxPlLeOI
aHBsjgIZJK/F+2Ab/AUFoRj+r2hhjydUOdP1WANjsiCagVdxxiLIDu2a+7a4HA6Kgb3KGasSJLYa
7pNmJu8y4jJPZI2coVknhJ0fm9SqSxdHYwAtmsQm3vJQ356mahgG/IEr8RF6NuACaV7+955gunE/
rg4W8fLVaxqAb2tB5oH/E72SuQvDF62+Y2OkmGPMm0nSyJOfBrsD2W6FURvRZtIaQLEB9vwEDLS4
xGfSsEHUSAMJskaNI5dyHKpcs61T2D+eTFYZ6dpXeu0l5TKeXw4DFcQUU6U8bGFff5mHUq13qXqd
kASl6e7ukpZzyZ4+ZZkQ5jHj+XcQKn1aEI1cJUQG6iNkVBqeevHJjqJ0SN/14w94TQFk9wrXQ5jE
FpQe+3pcpd9HagS2F+xIFhQXlqr5oAUD68aZhHPxJp4FYaDK7+qEw+v12VjhR3mrSidXR3yMmM5Y
l6k0e/pIPy22anR0SbKesIft6OJsNLiIyAb4yr+4X37q2Ak1LG9cajKLsYhSywA6vPUsKwC9hJXp
DtpIOjpE83jmFUOHsSuNb2MRYLUnteTVy42OYU5uJeQ0W1ZkunegW/ocBlAn/3JD69n52MUBSdSf
bvPtkiyJu1ztBX3bbjT+oWHmDQUvsWpaeUdUe5xt5RRQow/1GPLoxM+xPgtkXAbJunYUC9s6EpWq
rLuqtzGm7MpAQOXwme0zWVaS+9IdoT8xcvL50XOtZSeZ3yA9dGkCZYy6Kjmog4pUtsjQZ2nR0A+A
//ow/aIKJ+EnBvm0x2XhKnWAiFjqDnf/b4xBvRsfIhLucLQXbGfjeXwI84gEIj7WyRQrUhlPAfWW
IA4nOSB0PWcIEJ+lRxF5l7PE3Bf3+gootPBWdNYX/bPoxQfNiO6MX01L0GhkDIwgGexriAXvG0IP
9PC4vxMj4kjyt09E1k6usUUNdAHraWnpwZDRdWnQpytxM7Y9ODklzacbUaXtYbCWpxRq6VT1Az4S
2LvxRDOQjInf75wdAaspgPxpQaeAqzyzNTbEX31AdnpnNT3Z4V2+dAYwTHPVPKNq+5Naan7NkV51
1NidmN+WiEJHAz+YZ7huZY0Tx9I4jAlwoFAeuwpG+uF08g8Eyo4a7MmsWqDLr5r0t/m5KrhdPrGU
tiE0mjdzp++501HJzeGH4VbJMlMsGMr+FggGemJXPgAJZH7hnE2dWLDJq2zNMeYZmwXYNz111OMh
bXjlYpDrxmje8Aj57Z2PNmHbtaeLJoo65IvR+PrhYLIaWOcFufwtTe69D6KbNrWnR5MKjblIngXn
y0y0xDg06l5ZX7w7WyYdjuiqEl6LbrhVubUNQwRvzkKRngbj4KrarP3ymMS+qbEvoQ/HonvF9wMM
X+L+cZwTsXuyHo7hc1cq6kQA8MXPf0SnU4hmQ4xyUZKd7ZS2rFBI9qd1uc07RvvzPqmbqOYr8don
qAU8aYUuUzZ94d2xnfJ1pjT/Y3Q+WxDVmW6/uH908fM6ErtS5kdBkcRrn7wQsGHLg0ZKvIEVdDoR
pOm0tEPwyEw7VxNjiMAx1fIYzOuC9sbHC7l5vftUzbbSthoH91zBCCY3+F5JuEMaeneAvKJ9Cd89
KR+hDG+nxn1onTK3UVqMcWzTKP4IPAnNfaefmL3yC+QMy38o0rdinUISAFg+oQTnw2BAepuqftST
8gqm97iGaVIfqKVwG/WsNX9zsLhKLWDmU71JyCexEOuTlQyoDSwad1qKdVBThDbjrB/U5jksgwYJ
KxZIL0boNHX6W2R7+K1/zzxfuygK4vFWRZj1rgmmZKe7wS9T6Z4cK9pY++x6V5B+XZIqIOxoMc3c
xIumerv6J/eTyHKE8WW69J9ZzjET+Wl+L7yITcjTDbZV7NEinafQzZYAoJKMd1wvfJtit3ZVrPje
x4CYzxa/AUpmMi2ZLYXWnYE2v3icv3B4MuIl6nQ9BFPmKhIeBwZNEuur1C4CGMzS7hf2vttKSAaq
DQkeEBpETr9AgjOS4xLG6UmCISCo2T/jIQIIRKQc3YoaDG/oCvI7qkO5IFpTKviCkM4398UFS2BT
9bGj1ZLHSSesQTB2f3tIJbvOoH/vgV6dZNTm2eLVxx3IsH6nepKlLrp0Yvkdj47EgB6ZRW0z05b8
REjEiOAJcK73BhsjVJYsoKtc85YqUoEnHAEW1b6ILZLClZIA0RG3WGix1WfgQjSVjFOMebTL1XtZ
YVGwQiCR1hJZ/EGU37VM2fd+aFImkeLrN/vuNhMadEl/m7o9dK97WdgjeiP6Va4Pe2CvAW702v5p
alI9c2kJn3qE/QogMhEUNoEqsbU5iT4+yPwoWwVy1o5EsmtuS8+DpIQy2lVa8dA30AkEmISTYtvL
WoqsCJZ6pi8ku+4bAG7COhp0cADupR8F1Asuq5ofRxUewLbzVioqx/y77QbWAjWjbJljc98B4KKH
EVSJHVr2XAtH2igMXLNIGoz/qfc/L+N4bbrhYgi9jhAyeNbeIYamTmLIviAGpTpRPkh+2CB5JSQ8
Th3rY5PCLijReI0YDXK+fVa8CGh8gL6I2VFX5D34CF2hRFtnIgImL0wJLaD4BPmgZmNOF6AON/kV
gilvnZGDwPwyVHkVYKPHlgDEoUTbZCIQ7JTHxFKX/1TZnaE3fsuuN3en2GluoMdv7Fw63NR+BfMG
6Oeu/OIJViDLL9KuVTspgYBe/askFTbyDGuC1g/f11i3pUJuKYC1lFT8xqaalGO6dxqyhZhllDoa
8nFFw5z9CD0aJIB58GMK8KZGFL9xcADbWRzV4llaJE8FWfw64n21P0ax5r64I+9emuYAxXY3GMR6
eKxrdqaOO/ypUOBQE7lCFIoTNoVTs9PHaavpmyfq0q/V94nk1yHU5R/4DNmyhiC3uEhGJSADfZiQ
y6AHqAvZHUI2+4Ixa1psx8uv7tyNbl87b6PZVFfGjCfrZsFHKtQ6HMbFBSaxw0/V2rTgl+IHC2w4
hb4RSRjC5XGHgRfa0j6rPf21BX1dV1s+11RvnI1wmLO9VgouwLobHGd44mE0D18RgGdP0/W9TRlu
e1EyxqblND95Bps6XBmQMwtGAHY92+9pqSt4PcBD9ZUA6LtUNN78MONMTOnGdvUJ4u6MwLlnUKaD
6B6IOC7D06mCbQxf6+0SiOj4+t43x2Ilopte3UEz5nwqyBWz28yHafUpKcHJlCCJHCz6Zr0ntIMN
B8wMnSEfXQGjuIfJNg5kKSQcdQNI7j1GU6vAbsmarY3kCHEszZjQBNhaCkrrnfkjraHegk/SzPRv
fRdiaNOTn7fib3hpf8rKSMXwnwFUza7YXOQEc2Uq1xoff3WpJWLV4cMDzn+gXcV35seSrIId80Tp
tunkCoAMiBqfW0tT/vG/XksZMYZy9z/XvBRRnypSYN+E0hI49UpGA00UUlVzRgXHzTIG7O+GR+I+
SPfxV2ccYB6fZQyuGLYDJc/0VDjaFRuGSzcMKhzP22QywLyjG8DgAZMJ2hV4Y89sd9aO+UUbLQy1
1lipldd8Q+zNzHSS7Du2ieeKBkTZHO3RSCcI74F97wtEo3p+HMgZj1q8fS5pz5BGdG4Yj7fyUOO7
hr3xRZflYZj+bvACle7a4Nc6ORxxtg3csCzWF8lZuZu8vD7CCd4I97sAjME9/C0CUMZ/XLpdKaMK
ff/ojNGdbiHLGCc0v+htlcXLY7TWwLvAWjy5Gsi622JyJIlnOweMXklBYJBo5gql21I7xO+RzkJy
wYnOFEl53VZZVoUnPOz4VBJH4nM/eq89+KZIuHI+61wRK6obiqGyQBM8oeHyX6xEH7kp4LJOYrNn
GMmX7vNlAvSZ+lZFXaP6SMsifulswdbHyPO8a1pqkP0MpNW/USrhCOUHGZIf+F8dN5bQYAbPqAVi
t9eJlEjt6pUoF60+4Lq8AoaSVsPEd1mD5ytGvYUEiWCsH7uxfLqI0iN/HIdAsulwmn1S8OTVFwcO
VFSspjzLFdAFol1WCcEHaISLcURFM5kNqmmu0dEZyqVJSnE3Q3/soH/bLymdYY6Sad3mSLsaJWOr
4fWAL+JKJSnlpcSZxXxXoj9sCs2sBXdiqK7tY0KKa/2Izqx+Xh7rzkk9pDE69allHffx3PMyXNRx
8hFpoFu49sCHGHxO8KtfrhgWVDw/xoxd6O/tk6pK3OoYTbG5bJ78xsfhjv5vCDblAGMPu7OCeHve
av8theiX5QbUbyrbJB4Q1YHfFpDg52XPCa4nPH7/vXULIoga0Znqm1h1TvPsk7yvgC7dvO0aT9A/
DMZjq/9xVwhZOoPupyY0o8Bj7Jq9pzJnNG1L7MZd7mIAivi9VRfU3uZ396MW93FFsHtQIvPy5BZ8
cexwwePj0aWJl1KdvOsbnZzeEXpHI311burQ9jsH4wG8pLQAUaARGPrLyeU2RfrIKtSDU8nXZHyg
e158y9dUczfCTxHP826Llio22E4B8tkz7/ci9JDn/43+WvZ0A7CwfKE935AGJrIIoqRFIhDgq5he
KJFsD2iOJEn7eWnppq6vs/JzO0n6R/sXpwYlrrvO3QiLHK8dQ5PUOmz2Fbdl+eRxqEFQ1IkiP9Xy
jvvxDhp7GGPwhZNiIyFku3RzLNRTUuU3LPq0m2p0JEojkXzo0tw/PdTVPUMTZl9/Uu6moIu1iu8h
86b/6x6yzK0DLB+dtunTYPwxSDGY92wJkoV7vu02kDMH2eUlMLPVmAuSgkHJXo+bWH+OvklCl5yV
K5y1Bcf76ktZz7J1GjWUy+KEHFSS6RLGbKmMMuqgb7Zfv7NlnBGVGKAhNVLZJUzJ74buB6mFDEQB
Ul0OAn8YBWUjjvnptqzlc9nt/CM2I39u7hhaEPb+3psjDqEo1+8JKMz681UimwHfE+Io261U+DO7
kDG079vzWI0tbUpwyXRQBepbiNO8cFWqqcO4vW7hdi1+kYqJU+9d13/0A62phncl4GC4zSUo/2aU
uOwaGgTJcjP0q7wPrFZn6lslk/OhBxcyhuIzjgTP7mbuFnMXDaAT1U9w+N+66Q9ap2X0D6u7/NQ5
MYXaBqOky8SHNkNj/WhDqx7Jk9m12nRp1BW8L50fbhge6DotvV9PwWjS8t6zaAdDg9FAomCvXlGk
qgKUqc7JETOXi4DRfpon6emd64TWDVAIW5LbjllJN+M8njAk7qW0VPMQahuangVMsurzgmvTYJOz
lflOg854AB0QmcEPkcQVWxcl1HnIHNoIDWrlKQmnRD8zJ3pks+2J6B70cHgQazlBCA1NldeYcIMH
5sFJnIbur68edry/HRWE1j2oz8gG0mxqIJiqXsfPfzlFrYcjfHxHdNsr+utCC6ocYkc4tLoLXNb5
LrmIHtzvG21qcvErZUAn3yBtgf8lX2ZHh6MGuAS6YL7v8HzxTcj6fQr0Ge9uhcyK6/p7PYAlPLnY
a+9ZuDe59Qk9Mps6Lq+aUx7kkgbqvHQkJ4m0KTQE5HS7XG4FFevp8SB8EXBvKBO4yXncfzFSC/tG
fOTgiNDvpWh7bmMEnDDHFhnyGHPcH6ahVzcbm4VX3yViXKtKmyHdeJKzvC2ClLo1q/teaEQNGSJf
5nHEtl8yzqHqbm+ntyWwHN0/q961oBiPjwA3rpMmhus0nCu7oSK7wLmNxrEPRriSsul5XWek7TLV
JVPHXtQFiH2rkpMEJpMKW++AJTOemT/OCJgMTe4Nd0BaUBBgUxuRqK/oX9dFVb/9nk0kl+vk9H6e
0eHpQIpJ3IV5IguBd2cKY/uQTksCLeu4U3zrXVZuO9lpDyfdo3vR1+8l6NW/OAI/mxr01XVuGFZj
0HJOe6D4EU08A6FbLIvMFspUS4S7yYeJhzpLY9/0H29Sm3ut5jIhrA6786VR2ePWzbQ2FXC1ewI+
koKNLu2IRgT66rWoCK6CtxzMNUGKUH6ayewtzZS+rApj6lLLsfjeM34qgcQLfxwxnTWjoJ+fFFCa
azPcJI1vP3Aks3j2sVtvGIFRWQHb/t4C9JgslD66bVik5G3liFU7dUy9F+1YqtfmtTBAyiwG4d17
zaZpSxqeu5jUd18tg2OoRYB1mHJ276GJ1w7PuHMVhX0qrU0Fcyb2gElk2ChI3PJgEYloLed/iEeE
7b8tmn+ObIAvdTKgLE1RtAoHvkG1v9PAeuMjHHMAyvymuXUXLOtHATGEnxBnsyDY/eFAiOPjSBMH
Ak4XDGf7yuq4I5dLTWe+HSE/EA8ic9E3TKXqvBnxWJGyTXIZV+m04/9dzzW31z++Z84CyiPm5/et
OcrO0bPgYxZl2S8Vxp+Qmrfennvn/RzoL826fDKkqYME22xC45m4S2gG24pxTOhzLK75LuQ7Af3c
g2AV8XTPH7hnLQPYdAwyRcwZdI1LAqIxLp8L9hsT7UrUJuH02pyRa6ACNG2giluUVVafsCZUIui3
KYYHZgWiiINy+eoeOFuka1zFOkQDj6K+Ku5+IxTv0mkCA0gCDol7p0ky+v2grTfXwK0dXNmuN4SS
XofhGVUawnJAMXFFk9RihmcUsn/jrvb3YusCwwxINALA3xhwa4kSanfg3yV3tw8Nj9HnhC7HeYtv
X8hwgq/Q0bKi82+t7faqTw7BiONcyPUXxW7dpGdhrxYf2dGq0lUbdqhTQOOd15GrASHFN+BPFcYM
rfLWBYvj0db8Y9LsmPDR70AXS8RUqpQY4e5P1+Ma2kAqubgfQAVZcW3FcZu/AS8JuFIyJ/aSsJAz
s8fzPVgI8/0p3JLDdhzwg/Z8/DNQSD6tnItBiNpadztwiqpGimwXvfTpC8fPIuYjZwb9nQ4ETD0C
CgQrw24dXSlgr56AZrel9f+bc14qGZfIcIn/8Ehog7qShAtiriLFl2q15DG4qDf/vw9+1BKBP0X+
6ObT0boOA6WE8wdRwPz6SZD4qhmOSf6TKiNOj5CsTDQzcAlCi4aexVmeodTrI5I0PdrkrSpVur0e
gfOJegmOOFwBnK9hIhuaeuKRHbYZ/7r1YLonh9QpiqqleZIZfMJBkgkzmxDg3E5JTFN6TRalwqY6
MjUd+hpg+n1lwJWrnN6S+LZ2skUoDWx7LDm8zvXzaRC9p5gGism4S/6RvEXj5Rxdfe73brC0j6YI
PR0Q+mTG8RJxPQqkKOwLCkJb0mHnzGsVlvgTqoZvDNyVUaZeFzAvb5J+UmuqQiecZNiyX/ksZ9hx
Xav0iYiHF+1XG8wUSVmhyMTBZenwnZxwQ98QM1A1PL3rJm3N6Op5hePsLj1DhzHFTbdTIuGdNhpI
3vXUAmMf83kAA5URcZHm8IR/OBLBgLeqvyz65YGKfwZ4r6WVtAcHUAKJKiSdwKVXLGI63rwetgu0
4IUm97z5qQtBf0lMEnDAY0GBKZPjtjUjnzW0+qi2TPGmbr8uNt6xaENWMQiCsUqm+ZI3R/WwNqSW
XywGIzToz2Ph4K3tFaFab1Mrg5tN1vl6Dhp7sHc1yph0eEmwDUI5sxk6RgYMCbE91oID1Wmrf2pY
PGs2/7Fd6erwESPB8JaBA2PsBBCqzdriMUn5Arsa2yZnvoJWZe1aCJgBYiCTHIQcKNlkHB5TyPGP
32FG0NLP7J0sVsG/788H4D2xqOnhN7VCwPJJK19Oap6OHmeQJl2Z5FANqYf54kEL1KHc1Nro23cp
OaKPVMoMgtthMBRNFBOa8K+uJMwmy9KyUnejORSlp6kIq0BIhye3u3ltNmZ1EwHxmRc/qPEPH0+w
6kJHbmxNor2GbKoVXvxY3dpjOorteTalbffpI/0g0IudvHFbGF7b1z1E62EOmm1vich8w7wb8E1r
nRjJR4+HNEKqxr5n32A/WlJifDpwbZzibCPfKUvrjQ3HAmaREdrUtgyl3g2mHmH65tGZkyDHRNkC
N1XNB2t9o/fL/WrIuFUC1wc1Y0ZFpXGI0IOUSwv55xhJVA91u7zOoVX2Ni5pQqPktVq71k1AD908
X4yxmy27ncBszu73/6dJSLbBFh7J76zXO3x069ZOm0fDg+iMwSHdCIdW4AyNmAo7Olf3Cb/qVb0V
m00ADA7YOF2J95wcNrU60BO6PW9QToJPZdXPAXLZGZ/aBXuorVDvlypmiyzDi9jFdsu17+GgG22V
8nGvGXI+rQX4NRCQPl4YaoVBBjy3mQzuqOb6QbMcbkMlswOhz+D6hK4IrfjVksJ9yiSVhLZu1H6y
ItRbVGzVYWvY2sFB8drZQL3J+uynjnex+Ynew9Gx8U6eQZzCm7uuYtAhE79pkqQK4ufP6+mpIdJR
OjUUZsN3CktDQkmqNjWmBqlhulzC/8cU+8/3L6h1ejAt/Z6kZi2WPZCHno4zko/YHscifAqpiHwT
bScJMXX/MoX/bKSFhQwsksx8lKcI+7R0sBO9pCFbHMHqR16lpQXhTzBvNsZrx6qrYKw1lnRHeL+w
hCse72mIw/BRzNZVWiG7F8jbwoMQi3PsH7mGVSJc8Ie0p0E9TFu4gy+mlNDUJfvi9+GNPKbLGdU+
3q3ZdmpnNiRUrrXqdNZ5alA3XP6ifVEtCqh6y9038brJ0hBws1iXiTVCaZ67rNe/MBMiF5MkOBgV
sgFoQD5Paqw1JNWPF/fsKjC1Zeg3zqc5FCNTAOwXl1Erxf7IsdRCOj6QOQpk5IJTYoLXkAuF8zum
LE2RGXHHSZfXIAi6J4OivFS1iu3YariVjny/ZPtDGOoXDJJs4zuQ51HU/H/JsWHA9QE1hoviKUUe
9Yk6TsRASoM+Az4nkSXyQZgin0aw0v3nrM3hKCduMxYjkrXgMqhOSf/WJIPk8/jpfF5sv7RfJzVa
jp2lemAb22/ws/B2b5ms5/j8TivImPYBkRWBjqPky+6imVEDMsidhvJ7JvSQi0zrg6h2eW6eqfqk
54S9MErUrAYLy3yQkYFszbZ/dx7MXxhxgmTfybKHslFpFVIkRq8RrRTgqM06wQop8glOjglQB+22
6ry0EzJV8MSYOfI6kRlTZzxzMo6x1CuJS9AG5gA4BZPFg5+6jhbBNfEX2XfHzcVAK4ECA6eWJ6qI
6T3KDUAgxxXJFF+lRDuzAGT+UWIFq1G7qjiUUxiMX3Tc499Ooxf/B8e8K0ocbh8UsXM0RHHYE3vS
h6XI2BvKkTzbrjHHJyin7thI1m3qylYNGL0YOQgCeuMdkli3M7izF6njSon/IgTSRK3jlDjrH+Ul
TK+mTXljYxXBFwyYdd6epx0SH+NezE5umo+UpW3uK7MpmvblCuCRRiDNF1beARI4i6bvPk0uX1pV
nDIy9yTWJw9IKO2xa5g1z2J818k+qIoAXyhQ5i1Tq/kmeb7PtklWKzohHZfGqi50cXbVY6ykXJk5
Hu3VAXAjGbIGT4SZdFTFP31NzsXNGK0XWUBJrahsXYqp4cZo+LJmB6g9/IfBBUeArrRm3hy0V1bi
eApuos8TRq9rrPhGzQjWEuB+GHEybMSg5ABPGqfDlFnRCPdn5q2Oytpz8eZvVU8qG8oN+ts/2UeZ
RQskH6IEft//MZMBw0slUsOnxy+6fJdc7vNGJzDKoGGRu2XUkZ2cgJrPncvE0yAiV4xZc5uUSVTo
xPRbNzhPqfg29Jf10VyJRFt7Yywhuo9e0BmTWPsFm0piCfWG3Z2OJQYlc1nqIHPfeiPnW5dsLcEI
x48qp5H6wVSTTTpdjavYGmHW9i8bM76rblEe0IDbnIZu0/NILu6f2VEGzTMgXXA6COplS3DabpL4
ZwUbPVhykvLAVieVlFhZUcrYr99E54UMk8ScdrchHsKGD1knM/yfVQAqLSFHhM4YCWCWN4zfSO1M
bl7tZke67P3Mqatttl8AmjMFMHmhSofyRZeNnJpBevXRoh0YkwFhzk8J0Btc6KepfVKJb2PA7yeM
YrqZ96PaW2pBkmTcShCJyg0bGexCVxygjRi0IEJGxsjzNJvphbJSSQBciXM3vubpaftZXvDOcqGR
aimQLzlX+nFMmhX4QGz19pS5RuMpCVhF2ASp2qlAWv1QIybjeMaPlJSgBr+a2FAFEB5oQFEkY1Ir
FpUM8ToRVvjf5V8YZQt8mmEZK2i082ryTfM7Sz1L9sFSTvQ+OicG85bBPA55WKMG3Zc1qyOj0t+5
60heI8y15exFw8JNv+2e+Isibj6vT6NKgI3vjU7MYpp8M2bGlHgPKqPVvA+fDuuvfdVsdqVWqO2/
DyzjyutkRnY5dofR/HhI/w7A1ar6c+SOZFAOxZg8iwsbBZSnJLOk4P4AL7IkKqQdmF6AhSlN3Uem
ZB1NkpufcEPygcOPwTDA62Yi4m/Jv8tuOg3+QJZ+vAexluCS+9lgiVMVZU8WLUZ3Lq841jU8A2jx
4doazK5kMQhCPdcDSmLivQgXrWfuuQKWGLzZsPPT68ESyBvSw6AIkWQ4+AK5Vlq/Mrgk188iNchY
niu7YhgEmPqc3HJhlz+XfcdPwcX6HubD2YVTLYDGg4aRMYtwiEBGnfp26utXPz0a0Le08C9m2Aiz
T0wnF1bXOPMRI15XxJb1DDYOa87wkt/oGb7FpGikK6PERfsrDf6TFsiK0E+10kVYG3eDgYVGc3KY
PtP65+RaE3B2eDvEEjZLbcMUSqfg1sBKwCD/YlGBc42hahBw+4xyadWxNYSiHuleQEefg1R9D+oY
KsKvgDnNb7JF0k97Xt8XdS1rFvJ/cYUa/xSpfkjWgPL0f1MgUO7x3idwkJ8PGthuaa+jsAglVRNH
seXJaC8Lh0La4vtVtpo2cH9Jq8kHW0WmGHDHaVrsrAmucAdqKnYc2n95AIvPdfEphOnCgCX4WTWp
P4jRXTrstchviEvzRdthcAvoZH0+gpyCsUT/Ya04OsgiuCEjSXtDkTZ1e3kdHOTXT5DK4rf6dZ9N
/9beSAvR2arxe+dkYtzzy34pNw8aGgzhIIXOVsBxoV9cGk8j04AuZcXa9KoArG5miEG0ct0trAFf
5HfseiINtOY+yRg7Iby59t/HypV8J/O3Rcy5hWNFOFOJRZE4cJg8WvoLn7xdnZhGrSshNtDDDUag
lP/T/4EQGUQuUdPGTtzuBfwnBCzJi+sGuw7Q1ZHkBuPzgz16sYeAiCUsm/xGogjp+VhMYgPNdXCK
Ohupx9HQ07elpnUcdMJuuRNuY/t8dmtIbSsz5WSMsGkYYhE0+nfuvNKDOsyjpLg8wnZHTY51qg1f
FXs97P9EAREd+5IG799kK9cgm+WzaOZ6DrJljsvjXxidkWcLm518HZfuQCr/rAvnNQJN6KdDVMkN
Kb/ZFcE4gAVWK2rDbTDiXvFzSrc9LKHyXCG6lc+IyZ6xG0a5YrRImcW9hsjNVs4XrWf/UK4nLxKL
BkSmbewG0rnRJ9XBWPBCfnKraHBUK2ce2vajpoXxrKRA5JrXyaZu/Kdw/HuClQAJ0s9iJ5V/C1Nu
i3tXi8Z1n6hMesX96/sotuEj+OceGjIXMsaiYdtdJYpmD3vAIJ2M8VC/16GmCsqSK5YUu5CshvPF
VYIYA3E6R/PBX/tKjqCGYft7OjcBKHXA6AJLjVAbFj1/h8e4hx6hN/gQG/LB15eVpbzU4KUBfxLo
YiW2dlzds0CLXPzcmPa2jGdv5D31mT3+vP2lddAlXhifdC+dfx/TG9n4vEwdVCiwJFrcq4cocdkD
OVFpgVx7QEwhHDkVHqStEuj5ZYjJESMH9iLk28nBT7xIiXIQCbFfPn+qWAcyWVOdlu2Nyf79Au0Z
b7ORinVugNtpMwFhHBPl4leNys42+B10TColYuI2FbVLkl2u7AvZcq9P74OsLJ417U5dFK+h9302
thUkisTeJBg5069Wlm3FrX0CoOSxoqrx23r7oe6uTPcgyaY/ZTkL0XWOBPVYj6LSV4FtBfM/1YOp
IkOXripwvTMvMIsBxK2WLCizIr9LOo9+O2yqjt9S/8PocbUVAEu3w2wJPAwhliMdOohaOXqqtzxk
shiSO2z60/9JrKc6u74t9ExFlSXDzOTNx5s1oM65soO7ZD2rZ6EFqwIZegqX4d6UxQk2up5KETtc
hmAY3JIXwBxwD2kAExzKY5ZBIgUECd84KJ95HyYC1Lgr4zgtFWH5d3G8Ap0WkZzNWg+gvehkHTE5
XwOCtYdrq4/6Y23zIcx09vtPgLWff1bdN6OhyZxMOGiU2JHeYMQzuB4nJgwWjad7+riF2vVXT3pB
1bHqt0T/xDY6QReToyAYWxstnFqkTEGL7n2D+J0QEJ6T+L3JGBYRzexPDJX32RNn5xUerGZK8R2f
ig7/8AuQePIm1hi/E8wjjHq/eZnS4ombMIr5hkTU03HZfRtZjXYjWI9efWMtFmtwDWaZ5yEbHNSw
h2EkhKCq91P/Jrh+apxnKsBI7ACem5wvAVH1spK1zy7qVmMb55FaeaHZCqVJR8LHDrGIoRNHtXc+
rJOq9rP1X7W7/1MGjL7wDE3K/OrubENR0bPxK7y4VPnWKctHVfNEKLY1kDZA338LLkhhSDGbkDHA
kEraAgYmQ3cjN2mGVdK/JuzVUc0mifGp2Cb6tfO3nYmyd2JuccKYD7+A7rWutyNSjaa8N3I+CVJ+
93UQGfUs1fY4aNGiNFFSwVDxV9BMJWUBJjBsbYSZ/CRykLZVoS88StI30WWsiRRgzkpczIDbh6gh
AisRugaRxB+ojOn3QQxOPV103fEhgQgf9FyKwTp3YZ8vUqOxtJitscHN/azen/ISoBLMAi4CxfFF
91iQHepfOWj11wzdp8nZCel8CLwkj+dKDXO1F/I2lLC6/8BOt+Fdi2Yb7Ny1a7g3UvbQSyDGN/ge
7bYiTkSbAVrsZGZOME9dfYUeQQrCeeaAGF7ObkSvG/j2AhpCnAjRzZk9LRSe0P7XVshpyidbBX79
gc88ra/7TJrCraf3w2vR6dSJkFhkQYgn5Pkncxhs3jD55U4AjL7DPpA0A2+NKKmdsilkrrY1WSz4
Urz82adv7khVLK8QJxY9RL+oalOerAr6fgaPyfbkxkd0sPSA/D628CrXOX21R06yYRNECjBwwGol
ENL6J9phQAnu2GqFeIekxoBUY/Qco73vrdpYZoFvwpWlWKJtc7VvY7QSvHVmmcSGq6Y7L0KW78M6
/xKvYEjhjXi2RJ9N0ufxO3YIAKG+y1lwTRL144fSoB5Yaidy2dNRY2B3ZFzAd63kyQeTh8Kck2Ra
o39VB2al0mo02jz8INk1MIDKqUQzfvDkG6/wT3FgTy+keuLlPxcrGCODifrUQsN0lTGyG56iOEvM
inzvznFNRzn2h6OeMmhvjHjbefDQC3UzUzohNZSFa5+aMcH4g+b0MfPNK45Ff1r0J+MFXmCDxhEK
1b+FMijhUe4/ieagEyzKi3BLbyygg7SdnxIc0LQeGTcOSz06509HYAuo9+MDmpjxwMAKfkz8pIn9
U+hskU9vKZbeRkw39K22VyrJn4oZTmJaIxU0/eJpiC45QAtn8FToVXAEzcqRE6hUOC5fMuW2W+kl
n9DH2a1hQIIuonhWBlWM79vQ4lbPg6TMHyx7xkVYWTDgA3J6kjOhu19/e64KPHlG+28szefeNl0N
+Z355wVEdKNdHXnF+A0aqvtKD3jEn1hYyZZDuMaWVVX8vKFkBi+63oFmRBDqY6OKSAvBn3QBgJSs
KIWR9Ugwmdg+XQmRbpleChwPDZwGnv72dUptTTllufbBFiRMTFgS033DQZO1M1X/ZQpY6MhfMnFl
MK7REUnJPJgP0Np5dU6F8atBehBROIvvQicEKg6/1M9lD5nsL0cjxBD/FLNxDGEcIzI5OOq2GyWJ
sRBo2Cd7PO71s+IRN/Ou/0jjwUwJQOt4C8NwfUYNyN8In60IsC/q2IZdFIcP8poL4qThZoXhXwXx
Z8HdFocHPsk6t7CiCIXUjbp03HKL6bsoivHR3t1iWlo5VdR5F+dY4S4P/nC9roONOsg3ZhXhxywx
Fx9rUIbIKZF9ndJls7B7Jx6YYF2ju/TxvRgIvmGLRqNLumUilpJW9fhppenQyR78RYfgie/bhZGl
GIbiVkD8DQ5eHzVZbpZhrkb9ToZr1sdPi6RFL0IsUD1nlXWWf6gddFak7/ID2b0DbwVM5WLDSn0K
2BOoEnkIBo+RqByXhZo6TdJu8ZMaJVRtg8d/s2f4SYDocEX5E1e2ctRw7TES13XGDEFMXOExaqpk
b4gNE/ohFuFzxUiUn/8EaGYA6stch/zIOOZFGjqtRJMJQQfooQ5+mnmIWPehBkpSYkHelNimXrn0
+la9GuZ+7gIk/E6qK0bCjYG07OWx5QWkMlYLSaZ7YDBVcQeDNLFWH1ZUG4f09WXs2gNRtTE4ugAd
cqGljVv4hpuwG8R5yAT6J3CItVuuDa6cF3SmIwZiOsuuYH157zsZO/Io7TIn2Om5iBmUU06ehaQ0
1e9KJLMVZ64eAYqmnYPpnzKWZNxl5tVyRdQLobSmk8qjYvQxhck54oclcFwmi3+9Aa2yFDD3LvJS
rFAct8uBUYsGWl4KsYeaZYemfdk7B/brAqpf8KiZbTW3IZCHpi58YkIcfCLrap+e/9yWABR91gjq
MsrpOHzPYzQW/fwZDqb24CFAUQWBthbx7C976z2XLbPTNDY9qxrIWIcpvzaE9ul8bSjMfSJ38czf
p/wEA+h/uDkiCZGpr5/gnKnUuys9UupiR1vhfwkzPRG/QFO+/3MqDIvKbq3FxEhKyhZidr9eK3Ry
rabbQgSBzFLX7MQkLc5/s2ovW/xO3J6W0cNjATuI2Y6HW7nDZQcw4T4ZE2rIAzlgfIqI8qfiVkVl
7BJ/YB2q04jra9iA6Kxe9BdwU8xNBm/aL0jIKSlzIh1skscJ8Do8BVsweDBqbJwYD1Jkv37b0IbS
RDMtPkV7WnHeK0b/0e6ABY6hen1SWrGtMZIez/hitwHkjzGsube0FQH+KLojXAl5wcn7f05dNYy4
itzM+SL9qA2wdJpH8EzV2vm4QJS/Xo1GpJkjBOXM3N/kQ0meBQVCqc1xILUUS+ZHxDLz7Ka2fQqj
pNSQUN1jLFp6wek4OMOY+qNFFGo5ZoAK5JbKmyizpiMRbLOXN99OnVAysOu/WUKiFAaJjvwvcIrm
uvx6YBjM6VHKI6RUN+CCAew4gtU/t3rYXCywubirOm9tyIQgKsB2wk2Fsx1Cid/YxpPuC/qnoyIc
CCqm9fok1WUqSavkFeQ/RU6zagGJesHAco6b9dOpjvnaHG8JdoLkPJqiDyx8ts/Uyx55A5G2WzkJ
C+NBaUHz04NEmSJ2pxEFHiPZF0udyV1lDXypQaQ/1m2won9QgXcGwYgx92cFSP6FR8851RdBDvGq
wE6U1FXTZHlbWpjhk2huAx+tbCloAP1/UVpJq74Z+H/8EKi5H2scD6qWOx77IkVYCkV7QCONlQMz
JYKr16i8VSoIbgqUK3KvOOEIXRGuFWb4YVQ6Rnropl9zJlSOcT1frGMalHQ1bs4bDVIS428E+71L
uYo5F/sAeX/KyGVToojy8DKXthZ3iHgXV6yniKf3SucDi5o6Qqe4R+XM/Ol/5sZ3ZCyhIoq+vC28
LD/EGUFC4tHf9AfjFXlFs04K1/tPO/xWdyM6o+W/ItScYcKjhVNoyd9SzV9sNEhNmdnQ/FP3jtT4
MdOphQJ3LWrUMFiisCHXn97boTOelm+hC5WZJ4RD40Vr1afQg+XcI/pqO/eqmQPtckjrTRKo351/
vQDCAuWbOATap5f9yHKnXBx9OISJqEvMR1PGfFvhLO0P2KMZz2M4tk5cr95uDJq6U0xF0pmJXTZZ
PlqRzYKpQcic//eq+6VJNzIVwfLzpTd3+Ce6e6WQmKV8T04Xs0njcbixDQlOWNujtXNzjOI0/qAb
4v+GC0OFtHl8UQ3OLwLvtW2ZN5xWjXOoOn+R3m15t5MxUMrfXEJvv2XklSSugKHEHNgBygjPc7Zm
makxOO2GKOAWxpgK8IXj0FeCYwc3j1DKeCuESNZgptI5nY999tlRz4poKN0oNw4Jt4AfSaWoRRhd
nTVRVNPRwntviUwOKr1sbjohlEF/w2Dz7DFPOGSX0CRHxchcEd22upPm9EjXoLHdPQEHwVtPIzr9
q6flzbZ4zvelMbeOKgUnsH73ZPwE9RY50QF0myd4BiGhy6agYXB4TCxDVfiMZcpFHVaK8T7bap6C
wZwN7ljjNapezcszhATKfdisimh/ymez5KNK2jKbfz6uOSiUkD6rTdKh3tXdNCAoTaL+VFdt4TX9
hs7lJ2shLbpbJkdSQTRjJapTYpdgH8qAl+l3YTcz8X+fPEjOKSFQeOi7iSSz+EsN8fLEEKMEAVYX
NEe+YgFgoRPVYt7OOHl8p31Y5yCo0f+bDpg9iHv1BK9RH3C1m4wlOIHMJe3BVfa0mf//RYBXEQ2Z
9xuUSk6flCTgO8liBknBn1vEnWxI32B1IFBrXKtGdIGszXcTMyzz0ZhI+yBsq9q/o8jt69OmRWke
kSc9xj1yD7lBiSvefBrk5B4pbWzda4K8dkqboXPnOKZzi5vHjnYBVddfQEQPeH3F4JF+DVxT/0/k
cD0+KxaCTPPLi8B9JUsHfkYlhZ6nK2t69EIlXhUhIYPqNRyDoKwI8njwpccJc4nwx7RAwsXfFnr5
kSYFk+7gi6Ht4U7tn63tvXb5sil9L+GZV/3uqMbH7F/cUxh6CiU+/G335wG96cd0HvSU8+YeG4od
tsz5yu1+2iKP5B2v/6swvJWhbNKZYFAVVgLmE2laUgFaEnhT41k3w1GewaFFz3v72m5sL8DlPxBV
XC8oKMhZsyxhdD4w7QCaFwruImAUKLyqbRLhHoAmKso05ca7JMrxeV3yrdkzlYOpkzoy2eFDav/6
I8lJFLOMmJ20toqwS6ScdukcX9IqT6DIpA6xRz+oMs52KJsR/cKZCgD+qB3uY/zyZg40z4XyRQq/
cq2LygR5DdOmVZa2XX4Llcld1OSS7Wig2hbnKB7R+O1C/a59OtWmaJiK0gJJN4dCpfOkBEYu6maw
qkA+dmko+zLqfKPYR7yO7BtrRhavDCmMQSvQYIlp6LZ9PPlIw1UKTGIENC9tuWOoFJE2cylPpsS2
vBBUZzIrBd4cSMLCPuz7H0O92bTSPn4tRDjPWqVHirxyXh9wT8XiS4tvTUFnjTHNx05FkE9Ru43Z
Gl7x+pCEOFF3/VUNCNJZdpE2a1GcQcZYcg5tAiI8ZTR2L2efrvy7BpBUCREXdz5Tn6rxCXwD0WAZ
MvECNkcU5PJwKlPtndHnQepsTXp6dD/BJJQFORmXdWQL+bCbqs0tCHAY8jIZhpOfLvrcYb+yH6OK
Wwoo/oXJnuA4dWVKn1XoF4AyPURv45o1swUoEeXG4t3FBwxiGHL9kF+30BPJzpfJ7ripLmamnqfb
zR1AeAP1mPyqQHsTCd7TpGK2KwKU27cP/96CvQ3hLeKLYT+n/15Y5Hzg3bsyC4ZSLfvUn2xw5Kh+
4DpFvdOcN0C5aYHiivVkcHyhmj5wRgmVnqyEBC7oUtfK/oPrhnW2rJT9oJ0SBCQRSib5ex3e+3iJ
lmDdnRkDbxbwmuUSHlfkjFPi3CMUpUy/aHvYpVGEIzfz4fBPDo5STtPlenvBekkKgv20gIQ+NZNc
4uLGmLFXlk9AYB2BYNJOoRtklNtPLZx9e/kqUkboET8wgxlkLOtvB4i4Dt+/xegzCjpUgI441VdE
tp8kKD1jscw69t7X4QjuqsZxvx0B/l2d2XTxbPh1tzYz0YsbSNoRZFWS+05dRnpoDkdLqDupDUtb
gf4YhkHkgoGfH/Z1mFweUKD7dLUS73T5wlA2kZv1W5himz4WFvnbgDcGZJJk0NI3OxPzlZFA6lZN
AP5VLv1EsZKgJ02vvbu1pZmdgduMWikhBl/9DamzEjW3b8oilHG/DjbMJhQAlc6ouyiQ08rHCYdg
2GCcGDfoEehrlYjqL1E8md4R8Ulht+lR8iQqgJkkERIXVFtd3JA9L4PLL7XMvDuLIe47UtB6nvye
yeFx3IVKIp3pfdGuzKDft4qltpCf8Ihft3sVgiO/N53Op1rbxWdyfC5jsu10O2ch1UvPDKbKubvS
K8HErqE+EWtqG20gS6dsJjforGUxKEvBl1QPTdtEeAVmlXjBNEzt8daiQRP8XVO+vtW8mHhRbeRZ
mq51BvJsimBHk/mhpRn82P399b/yJqpXrR4vxT4956zHhmOfnaS0PHn+oZPWzfIYkCoDZ0iQ3IHt
nqpvFN3lY1QE1tp4Wqd6Y5trNC91IVBptrGHaBk/oB62j9YV9mf6d3jyAMqJgUIBOE2OzSkfnYnD
RUzlrcyEqTG3jllqeiQk45aRygVuUiDxOJmLWEbi5AR+txSuO23q1pGloxhKehxMun3z/ccckBKv
or0in9thATp+si9OgyEkjz7zAAzxlDBcS2no4WARkQ1GiXv26HkmuCdpMwiEHqTdVE1/tTVmDC6s
aT9Y2BB8g3feY8DRiLWkUQdfm13N7lHRwiv+zP6zpGqw7JDwv849SV3bKR7KhfMAvzI5eaWeW5Po
dzUiB+gAyMMBAm1tX31sjLMn06w3Ib0yNXF6MfF+3l29wl0QYjzqojwVvZN6ieiIml+LYloV6QCg
YFxQQzqvPJH2ap0JGfg1mvhoW0uTplCshYID0/S6bfLkeU/or5ivqd+cjfsdZClSixxOEIyUfule
rbth5/w/1EeVuU7lH8W2bNnNycrdXryEs4tsnIIlRhk+E78pCPfWNVGySsi7xNHbylRoRMRlFmr4
qHBN/63GrRRlC9InbbC4g3BC3CgqcrEoN0y4f/IwjIsaY5PWzRb156/0f75HNOgw+uYeGVnO94Or
NOgvRLnejXdDQTnNRylqL67w+p1lVNkTKypBet7payPv+9YiI0I8/DMVrMy1bTbr3jOBB09AqA0n
fxjRuNO7liX8slqos1IID11A1OyQzVD/Py9cg6Kvk2tsAEK+4AATA+kAJG16U2Q21VsKhU0tV+gs
pJD/ly9PsVjkWeHx2v5Kz5nSLR71P+E1KRolze9vl8fpCoHGckk8s+jdzY+j15aW65wtqSG1wVm+
lgOMQ9rLSwQpZoLnKhttzf7QNaVgZAIlf6GwNInr4mUx6+6QIDcb+o/2UFa2/NpcuzEeE2FhZcKN
J2BbYUoiGclVa2IIBQaT67OpElR7rfhGFHsqSBp8W2BBtIngE77ZJUB0M439XyAk3bGEJ4uoGdE4
UnjlORHI7OqXZNligW31YA67LW1RHuv1cEUvJNeOYrB0QXrd+BcdkfSeB9o+kj+Yr30XNAB8+24j
XcPBKxi8QWdNu+hsvY/uOTag9x0f1jl4kZtyjTWcR2Ma7XYv6eTtVqBbpIqopuLr0E77l6uYM0NR
NdVXU4ggjQKs42YIL9JPX7mj12bWVLU1WgWquKl+1NZkMJUmxdQ5yidXs94DIaFsBwbKPR63JN/Q
EbX4bPQQ39bBnZUTyr0uxlLT3+2BQy3qeSgHTJ275azqmpidu/EHx8qTSklYTYvpjptO2LDppg5j
NCk9Ty7Pr6Yd66t/3Njk52L+o29AKGZUcStwa22JlUbFp3rTvzbofFxCbbao8c4EBseF7ZFBV/GH
w37EvxlQUQXtdEZ/9czX4FKehRD2FTSiYq5jGLH3NdjtnVMhuzLyLevXyWBTGilhi+7WNLlBLFXq
8+nY05D2i6sSz0ZCeJKccSgIcB01J5qGnkKLPKXiOrSZwc8el04xWW154ogGd4tF8qzNScN8Wo1L
w0aYIWwIuYdFz3hdQKppzyYnuOR9NVQ5VVw8iVRDi80Vu09jVUV8H/wgqfzqnnfz3CPK/CCY3LLi
oF71BIKM8ZK61tycaiY/uf11UG1rrAkbPY1wm1TP2DJ8Orgi+Yrej6xeFQfzjHq/SHaITJLsnKR5
0OK6oXVkxQzcZ9nBhleS7XEANJx4Payo2d6jG0WF1NroJKcP2NXma2GfbpDjtuMpEDgzJ4X4jJM0
WHCUWNSfxLyp70AXb69MF3s8jjgwtBQvRodCBXaOj72NFtCDBdjFyuhcNX1fj8hUl23pdFnOgNf/
YN6n5Ap9ji4C+xcEUmGYRw+AxHTQPL9teK4+yPK+lSMhkLVmxr3VabMpveQzXjDdFetNlO8iPWj/
g2TidmG7ezqdYwskjgqNUbyPmT8YlGRK/pmDfaYX0w1U/V+D4O47kZUBZB95PLuVpUxzq/HEwZX8
U5FkhRt7a55Z7LUbzxTg5bJmFhHShTR5Wfzl/s8L9MrvXquDi2DmW7fWxH+qL3u3L655fGzr90TL
yl+7vi99Lz3efQyXqVpKwiHzKweuBSn06NqfpGdle5RN+K/YJ74lUk5yufyyO+uw9EyLqWgJGx0T
GoGNdyLZBXzeaoAA8+tSIoe1o9S6CZQHcfwrem3S56q7lqXERWNcZn7vpomfW8AOfdTmdd+7cpW4
MbHCDFtGkBjLiUJpdZWnsfQrtXvBhqmr4sMiZBTshrSW5dldHNjTbOiFfzDiDqaGenu7VmstGsEr
c1NR6Um6KbGRnF3TQp8zcQioizDEjVf2ZsPedmIYzj5uavYuiADDMvXqBO0JB/K/e+e5ZJw4CX3u
Fyd9UTTkAIrHsAOibRc0wbmbTP5z0Cw9B3gX+E44gvWtZBdnKy2C9LgI5SfjD+B4HZnbPfovoxdP
IZqCWQB3fHdmQw2TMQvfGMkedg3t+K/JGayCcxWclhU0j2kSWKHHcS6ptMq7lrOpH9hK++ZQGcFl
8ZhcCWgcbvwM8MQA4Tlg+fjvCPFic7AdGDpxkk4EWzjYxhOOqn3bdKkdTsIGNBW/XmGoGh+9ufC2
v9OqWlhUl+Fv52a1iOT7X7KYfRjTXF8Fq1r+rS4pxMR/1MisXbL3dFc/QAkauziJZ9W7lZmLjinO
G295EtvG5JVVJNlH9IyBMwWG5l28UhXSQwpmafgevgrwgJMDDPynrTJcF4G/RWAjl2usJJmSaA2I
bLsmNM7m0cvN4bIJue2bNksTAs5dhXfvWc0L/daNgo/1gkm4fU1lnmrdEJiCIQNFT4aUKfKshT35
N6g3hEEqqm/Fs3yEfCx+r0SWpS00EdfPmI+MXuyfiYEyPDMZ6Jvn7sgMCok2tm/O8ptD4DZ3POrb
y8GgSXYhJB+AEvo0N7B+aZ29xBejg0XQc/6uoZnBJA+iAea//bk9KFeQFq6ie9ugjc7p0KrZgvqc
0MC3543W9GLgnJu90/N3K9Ch+LYPbxJs9K59qi+giO2gQEjWLcsyJP0sF6TM0DxqqK0VuOsmTwGr
Jc3dgh/MwYyEU+XqMUHZjbPWMWaPBdoOorCDiKOKD6JVJgovslqT5V+ma9Ycm82wdwrhhkl2EKmk
RNaGWAQmH+4oSIDb8WtEwM8hwTN/YrpHV4HO72TSn8yBqAjAC1swaf2/wdIKdO4x+Awm8y4g53i8
SHp6Sl/bzeEoOVe7XqXpho+krjJ0ESxWBFqTCSjtmBdcqdrJMqNCiJyChnyWtYp7lFuxXSGIIKuk
On0wJxEDqj2KGpxUCAgFXFJVpTj34SZOOzPYOZRdxwtKTl+6XSmdAl/PzcptVFT9AM4pRZxWEYtD
Gnb9TBARuKRz+n2wWfO4k4vg2PLM2ft105/fNr6dw21yR5Po/7aTymHWJ7wpL8XSUgVXHZTEOUd3
zLOBwEXPiVIFTxPhN/qwbL11Mw/+V9jRP4Cx6Ca6KgVjDwo6z9YxSXkONei8ohKBNozZHxyosjjx
+MpHOMCcFaJ0EyXu5SEqYBJg6+SB8hYhcLCQjd2ap3ilzAU7J6dEN5o2XFumNLJHbAG5SPJ9qTgJ
fA/W4P1yK+FDTwOXwCnxSvfjs6OPljf3f7hI0OKyBqk6fpbGugyhdJWZIn0CAkgDo/JWnh4Avm3Y
cqx+rK6/50ybJK2OGck1qSQ+Hvl7CzPlvDXewrCHCo1xwB2250y5SIHsS3ZWbndGhMXglzinZby7
BmUmeQ9vuRKob5injOvA6vuDXm99QpOugPUV/w76nXrBA5/TiIthfaWUdBF0PzwdEVcr1pl8jpeP
d/tASLov3EssU7wqHF5WWDWoBxYeL7SSlYFm6iMy6zCFBZiSNi83abG7ktfTfca/cxKIz3A1+tPA
DRNH7nd9qV4/gF32mHMbTM3OCjQC63ZJ1qhH9CyYNPYcOPB99qaI6nnlKZmT5rTkXd962cc5JOUc
ij0pVVZXEwo7gOBwIF7i7CoEOt7vvUyHuE8S6yJ8P94KZdSS5Yw3XYPoGXdT6UBVA5dnxx32MCJq
q9tLnRR2WGVdfNakjIPnR9LT6fZ/Af4JFdoRC5iLgBMC/XyU4lFuJ20nvQb0HiN0eEkchqVlKV8x
T/bLYvhR7Jfx1gbwZF5NYmbvMJ8YmGc+5+lo8HZ9dL6K+8FPCTOHdyv3TMfNE0+6j2xnZMFaqWQk
9PextUkYfFpXsAyQLkfJzzDLULJveTAgLBaNceflAUzcTwAD2bfY5HbKTGnLk/11yvwnzC1EbScY
+OSHZn3HJuSa73g9Rkh/noZqKQL0wdJ1H6fc/lQfBW4cOrdoKkPSGDfpsYM4PErydFnNn3vQpW9Q
U4h+D372z8tjcwQVCmgs5Uqf8qm/kh0TOkAcxb6lux3P6GBIR6GO3hsVqJ6tTOoGB1nWQ6RJhIbN
MHrvTsPt8DSFE1Qxi0/nyek39117yt1WqWyYpCT33KzrD5hPG2oH/Ry4zzU+hK7fB6QBcq5+T9lV
5PkuHmK68zIDy2b1N8GdFKRuqmnXgEkHceBBLWOLuBOCS7BK6iBB4F1pBb0UPsM57aI0HkqXL0F3
H9NwG5ErnAU44YfltJOVTrBYXD3W5nJLlo4mbGQdozL5jEx67HPYENzxNEwxSBt6g0ppUTgBdqpG
mu0LWubqPD9Gpw/x6eO+WKG8+0xbS22beeHUZjvUtz6nxSQkmkxcuATvh/fOofaE1TGN6CDkPtw+
aUQL0nvO868QbtEGGA0tcAwHtoyzxPDRj6jwCiN4vovIDuFlhjm3h7p1vmOXcQ0avXU1Ha8jqLlB
pIPOjmeOwUAeK0VuqvG7m5FSfw0xe92y1ATTZcztE+uUQ8B8n1n+E6aNaGeMEjJVRuSkqT8rhsT3
VKSrsrFo9G6nzxr9hVPgaPsdeudibdp1AyFcNBb84C/s/roOaLR1gVgVAyyy71IW2hDabn9Dp6LT
7Z9b3pBIUIhmAfOED9JzFY1gllM+IWCRbTJ3f0Y2scTFJYgqICfKmc6WNG9edxTuQGd88AR5Suib
Q3JUxLOvtyBY4T16cBKo87K7bfnaXuMZj6nbEFmn2MbDswMpmSzfDvQjGKAqEriJKHUjhWwnT7dj
604z9NGm9BndKgNr4O8z59EUOxvbQP9vQD6cwbdTcChxfnJlsp3YIUHTNOShT1LqKAMZSnMr0JOq
baTSY6OxnqSpO7hffzb+bbgAjJvt7vSFzJRAhx0Qvb00NC4isT0OgqauhUp/681/9YRLhnwyDCjL
8HTqHKGVfit8bNl5xintbsfhIXfMc5OFXcQSCygktH8QusRiBr+U/tgP9FevEhfvdW5hRSa1aTfv
JfzwdLz0wSSAFqd2CjjmafwYCaTt3olhvVrjt6SuPJeOHEEhVRhSDz2h5WiloclC7+waTbjbxjRZ
CEyGPf32uT6PNWy1YQdg+V4yio+ISZMGUTGTHezZ4Zb3Mmp+gh68bHNWA6LC+MyFGLLWRGvECF0d
vY3TutJJVUeNVR6KYaLoWU+tAvXD24COouatHcCORNNJg3YXZC7xdre5eo/6WgCWStyt7YeOy4Ml
SEhNqxi9YIrneciYbq3PQRnD47bTPFmLikUD9xpb6JYDW6eXaOYPtpQ15Bn8HmLTWLjiq36C8N7G
LUMg9AF9DiPUmDfC/vBe4QrJa11KK3ak2uXC0Pd1JPKq5seCC7hNIk/w+c2sY6cf1cUqJrgq9lWi
xztvxP09jfjjyHJU5u0JVhMpSOGIwa9TBNoy0MzVsN/ub1mII3k3lt3cjctVevyhsEr33tfUTlTn
uu5yN8gE0veHL7L3gwcxiHSzGNp+3Wl7ws47SN1srxDj6ZtoI9GBHDGRLhuO2m2FajFYxz+hCSlw
a4Qb0EoZ5sWseqlsxR9vUKVrWW2jQI6QWjGeHdU4DnKU+wqULZTIikEo0GIiigXMnoNzc715WbJv
0UyZ2aAxGPlrKGmvV6igN6ToZ072hRqrpCVnXb8dAIxFV7ym6qYZTQDHLUIX9L07k//2ir2mRgS/
EBJ/Ef/q0ThFp+EibWMsXpN5Q5wBqY64Dj1MS9ULvX1hQonkunpsh8GaxJD59C/Jo4fpsiW02z4z
3uD47Xw2BEgsPFU6TyWqieaemqlwPi6ID5QnE5DFbKkZF8oSk/Vs+72CEPhNUMJWMmKYa7Uloiun
W+ogoIA+K4WBj/maiAA5REcYQuuLsSBax8bjfEw+hS+mrLizBcMUwsIfuvTUu6ENWHpdf+lG79im
2tDf403bcp/v3XdmrE6ZUVqziUtbYWye/JSLWGmWio+XMGlNzFEYULoX014MTaNTSTk1joxtKNIn
zILxiahUEoRTe0+wpJ4L2DOzeWy9tYjluzPsx40rh3M37+cKRzyYh+ew6TxQDKEZJuNNO43E4ZPi
D3YX+tcN6pFm6QGYaAEbr9t8Yrh9gELd4DH3jlyrD276fyYrfNB6NjJq8hF6ONvThxaVmXoWsQ5i
2b+X8TZySMF687kVneq6ii2nm5SwFe1A4T9aFHQ4DYoJc3ttoHoFGEjFlwD9ai2ZVzc1wBP7SW7u
v33TU3Pd05UuI8+VJNPOQOnyD6JlxIIlJ1VYvb62mLkMCEGsJV4bwJDfx71XLjqtz3AmGajI1xNV
vwz4dHFD/6sOjhmiRFGuHpdl6hphw8R5Ry7DVqYCllIfK2ybGlLkqm/XSzC3l50UyHPBHFjI5+vV
KV3wWUljbM4llFrQ4ajE582nU4PuCtaNWQQCwqEbb3ORCVTWsAVMaFLUSMe9nOeBULTdwVWBNylq
LvPWwgIB7IkZ/gKjcuVXYFcIMQaIpcqMsWCyFE2c44krmZkJ/z1+FiAavMxPJm62edT5AQBwG5mg
+yyNVxE9xw2oq3BXJoJ1JVDf3g8lLr2UHun0NB27FQ3hmXls7htPHTKkhJf4ZkRqmCTqJE0bSS5T
JxJJTbh0PZ3LsE888OzLI3P+VXfeFpzsYmsf1RkIjFsDiGvSYlvDxbUQ78sCUag/5K1zBjAYPZqJ
plyVcJRY0TisEXq3b2wBaSa5zU9feMG4Qg/6WhyaFuP758xJYDxwniFRV6rf/0SrC8Vx+kuuXIEv
KOkQLfO8WhZ1z2Gdpe5GvvRxDCPMMLeYR563P14+SLm9AMtAUulQBkqi7dqA9yAlDYVoH2be2stu
b8jVCcpNJWlzDXQqopa8WX6Kry+6Cjs19v5WJY2AWQnbCsYOsdG9LBO5WtPwXzvRNbrQeOz391YA
VyofKHDf4zauccFFtsQz0EiPECeg0Gmt3ZesBRUdfNEvwKmufCSP1VMAq46XtZRfU8+sYmfQtwQb
7wCxIBLj6Oa4oyiufN9TvF0xcLowM/m8jCkdoVnMBt/D9dMtJiJhdWIt9ij9h5MjoZVaakPQrT1t
r0X1JqroctL5rj4wQAt8rfb9zKBZTqrj2TaUIIHqUZzIpjDOVvFfA+PM4S5YvmV260H9LwC3FmIF
5snx0GFBDcSfCTZcE0q9DRLHDQu0l/pJtDAx64aaWGOkHkHb4AEakN2fpRSFOMpULzFC4cA/u5g0
/yu34FbKGGs1QfcEdaIAY4O5CRNz6JjE549gzL63k6bu/laDtEcez8pgzYZqbhgG/TsYyuciPdmC
Y5GE06ZKhccHMFrEvJtVUfFsJ6A1OsWlCbqaUQsmdBuC+pxXCViblkIbVoXx3idsJ4+BOm+DXGPh
LC5CDiSWHfdfkswDAMP1iHl0i23Io4He6L4BEl7vJmq/K2Wzqf2I1ZLaytMVwEesZZuQFFCF3Ias
vVDjumt2qw4yrGOPOFlkucJHCfTp0ee1mFHv9BTzml7NS/iP0HPRQdyYpURTbyLLCGPqFQoFKrx3
/zB458gXKr7UG40GJMU6DjYIPj9p7nlX4aJeaXsS6WudWemomMs9WgJVAXsY5R2FBFi4+HtINYYP
rlh4B06TCms0KgShsANVATCzcdzH3cUcVSY+/1qQnKOMdFRylW+NmPP4OGaFCwVITAeere4zxR9i
Z64DrMydKH1HOo9FjWzednVG1htkz1hU+4UaN7tHS2+4STi4NPafiEd6h3CkeJ8ZkVqzhZEawj2q
YOfVr1OpNvkClKqDFPGKoSF5IP6ETqCIzS/zbPXwtkqw+hv1kmPz6mqQgZAfVxjESWRK2508YDnT
F0DEdauzjc62SkHmRMJfrc18CHn70JsqL0RbvU9u/AoFnogrc0TMK5TqIJgbcnaYT/bijfm9bZWe
Kef9hUR/eRFN/o+6Ssg0mZrSLkuvJsADP5bcWSx0bUy4vZL+2zOOjIEXPBIZ1CxB0MhUHs4Bm8U4
5jLO7VLEXPmY9u3cjfRecHZWp6x9vikAMyRdmbu21PEd7P4hBgFt0mE+41vr29ckhnWDtbVz8Tsw
55ej3S2m9QfC6Bw/zUroEHt6VehP6Uwyew58Jbh2GyhN0Pf6z1JQ1DviRkUptWAPLeInaBnT7elx
t5lANhmZ022gXOfy6cp8Nn5qxmFpnux9A5TMHX48ex3UVh9qiEUPDRrIOXTxTwpj1T9CBuZ+AFK7
KTDE2uWGmu/L00YcvY6hQR2uehd32HfVHc/TrewS85BCVU+fr8yU7KHyw4luke68ydV8peXkDexa
OA6CKOIbxsmbOTrX7iZ3xnGiNx/VfW4s7SW2YVYmqMjDMWftIMV8mjO2VShJrUwfYnrgccfIW1s6
gTDoaA56iwa9JiM1dLWDPZfmp7CsSvzOREFKZZOFCgvQsbO15gl/nnAKQxPqoh8vbB0GKSBBas0a
tm3DBtm6JIKTxAU0PF+FwXbRXpckxjdTg1uroI/SMdk2mtn+TQZzFfTiwlsoxSs54urw7vP1vvp4
2NJfMqkfmXpcflg/CvDfuPVpsW57Do+YEc6aZijYBYhYnM+EHZbnKnNFAz/kjdkRofKYLKgFMs5V
p16SJm2MHWIfBsN6BRvLSXMqcB/Hw/DoPFGZzhaxouHSC3LmPqoNdA+4v1DZec4xtjrk/HfFXKTm
0pEkL2oioL3LzTc0lOcbqiCemuYWYVEp85b2osNvxIP54ZbBaA+DSo83mrc77dfxxWsQz4sBcmFw
IQTCI8ep1bHUHfSNsyM5V2mYHpT7axbMs2sZf41SNb0qjl+UzDM4DUwPyKb/VOxsd/vTEHqrhC29
RdlvtOcATsfuf5etke8gH8KLs7rKRsIc6qqq+SykjIhyDVge7YBmE3IzUA25cRnnPdMKrvvII7+g
FbnPLEIZPhxwI2ZGWMXRtRqkXc2laFTbzGx4O+dsnrmCzc+G89HDxLh/FMzgMCbBoxbrO91FL1cH
SngeTJJwZjp2BXkT42DPlN5lSxO33bCHNoOnwGr3pA0Onm+DxH/P342VSaaUnNwmODJOJcD8U1mE
SBxizgRiP8Z8W2ZEsa27hE+Z8UtbBm9dZStwdl7luRpyqdnXUJBQKcATlnbEPWCdQrVLuRK/NAZ5
a+Q0rW5DHvnn4Uj5XwzjMsbE/b7tbu02BkIB/p1MqxDEr1/RPDG8RMJGf81VXklfoRsXv9ztK+RR
i5sF7Wy3bvhRZy7NGdJvA3ExoUzHJb8QHixyIQ/d9FJm/hPIPF/F9UEzKkJmcPAohB8osDmM8NDb
bYQk3cvIdQq6vPSMr0GiZnfbRZsogId4Yz1b/NjMQvUTCdd5DM5N252HMJuA0E4So4sT7Cr+btVK
bPywuPtdCBxNhGdP+yMiDf7NBUeh9PRzLOESQlhSTE0UC/x2MatUOJq/W6LWpEG3NIlNCBguM+aI
a4WPjJr1dPCSvySutBObuXB7FiQrVZVwz99IUMrBO+RveJ0gdFKXFT0jQYeg9nqptUKgIeddDJ+O
qOc2qQxL8osNxkOwmwmQBVA+xCFBEQ1iT1lTVjBe5T/ZogSdYcZPshBoIGh9DFj6TTQ+bZZ88LIK
k8RJ+9voGtRW8TNLxWKNzpEwIYxxofmbO+63pHxWIkwuK7S7RtrAr9WidTRaYOgd4XDCdsaDAq5m
C4I6nsU6XTcvC3/rQcwIZ51/z1PN+8xRmfAVsAg/tzh/Ci1lsJ+xBSgCA1As3n543E5EahpAvBV4
ny/B1BrJyxF74VCtCLPRZzm/zKM4XR5waX6Gwa1rp/yImO+962LisklYljhLWiIrzC5qd5no6wCo
QQe46w9KC0bnakO7PYaC90H/Dz55Nrv3/S6vExVZmC6wZUoGMA2UBAnJdCgqp1w3s0zvyAgeK2+I
se21UjzKIj5LrSTLHA5Qcl2Wp6DtN/fQuP8imqHuztG034V2EI5LA4gxBv7xeickQ89Gea4jFnYp
yLIqc6erJBl07wxDlxBNZwQhXi7gO6bLrjOWdYWmT90GD2EbY1vBTTWS42ARE2IMchoF836i0BnC
0FRqbcl27GCCJn88BHe+m3Ig7+yQ9/ym4wNQB60w0/B9H38hz2Z5OL3H5m6Ua2MgtC80ZSZUC3DH
mWl+yMarbNhAmT+OqkO5tTLqgt4uGCTmIO1h5x1wBQ87hP0U4S+d7kNWlPrMIFfiY5y+/+sYtAZW
UMBgZJEhfLXecT0VniGyc47ItI09HFA7bi8vRw9k6ASXpmeFnbpX+ZIkLAh7PbycOLDyeqF5/pbd
j5FcyLvc93kUj79sJVGdDXHCkdR5QnAgdsUxVYQUbhI3GtQls602E2doE5RJWsk/RZbFesTIb2dz
hLfhrh9WrvVmJip4eCwhS7n1Kv+tvs8w9XUUm5H8sUGsvkZ5mBrcxM1TnWlDTgcuOGnK6C4Bbje9
8S8Zln46f+fwmkPKFgS7uLymEHmCa1fONZldf9tIwO3gW0/vXze8PbOqzyiPNK35B9GhDwT64JcB
41mp4aeqDFFF/soSudIG/83WF9x0SDQ5a4vgu7/ml6qEHh0TL5Q0hrkrhbALlbU4ijYn+VoXO1VU
VIFe6X6ef8nOjigdlLeCy0keTA0CVYF5Dzx+V75ntqfezBIurYtyr7fAtcCozbdIsCsZcDg22xUy
o+nF2srXU3YOazrUmG/QK1inD1SeBdG8sDpiE978dHKrfZpsMI4qleN090/pweNFarWPShHPHNbi
K0KXt8Z27aB86o5x7/0f1eciqP3QlbhJVqTfEqBfarvxsx/4HHWyh4taTs/erRrfI1QUBrbfOToZ
v/T/LjImuEsKGuI0Ijg/F/YpzK6uO5rSQdzhHTs1epRfUtET1WzQ5ZAy94T/I5n0lp3gehPmNPVq
WVacUW07m5sBI5wPpKCirY2TkUgXoOtwNQNHX8NYZOtz7nwNtUUj0ejVcgummnklS36fG5/dVQd1
JiOtgQpBhqe0QMOd3/ZqnmcSo84EBWj5Qk1bP3yBnvCxzdSuJ4LqC0yvb2sM5oy0TvDWmhe+G/SR
EdYglV4Z+E6f6iklv4oRNYHM7qr2Sq9i9ZIr5E1XHXetb7jSs3vmJYbkrdPvZt2+1i0tJM7hy6EW
5nQzqre4aNF6czh+NCZAjKjKli1AjYQp1EIiAxG7YIRbvl7gtv0hsbF6jYBAh4yJe4jnvpFlNQMJ
lYpFsVIwCus3OhEmAyEn1blJncMy0cnlWroC88NlyX/LwucoyUblwtfkw0f1cfM1MbFOQTh3QFXL
2K2Emdc3YyGaUYPEAUO8vhYE1Rp1RPDb+OkDkN8NFIRLu4ZsHnmMw12PPfw3zal7yj+UkhxgnqFe
ZWMKb2mZV5DjD/qwuHa6kI6a6ap95NaeGM3gYiXUbgYNsmIISSlQn4IxXQgcTgdgv/KKg4QdODYN
KbYJoWmjAXY2BJ/2EE5r84HYoo4mbO9Dngoz9MaeoVwqyM8KRqvXnmlF+BwaY0HnpNVffXjoHA+7
PTBt2kGfUdL2wy8ifQf5UrhUK/FLDgzoDkEXu7JnhcvjSlzk1jPnQYD/MMthHBHslRSHm9DNzxLb
G13JGSrmXGWSdoYHgsoHEtaSYXTPQ4dXgbFvpnGw6oBCmJvUOQ9DVpyWopBy9/WJCHCZEf1LGlrK
dqlVowxMCJbOlH0UB7HEyT0KXhMJoIVqRsHprxXbUIKlm+ZlnpiLnq8PNjdC2+AhE/j87Fs/75we
sDKrhMBxlO+XvJ9vg8G2wCDpiSMr4tpBqWDq1pyugb5piYQnHuy+4CLNqQ5xSDS1ugAm6wvxhlL9
gUxe+Dis7gpzo/F/PKxtQ0oIWyP8mBO0lym6fdKlw6o2V7liL7rhBAIvpwJb/CsBy3XQg/eBMcPY
6qGlkw8wB6gwmGU/u/moIaGfZ9jeVosEJFM38kbFU6mueKxhujsM4tXE4bHsl7ElbutbBu+NBqAz
DngXyfeXdHnRfEBgymQaCv0o1OuMW22mvXMAlaXC0LQiY08os2f45xU2/jJDq2Wtw0vGddGNanj4
WfPUQQTv5Evh7m5hsrkBZSHJd8/r36TaSKczTR+tvlnXl14svjmiSIREMmD4ZfaZjfcs3CVM1L19
V6NLs4rXFNgntx1bXMa9mjZK0n7rgz+2U05IXxEudH/pXgmRlDSjn8aE+JE/vQKOBHtXVnYjBcGy
a/EyPtLx0Zu5eMTW1JNv3ZYyQJEvWICXX+geL9eQ7mFEe0Pll3iuoyLBw8UQ0h2xRDA2nTpo/UMw
wRuD0kGxtQa6MHGfQZXT7KKSCxm66hLbzLfIP05Tqr6CzwNv4KvT24M55xE5tQ6c8Q49leu37J4b
bOjExd4397u2utmHNrrJG3qYHv8VNrod+WyPvpIiI0uw7S5WmaPaSWjJr/q+RNJdoPtqTVIRjTMO
NJL9TYww+cYJ0mPS/lBozQ+qR161/i25IQz/0TGUlyj0n++vynEmjY4jaRdAMClQtK0/fHdgEn8q
E22kJeXCJ2f8zpwuuovwTfbIJl9gM33awxoSwPFDM97djAkIPZz0veLsPFE3CRO7ipeetk6jm87J
IOcCuCpnSRgIOAWtDHFU+Ymo8EpfKTdYN09Q5kOf5JJDygR5QTLoIaPB8oVfrYKiRiWRjrx/KaBE
PBPYAIDfkEq7jatR9umyEEIIak1FhU++et41i6U+fMRG4UDK1LJUyjj85KMlI/yErBM3Gwt9/DdT
+tzE41nqaMSHmDs6kjgzl4ty5/ckWXu5/d9xOOeTzUgkNFOJEZ1hfshvt/SzZg0jxJkzC8mnlpLT
2j+pfRqUZq1If9ciowCBuxOPf+/hi9guWi0YIue4u16cG27CBa5XO3GrK3g7A3Hyz0tR3hCpNAST
ec/2RKbZ3bbkBjMV8n6McST8QVurb71FZcI8U6JpjT6IFYMHVVAYjY0rtjKc9YW9Q5RFDs8Mvl/S
fMwhqDLqZT7gWTReMbwKBW/IpMnaATxescP3l/caDqhoLZEpfLDnqYTxLgSzXMKM/0jDZGTmgf0P
EqOKjIVsfq+9Jsr2Zqw49PHM9SDlK/pPLwp/uj1rcPEGGwTwz6Vp0qe0nJFbTemmw57KNo5+zbTs
OLS4hYoNvhe7F8wfApb9WnRbxrtwPXYt97avznJlXK1nynIs7nofAMnjfwWZdkBt4bMiAUXHkJTr
pAioj9y3iNdMZDZeZUmoVlN6ArK+fhgGwmtPV57zcrO63RgUa+DmqGN3OCxXhHQQa0dm5be+Mm8T
QNRCh2360pnprNWDyAgNEWBfXdf1LRnRK7m+3PkRZqhLUOIgykRPeEam33NB5BoeYtUmn2YoU7Z4
2I1gIxdAHoN6DnxpjkRjJ2co5JADvO9XzGr1okJncbDo31RUbaTV1GyBb3pU2/QjsBCXX7Eyxy91
oohcohdghFD4IMMFceXXZnKx4nVpbi/mfa3wMyUNA7WvU31haWwA/75c6/vc5gqAu6rN+ZMJPM/b
NUjXlIjsRMj+FLU4o9E97y+8VsWBLtmoMfRbVCD6Envjd+bJiPf8z8niRTqnYuBTC62ol2NwVr2x
L7N0HWrBW9dE+Py2sRIY16DCFJRwBrdieqXWY0atUCD1LB/nbAb/QdQKmNFsoOewPaRrupHD5B5f
43qNQgyorEk4jUDxVssZc2pganaIAqdRSnpBnbJmC2nE7EBoL71iBfGH5+xeCK2kz3c4glSUVRXV
eOWiU2p+ysZBvC8QQQwxhJTqd//HJ+RAwGOlJAVPx65pYq1Xod/+Mo4eYsB4lOrSncQMRsXGVoTT
rURCkfpF9GdUpamZ2dc91VhQ6bMdU61iUXyTpYFOIQs/Lh/2kIZHRfXd3feLVvnKBsQVWNYRYNmW
QpMyTV9uT4em7o1qQ/RrJW3wkYLN8ZQBMf0c2a1KaFitdPg+i7pF0R76181+WIf9BTDkMqP+hsaM
3bG+ZJ40fZ864fP5kGODLhG/t2kUw6VEW84/ZC75si21TYGjIkZUc9zj1GkEdBmrfEzmY/8NAjZd
fw9wPVfwhUUg6m6uW3BuZT2brdyeYfmdBfE5Vr+l5hTuWMt1Vy7g88em0DAQtANSO8x4un244oTV
VYO3Ul6SFaV6NEQ9J9D73T5q4oS3d0NdHK/k41Bb/oXZWE62+0tRd/DR0lUTEF70CrQwMZMeYakB
Nhf6VQ4f94gY/nY/APScW24s/ZIipRfiwTcn5+teBt2O5r2xgq1sJUzoD2sBBElfqOJ9ZHI5Mffx
pHsNz8c8+8m9ZOlMXTv+3ebBnh3zSOMXF+yOrT1AB+I5MfJVb9lvcLHuX6LNlLnjpDkkDZ6DPSAC
+2M3QzQQwJCio1cehXP9P2xe6frTdDXS5cSqz04hq7BnB6Fjkkrdbdp2QvV68582ZOQy8NZkvrWs
JQ406yyu4bo5Ras9lwrqy7bpv/BlpV4HIJZvvNbwt1miol57LV1tIQ3FTkYgdqVxO/lmAYcLF8ID
FKs9ZqdVKYXMSImnNKxu3IopbdUWW0UKDn3z4BGFtP9z7R8ze3SesxjkL3p84zXYtJbk3xtgZ2Qb
ioq1Pvq/2CR1GiNVZ9xuXAbwmDnHdvXt13F7YFUSVpa5JqVZcpM6RRihPaeG1UOgix5yhR4AVhms
BWWFhN2AggxSDGrLtc2GuOYPJv1NKsB5dXh2B0y6gm72nOCMh7awlraytAzIqzlOcL55KH+caFv6
QCf+GPmu0Jv/e5bBrcIV/QcfhRaqV4Dl44JDSf0AigqVRdO4zVpZg6KgrRhpgWVJOqTjLgZaHe4S
9OZSnMd+9bsY9AC0FUxIW20TpmAYOgiCLVKKQy5Ia5fsHeZaCqktOf5wHdAwG3bJ8Eu3wh+BPvVJ
rVfHLUiqxTSsm7aIoQ4jrEcBx87yM4tQh+LBmofXT+5lttAL0vWYwspxzSKpxs7PgzI6hiBaKNoE
FofICbeasCixrMLnQLurq8IdAifocLKc8UdmFaAArFiHIWDU6DNYvPCsiZOuhshaXFGnlHcGG7vJ
cBXCGTsYb8gimj4XFxhWoR6eIGXY8InkGZL0TYyc70QBMrQsccaBx9oTdUXp1mosxE3VzJLnuqf7
/YOLpiAWJaNU5v1Fd0PGshDrW7VcoO9kWWy5/c8Rcu8qP8U3Obwk9Zmn7VpfhArtYBcQbMqzd5yP
2lw9ZS+KVFXmlx+i8NFH/cqd5u89/9E6g+CYjQlGW2TQndpsxDvJ8k0GmY/C43JqX7yyhM/g84Xl
eJ8j5jbEQ1jLfOxArViRIZZ4Y+sGFLSwx5ufihDR6pGO9jwGl5Dbm/TsIG6WovbXLpn7N51rpvYL
DJsOsqtQxcYc5Y+UTyuV3hlfMHb1I06FrtaZ85T6zE9RkGNmvV94AjQmnCI25Vi6RVvajAjC/zo+
bU5Jw5K1RQBpQaLfcoTVVenQ3MJYrJg0UTLufkxooWnDWpDEEBY9wpxi4k4INB8nQbJLrwgRkJoQ
npbkFkbQEKMy9AD1RIuzyBpICVe3MpvpGwKIanbxaoQ7B2OnNZmSRSv1Z0FQOzGc4y7FkzuJzDV+
lYrXFwaCsZ1reGn+tJikrCiCzqkUBQkcNLguS1b3r7zKXqjUGxPtg1IqlmRwB1teUo/kGMvGTsDp
cb8zjLsIs44GYxZJdqqeuu7mesUzfBgG9x+ot6x9hIfxdEwZki8E0OcfO5Qp//lkq+M/eWFyN4Hh
2yV94i0Tx5YKqoNzhwhfe7DjwzvBrqRir+fDRiUTxK7vezlXg2NNhUJlWnU3JxFBpqxSihFH34dH
YuJJmLtnsobnC06xdBaPJrZ0V3hK24j45gamWJWNjiIz0z85Q2tK52E4ss7kqhU+lUXAYuK7vx0m
8exaxDVqHU9MkPbqjpyOAyaFz4x2dI1CoMphCUeWo9MtepEBHwSP605ao28bLVIKoYGKA0+dPg+x
W8lNua/wtkkEDcqXMantlGFfFINCfWjoxzcNM7LBLyUvpDMsy6ASHCOPxq+3bXaOyz5OvfrVImIx
79zASq4cQgGNPC6fRLFrSBfG/Blr/GCYONOh/UaxbaZuW0qHo0QBRNN8wQdOscD7DNXddoekCPrn
Gones0Cw+YaXS9L3oE6Ez9ruBN9K1jjBKMDgytaxwlV7GJdjZ3BS5B20aD4qTg6W3p9PAjXywyuE
CHhGbb0M/CRUdyOW/oqHrkZUTSLTWA9r/ghUf9UBc+umuzmT32+MxA/o6GZ5uPwEMn/4Ve6/n1Nm
uCWn2uuUGWpOTxlhljBLxLICass7OIgRqq7ljAwIXw1E7dcScEQA+zLoCgb7psrLoAnEXEchpAI/
akksBupflvbqLv9GRn7q9rM9AwU6UB7ZjMERTi+zEgqXtEllqGviO+rGsKEVtQ8WEdY/3ZOs0s4o
KtRcRDARy4pOSCTARnvJJ/+ZNrLsiWkyFuRdS9Cv4zPXyiHYt1utuUyP9C+av8YAJsnt5sZ522iM
1bLNklPGlNrjmIi1xpXPN0oIVHWXSlgLn/aeJh0kBBhjNJu4SyPN4OaUCZ8tTrmvjAbo+CNmlNWe
PcOg2mngMflpZT5Ofaujgr5JnkWKArN6y19ePtROnWnRK2n9NzsFXYAp3VbW83pPm0nEAGqEqq7X
jLxraLOcciFDiXKnxgXIWQh/TdWKOrpfEyUAoT1OwkfqiEleYv408+k6hJr1PlooMltJeUh1i6ro
HuNK4yoEO4lbcerKWNdlcsSefcTH3cjX/3i1WoZny0On03mGwkcyXf2j6L7WIneGQ6YQwvNcct17
meNWRZ/G9wFYeG0mmtABLjW9KrFQh4Ar37XAev2fiIrH0wKnZyakYCyuvVE8B3ewYVcit35nyZXj
LIYPxBlOLHy9QWkHAVOJxlrtgX03K3N+L/WjsXKSzHv9msCJCBfdswpjmi/KICwXZ5n7vwW1WBOy
nDxOJQg0AW+B78EORoB5aaUb46j0OO0X9V7QMixBl8rAA4H7TC8DBZ3ccwH2ILur3dgd5taHGOMY
BulhOB2YyAiI5Gx3RCQ0FJVz6Hm9mKiGNmEctU/5SFy0TBOJDdhSRzD0xgu5RWKPtVSU+yCeScfj
B6fU8xBIw0xzRUIIeje8icxwDvMt6BkNUfFQol2lBIkALnKQC8o+R6Zywt6zA+uzfLK7NSuwExhE
lk+NoEEFWvTYxKsL7H3iKud4OMhdXTaXQFrmo+ccJBj3r2b1CqkZl+FHSiwzgboS0cvB8OryZR0y
Shj395AMlqmmFOmzfn79zao7NpR6AZqmR8PDyJkR4vVS1nFa7c8oyPBu257MDkY9w8IQwXtuk3i/
Tsw8UH5rmjZ1BRUuzVQ2+iYrxu61xiVU+xrBXMjUUbdRU3R0XUlSmD51UGg9wjzmWRCKX9w43cHy
dzFyb1sYGlaf4jHVkxzGu1VmOLaGw2dHcbIuVRDltnZ5uehz3uw1TpOtPyIFMWBK/CNfb9WDWonU
aBl3JDDPH+30j26Ek8UNDr1ZRhx9mQjk8CyY0nqjmD3ffWe2EmNiMQsexPSynp27yQyXXEX7mc1Y
PfGWrASzkYdcb0Zu/R3ngsqKdfhXOabxtyncEVI5x3uLe16+4oPvAWAwezhxWhMRiFxilvjsubMr
aIksG6PhC63Vcnm1NmQMGXXYanaScNAGYqtb0KuaYEjd0KQhqaUi2txfDeCdGmujkuHT5N1qIUSj
ypV/dWMl2maXFF+OWsyGD+QSdyIDhdrhGFmWNq9fkXwhPHq9FgSio9VlhcXmo1XHNj2Yc9/iBR0A
Loeu1e12c/AApmOSqIg1+ugBHJshVA4iop7hqjG6DjQ5iYJvfWV0+xWkzH6DZ+0H/1MKfqmzKjq7
3vuNclyQ5JnQ54wiDmkA72MbnKJx9FCTCJzyogbJ+rD+Q1Dg/vAdpTMGizRXWKGICFwH0jcRPIG/
/Gzep1a6AI8SHm4cCXDtlp9JASbnGKxs5hg12zXXkcYjaKFHkGAjfZX3PT0V/WGC3NJMreV6/x3Q
d1NAnc44gXHeBdZLB3oL+Ey4alGdHvjE/B2kxWEVBWfJl6PNkVIWCZ6GA3akuelaSHUxvnQPQI3L
7HRYxBmD7Ho5CWDvi6h5yvYFIyfY3G9H/+Xdq/c7ydSewwvnlSjhrOIx903KpFvTNoYBPMlBqytn
PAa+XyuLVFu3drmCxnt9SYqEsjrpbZYo1Rwz3i3Yi32GLw71Q1+sdGwH2SuSyubEWrc4RHF7LjO4
wAMKD4ZL/5JJj/44T39Szaq+5YtV+hiOfU2ZGps1ARmBhJ7Hko1I3x04L7xHGY+8f2z+wYGjfJuA
AYnZRml2FJ5US/tGWAIlixbKo53Zp1yHDirjX/lr5DN4gJAHCNaySvg1LDWwPRvDF5shCzV243Wp
xEYBsG+lg+WnIyr5jQgDUBFZH2THZIr4eGdhdKW1RQlrvE77SpFnV/Ud8fub21elpYtxS2za9ClD
rW9WTEyROvY0CIl7bvDJGprlyjl+dQamksCNvJFvltZ7mLvJ2bZqLOayvWcF4aSDeAT+3fHqXJTf
O4Q0Ht7TfQZrzPvPjpG47dxssbINAEymxz0j61kJu3XxQORTKb5lDCAtrgqssVAofJnkrw5s2UzW
246/+gN6tJrovyKiWVVElRMZUZRz2tXsfgijsaP7XI8cmKNWEqIMq24NDYrdXZ3yHsI+7CWbeY7N
EMRo9wmmp9gZOBLV8pZsU89d9Xs65fwVPnCCR21f/5UsgIO1CWtGWMtYtvznby8AirQmpfrz+RCz
mwk4wW+UOr4FUnFOOuwNlSS1+cX2Mdg5gwop+LX2x8W/4pJZRAt0XcdmZMws2CPvLXfNrSA38640
u4B0zrf660nOBDrtp/cazaEjh4gcKMCvIoxSvrhbltN370HA5j83z0bHWWOb4MscTYxHTi8Q9TKP
9pvphQ5ok7XIXP2KFOWMKM2/w2EgvwrR90j5ph52/+she7TE35IXazUNn2gsWdQP/UfCQ39sPxDR
7goiF1WuRCSpKoDw4LfCV1q2+cu9vROb06uInKETBxC/Akpb/5Trr/NgXcNLIKtZZCUUgd7dpiQt
6XGXftUV7i4WADNRAOAvVh0g6LzUgb2V/gEltndn0szcWl9EwPdCW28383gToIzUvXlVV5z1Jx42
ejIyZObDDzAWGazH2W09dkyDSWLg4KgrPJrjlnLgsKiSzkNtjMhrIwpmRQxZvAJ0m4sETI2205xr
KJf1HSxEss2j6mbtrrpe0sv/C9MlTyI1U45xa/uDD9NOPGqQHvr0t0LYyzGh/AF8vZAejGmm29s+
+iDtdNgnaH9+5B9W8EPx6TSXtXG/tj+gOypPMzPUu4c/FoIifcyqgr6BhCfRSn22Dok1is2PSCNQ
Eu6Ln6bO0Qo4LM9xnbHXJxVDpB9sZekGA1huecuUdhJDdCjYcd3WnGk/LUF7bQdB9MWf+isckxJL
LoLn+H9OBrE15jtkcVaTKpIkNP73pT5e0FYT22R6Y1YwC8GmqmfbPtBmIbr1OunzSWm1DozyqcdO
L3T5gzkSHfdQdKmp0k3e0st3ivh0AzsejWcv8h2kHOikFYtYwbTxq1pSWP3B8SOVtAxOFmvzISzj
eivb0cqP+uq0cSSq2HmMK2EjfQBQijqgwNljXruhnjHJ/fO2DR05qcbfGD2BVewrTIzwKGC9wYvk
Qx8HWViNru7Za+5w/0wqnCP7zC4ciXK+91XsZR3MjpMi1dS2+lMWPxNzFiMmqEAull09ihD//xdM
LEsEPKqtSjM7kxqMHR8iA+NAgDpnQ3Xs+FklopZ7NG4lK4Vtsh5izGwD0TibA6p5wuc5jAd88nYy
N4nzqJiXxuv6a5j7ZLyNnI0t3eb4ynNXTVlGFBYshCoOwE18wJGtMEzL15arGl99aVQah4Q8EXQ7
3OjLppmyjPXRw6V99ipToPeMqESbMHjbOPYMHZZb6dyYtqaivXybw5x0kzwxrC5BLdjX5inlyWYo
uLaqB7o8AJ3EdDMBZa5fB/+RX8YzaMXyCfHve0mkIzKxf1/3+xpomPL1v3smuAvpQiXyUqstwQuL
BhjhGT5utezf+GK7+ZVechZAyAmc8apHgskdAkgfJqgyA8IaaFu/nuQex3TPY936LJ110hXOw7cj
hZWVUnlnyPsGgiWrXBWrcaRNUjFHj03ARVQn6fFJe1c6R/ZXEPgH9g0SnlE3bIkbV2v91zlbu4no
1iwtwHTtgYsnn82v0B9NY+LAUMl5qD6DvUjDR6bRvs+rP/G97hegroL9pYy0gsRebzXfndso6ZTo
xCuNuLZOOiI59ZPajravSuSPwao3vyf5Yt2rxuQKlrruFdF4TEjFFZTy2FGsvukPpGujz7L0dKLa
VxtCDy7GyRZFz5qHN/pW2s/XKi9UWQw2/CJLui7SzN70+Q/ZCb0N8Praj9yBdANxn4Ms+/QbrevS
rY9yvr4nU8h68V7lIjBl+4ZF2zi+X5Hl5We7uO6rC8X6hEqMIaLpqCxQpO2kNy1ChvZ+46NIA3Ip
QMC2zwR6yhmn+PCyBQvXwrF+e42SCOnfibzbHODqLPAgCREjANd4k5Tx7NBMKhJ6w1axXQoPKT0x
f0ujrNAKYXqp6FvO61XSksGB6Nxh1IITnALwWxzsQ+dD/HpIl8iXazPw13xBxyoWjaOnoRruxH4h
57YEccXIRCdmw1PwyILdGmkecDt6V9YozbaZqK1O/H7BmNk9wuFOv0otB+1RK31D4bYLIQ3/iLYZ
H5dJ78RNBdaR/eMDV4xf1jQo3Ns5GrWCtG84luiopQ1smIYRy13AQ0y/Wk/82T9SHQan8N/n1by4
2nOso477E1RTwnbh0CI1SkzRw0VHHfITEgWBg5MEUAYr0kEWPiJI7kA8Pb1iuEiSmnipnayRbEQl
pTmbZ3ddoFcsH4/3jxBo5li1Ih5mYYxSN8SQJxOOdI19gloHyNU0Ub/PPS6fab0mXY+3LLfs+rPv
CaIDRFzVT4uw2z764t5iazQLpK+kJiaI0gpg9IP6Ej0h8O6/UG4k+WMkXy0GsP5OYmpfGUcSmVA6
PG1CscRhUWlb1ZUNohppYEQNoo/CSIhM4z2N6HnWRvgjwKwJk6KKASjbsmQ1re4Vay5edVSJ+qT6
Kg3oXt4Z2pXzpchwnTQw3+bM8yIcAOckhQlhVHOKM+MQNm6rQpln2NpU1v5w9W/PeYnqWzn9Uyoe
MDiSh3AEHRRM+3tWOcOBpt8awpgaFGHvbtkdXBt9pNXAGAPw1ZLqFw3HrFRbqxGphkYzHhrT0spi
rP3TAp76C332UH8eDI/pHnTB0/rXJ9DV8/rLc7+L4nnqbmTeegFTfsxuQl+i33zjrKVOypwda/Mb
rRV+/D/Te0KOrxtnrBhpfKPW5/dl4YILMvXtMrzSz0m8weQRLhOtxhEpFBOn6z+a6o3cwqJjV9iY
/9fHcSyNC8ALSmknUKaGg+Kv4s2VLVnBNE0AXU8WlKf1EtuKmgWNwlI2XHdGv8thrwb6rX1SlBd7
pRb9vXsUcmMbVwP4wTejz8Pev43XnBIcgCNGx5yoM/0dyuLl27n2o8r/F6vIcbKzis8H4+FycOuW
x20ty84Y4Dht+Jy6tFCH3q0amB/z9Na75gRLOcCjkT0Rn5tCo7d3nsGx++PsYKhK3sJuSbKTgpvu
FGa7zznSmluK9+8eijVRhcXPmdVgEXkQRLW7JSf/lEf+DFVkUEYnEyYS/YSShzViS52F0CgBIfDA
nWmgbAep8jBp0kEfOYkarG4lcfIFzZA8XchE1p6qnFbb5OQEouaEOfHO46bImhNQSZ3FP8kgKJ9v
Ql6jEI/UZdz+GbWb1ArgvMBJzqNYRpNl+NP8hxwPudJD41twqQ/W1mgX0PsY927Z+LE6jR50nDqR
2H6BFXb80wwVnKm+XO5xYMUPhFbeRtHsShZeKrmxJj9RkfxF7VNIUK4AoiK650gnZU2/ewp116yP
ghDouDc5rfL0++dTC6+VI+7VscauOtvqYUnTPExltDNyVE3xu8YROOxAWC90QM8XlwX2bWLg8NPA
xkOaJIBneTIa4W2xNgUsCy2F6MBWZEpLxCLoIMZuW+xTmjkVdol0w0wQ55aZvOfOlTQE2aDj5+Yi
LbaIb1a3YAfPS3ve4p4RW/9OWsrKpzObBrJBTLM/m1lwMfSw+VxPhIEXfNZZFx6kg5OSD2Fwr1WT
c+f9oJl03dyr3/n6Lk9iMCsU2zh0QWGIjtHRSBvO86z2203ENgizF/lTIzoie236+7QvlhNosqrc
xVqaOso7K6+dv+FDhw54W8lZnSbugqaMRi6uStkIe5MwnflDd/fS+bTR9LdOTgJiYoyqbVISNOAi
l75xr8ljOMkIOVN0H4VG/pxymNlL+EX13TeO0kDjWoievr62wYfFxvIa6fBT8/noZ/jsmuwgse0Y
4+m76nuaaRakb1dH3PALWNMQr6C3fdEfB03nYZew3D5n9wAV+M6F7etxKAp/4/BtFc7wqQlehD7x
h9kZNmRiDoaLPDUEos/aJD9BorprJNl/7b5vDqkCtSekSryWkmEKlQDBI1Mwj72C0Ji4wHWPngrJ
CpLCEtoLZA0s4o+e2IZcB8zMitg+6vKZKyZ7oUUGHouBasfT5dY6c5VlFBxLEJVV7Ey2CcNLM3d7
KaAxBK3uDRAMUgknV2XRjzuKTa0M0V7KCkFK1lRDDWRgSKLDpJ2yYhaiRFh+Dn1xId7aBQYR7Sz5
xyHsGzMLjIWOMhpQoOtVwATNbyRUtY5w0rHQFYPQ+LW1C0grX1Nz3oJDPzCrH7niEUhImrOEW/MS
wsPeFnOap7Rvxs84q+nMGuVBVqN/Te2VARi1BmhYpsvjQTntq2U63RvGFGFoh4XOofptHEVfV93d
yVwl4r4ug/GzULLxSTadQNTEdGkD3/IOdlNXWotOLsorzOc5wPjI7FJm0Xfy5uorJjkiTfiMeWBd
fFK+fpDHKdDo1BBMsv38FdaXw/jE9dAgyVRT+lpR9QxgB+YhUJi1nyT9vijeRsN7H/+D/rfKoPwG
lJVljCz9X6JqQ6gA8RgdmjPzuUF7BABEcf8ACSk89lAPt+EcWQnp7mqMDPsJPXMvFK+9Y7kom/+d
QHegDwIyDbRIEPyBg8dPqMKLeh8mn4noZ9vjgfxFKkuUN97swqfe8pY8KoWQWwF2q9CHMGl9b485
5m4DDQ2w6w65s6fvPPPPz2UbMTZlK8zFmMhXw7/YbLevgqU0IrFhWSTSs6C9aTOMqhKNVhh5MAOq
TBUnJpQO57jv47cjCpp+Ph7iIK/nljf2XFlhutnp7tVJvTGTNLAfmM01tw4MqkK12VbKXa1Sr+Pv
IWo5nFjqcAujhUyL1o04HXBYfsD78JJDeOdV0qBXuAkYl8VDDcimMXw8q3duuw2APeoJ2wU7vjAU
ILfukzOlMq81ByOUcqKW89PI+ge/Id1mTYEV2WuqXLBdvXiIxux+42c7D341H1WKr8ACCtunJVsW
kFi+i/zI17BImivw5QJRrMxMI0a5QfVgsSFPYlD0On0Clu6O34Ffhvge+urQQc8pLeyvrYvGJrUR
pG/BQkXH6okGC6prnTjAbc9rfC43mH+fhc7QAcr+vD0i0taHtkAv90PZm/jkyHImMRaU3zV0+DDO
4X4Iskr2mc5OJMse/FpbIJ3BWL3RQL7S1bbeqmojVVFb7NE6o0u+mHl/CCDNgj72iWV7iktNiz1G
mGySPfT7CmoJVAT+UsFAGEK+C9hXGHTiI8ov2xet2T4JwErkfDgmuZlGiZoFzY9n2rtLpCofY4u4
cixRvbA1r7t/+ZFrhPAtV4Wn3tWXdC4+M7F25XH0xDPqfCapueACyfnb5jb4DLP93YGsYcwAqTIA
RGmQI0qQoKGoCNIoPTAvRGfYRsVaJGaCGC1H9RR2rP2nbucoxeU+oBrK42CDcqp9lpgJUe2TNzcU
clfu58MaqJSOyl1/ZxHmoENl+C04zO5KKYUHNyJaYGGgihy2XdGg1SgRvOczpT5zGSRIL5NCDnxH
t4OtV6q/tzdla2vylxXwlBXPr88rS3e2LuqctYqqZ055yVOG2YNIR7NxDT2Lq8mHsN+1OGZum4Xn
GfmQAZApQfeZP8iBp06eU8updQXzJaGaA0Vp7LKDAxl2PfiKZMdL0PHJlEwXcC9p9Em5S8crJfAN
rGlTAmJ7tzAzmX4C7kQpD+GOL18fbCLuViROovIDYLntUSSFEXKOQX+CzOarFagMXPC3uAWp9E+y
XCDgNsEvB+otLWIlT3IDYRV4RXU98uFBmrNkUyhk6ICaAOYvIQWYoeD/peD82l1uxSjHbOm0fX7F
Azmzf5dTs+kjkjkDNlgz6Zj0Y+gVKLC5VDqn48HZCeuEipxuyMFlefdgzDq5IKFnn9DNyNM0dUHP
ZZnbkr43iHaerkqsVb8o16AZFCsrWAO/5lbDezpfO3d3T1Sbck7N1TGP5mIQYoEzkgs3v1F61B2o
xSkQw9D8C5i/aBpcrri9+Y0qosIWayWtspJAATluB16Ol5IW4ZToQk7zV1M3T5bD0v/uglcbUj+q
+ugl4VjTUXRIZ9BxmS61SvG2ZrYLwuUC9XjfT9qzkE3YnczSqKZJYuhZkOkIH0z+a4NnKi/bWzic
wK1rrBqays+k+A2WYPPNWK7hkxbgImlnh6ufsMSpN2ATxOY9ys2WzhHBRK+JztrSIGwCJYwElIbb
l2zqIRDNCPcXBMXudhblar/krIMtt+3DOaeForLVBzNqOhbDVYEoGsWSoDwPcp/VtTWzpS0emAE2
tKskFHqnFWzaawJn6rGGHoT75yg512LdXpapLq86VmMYWRKsnDCLO9khDQJmKWJr+7uRvNZtmMxv
VqL5PpGRfnh1o5+sE0JD2A00d8CZcNOyGo6nqtFC670OY4yTevSG0sglh5yhw3Za4gatG4UBUAla
+pZUCkRrffYXSedcvA1dq0QeS83xTFMza0gMt9QM4X5F6wALHq2EJyTJUywqrva+fm7BU3QamF7Y
PAObZjveafqbq/SovJEDpsrYeia0fpYix+0RdWCNKX/rgG3ZXWd9iYBJHuoFBDptrhdrEBxIHQHF
1NGb+Gmc9ACOH3x8xPTYYfBk0tXEGfoWavnNxeQSlO1/yYC75JOQeTo2QwUlLlJDuNkTkHPlDoJT
vQYGJiqz1Ucv7dbkYHExv/5oteTjxl3SpS/G4XvOPcAUlE9ikgjOSXRZdiX7WXh3V537SyRsrcVv
AwiOldF25+8gA2IvtVHHrOhEC/JfSgczeMBljQoyyHIX8tqFt6A8Dc+a2AZOBeiLdeYIQbq426kW
zPpciNsGuzpAJMCIMuifMrKJWt6sraO+hrA3TMPouUBJXH2MuTb4RKclk13TUcAz06LYbti2LvVZ
4n86JU/8/MiMaHXSiEHFCmVXWuNrYfH4IaaPwAUJJXdF4FyyFAKGKSrHjOoylFhLOwNJLcsv4O43
fqHwgPX8sdKGX0qxjqmc+L/ugEZEI5tFC/507HW7cmuwK6RRTDrulE7Ocne2Fo4qW63Ki4twKtLO
XWOEJT+xuz6EXyZDa4BAmFGEUI9l611mxPrA0jj1RuuZWgA8MPk/9UJ3CQr4dC3+xCILIzLusZXY
wRM1HLR3ymfjSRpC0z9Ib+me5RVu7+soA5JPCAdwHSP2h9NxZ2ODYAaicAQZtW/YAliccY/MI3ME
Jw6D5sq/R4XMlieWrZn3AG2R4tslzNBpxxkHi2R6g/fsFD/ijQbVNnwYaCEzVpLmz0EzN8y41XfD
cepF/qJXXLYNU6LgKvNYY+fa6sWI04ttrTpwdh2hLG4+SpXWXlGNy5NysSolj5/Gvxqn8uemaVOe
vCj6V3Zu5xCwJeJmS5IQS/id8zuJi+mPw9WnhhLXuFvsrGGurAR7gQD/LtBp/0nSeNAA2fExaSKb
LZZx36BQRmroDVxq2TUgzcyg/Gxjhrh4okJoSh2dwqKxPPA9HwsshoYY9HgtOUBsMBAXbgvbhSy9
rbwdnPBE6kQXHA/YU2SYMDFqNNBBOmiuLRqsIhmksbQ36aMfGfngfDIJDY1bd4fVZBLxwBeS2Maq
L/30WwTZP06XpKGgODm2JuX+kVBQK1pbxvwRp0FE3wPl3bXTrSaz14T9B4/8uGCpeSwHPDldbqrp
p1KQCFxSrJUAXx/S47khjF/Rgq0+6fSGPqjsgWB0W+IC61WF0H2pkn++Zaf5h/cKWdpJZahRWIE/
sZvh+zAUs6Sk/oqHrxvc+o8CYaR/mEmwMz6FfYkScwqWKbMUUD/xweEPWOpjY3Y8l1KQs3I4DS+I
w6dU5B+bLaqIJqj2uSZk7mSiJ1seQkmU8EylO1m8zZgppoATJX3V5Vt9U4ozR4N7GOdN7gGEAK9e
r354S5V+8eRhVyjiVeKMvErHIQ8FI/2hwrcbGvEBiwApqWdmUvKp/2HjwBx4VJGWmP7lpCy56PFI
c7sbTrvKkCqR1LGBTlKIlFXAVn83MgmSkzk9iIdXox2npRnfOEGZYkD0hhI3y+/Q/04sMs/RNH+O
dbGkL8Lve8vfG+iMm2oqepVpDmmEUBGq0yZQAKQenTzSV1SJd4Nx8VSUi5QCyaNIney5+69QxZCt
ZMeJFAFrdj+kfYd6/2ZQHod9HgQHUqAhfCnfcmG4OWBagTwiAn5j30TSL8S0pDNIePIS8TRlsB8b
9rPLkq23a64eX3znA1rSvpzjBthimDz3N5qe6lWgTvcxv1nY/q9LKEn/d9H/nUO/mpF1vqr4Pqtn
69Urk3Q3/j4v14U/qLj/S/bPRkk+d8ofs8MW9x+nHh4PWU9vkUJtoA1dRz9xTVp9gib7HV7j5tin
IpbGXsHzS/Hx8hOXpyGh5zQyx9hsBPPd0LD/KuNQi2zEZGyNRFJVNWVWDFG5VIvkXWUSV6gznJwU
id2c6HqsPVipK8Z+zNjHMOtNVkKmaZVMGhr82CB4voOUaWLydLUnpR83muMo+o/VdSZq2oxIHuMv
KUbu92wPh1ZZ/EZUzK7jFZQgfFv8FKm/keFQ1RPYZhnSc+8mcAYaUO/8+ZeveaP2jPgjqfAfAYVc
vKcVKw3YUwMPdwsKVrReXqA7Q93LWG6O/F3f60WjAHfmbzsEbGOyGbiRg/Bq7+tfOM3WFlFvS7l6
ApxHJX0wN0BeDtJup6ZG6azubdHWBH78uQSVpcuqM6QeQJ7S39KbgWIr2iLdn0onPvGDYlW2urXR
7SZIbN2/Bdz79+NcLtERMdjvYWYCIShUTFw5Wo846X8vFl2W7lYgZRKUnQi9w5CFg9OJ7lO1ZcWL
wDJZBgMjfD/fiTTW46x2Lw8/Qr3PlFOvLSPiLiOD3NMQmZrhu/nfGRpaBoadptcu9bGErCZhRZBN
UT7mZkaOEE9Rwv0QVwHjZTI4IWtFmyi7QQEAZqgzsCdU4f0LeOnue+5sjJ/3ABszBVJ1kBgudzjm
JVGWgM3JU1jjPtVhhkpbmq2ONkoIRrqn7n4TTXRAWnqh4YRDn74XUat6Qo+4enMcFJ6q9tgHRvhV
VKtRylBd64KLnhKGbUUzeF8dhZSEocp7b2nMQ4NDCJ2GRQSylasp1wJWb93jy5QWzJTUlMmpmmqa
lYvPV2VJbmkNd/TtDFIXhwxR3DsSG6yc03EVjx/m9Mejoaes/Ezra+Yr1ytbJb49jYhM43OLX019
KQF64IKPAOWKbQchFtTdS6jsz3P8mTFJevu6QaGjvZLNVbm6FjYgajyzXJs4iPzegNr8Rllqx91/
0eWDrxz4BS6De/odyqR/OA4iqXmKyMVOtCd4uUe8fq6Yc0tIGXnEJ3De0bNovQQjA7csFgEdXpbD
aczJXusGtHnyS/4yLOnYng2OWfldjCc50ATYI4KVzQ/13uVgwleUl7EHoEnBh3121B0vEGOcAKBz
V+ENfqs4eDHWNWJfO1LpmsIkWuB5rpZQ9ULt6hUpxagMSWPWvWfvrOewMf3FNF5yUgrcojEAP3ca
9Z6BudQ2A/ZbB4gZwr6uWGgOfJzVbfDk7fPkEzKP4RIlxBJcmPBhvNsfBWzyTzjTwdAHD78CRToU
1P0ggzI33DI4TAAVjzlICkY24An5Y+FnBQREI7c2eA7ID0m1mWgRlpfKvBYis7eGh8mVYEG6+bpD
xB1OJANCDad6PJ4YO1KfiEHzkhWNsd72l4KTbD1tgYBF0yUVbr8nfDkOTnTqFT2T8b/FH3NKRXGi
s45IRWG2hQqy0w3bbzwee6NvX2l2DR/bVpv3GWMklhsbo47oZlcLKjf1cYBKX4q7Go+rR+EeaxeB
Prpmvj7uudE8KfukZJcewH3IULo5ZF+nGT/59qlfaNgdlZXhdr+qiy8gKnTuIpQ8JG8JZCrB9Jk3
u7/u4oLtjarmLOs1jRyWBk5Hbup3EN5wALNiFrpkSFLTLXe5w3SFolZX7TbrcMpXq04OnKf2BXnX
5i6KE7ysrQ646h7iH35H+2i9xrl/GaU6cN9VdYpAIFqtjB8m6A5VPHTPaXeKzpIbAXGXgBfvQHzo
FwzO2hXOXNe4lC7ro7/A+JGMyWVJcwSl6iYwyf5ynG/GFftrP8yiEmHQhMdNkwNEPMNGV/EFaoq3
P/mVINsNKUPOGSjaTxNLfHNcRLjZfH5QK/XQP26LfrHE84stf1IDwj2NVDVX1IqshIpMhlxNkg3h
mNxWtqgAsvOcQ/UrZ47Xd45ae9Qf1S9Yy+qOf0rhIB/1Lesd43DtVhNIVcwIMNdWvQb49gMCnVw5
H1orxaZF0y+CdC7vzjOtgHJdKD4dulnJIVWCP75Tbot9QCXkq0PS+l4BxxbI+MerEsSc22m8moxK
QWpnhZJsnexJhDk9N506ScTRlPAijBGjnWgx24wljVlEEOkhPWywtL6QuB/eKDm55DdiyKJHcUhn
Ap05Y+XNs2+SkuYJDas6iX9rbkC0vXgAITBsOf1/HN9uSMaWEGv60EAafmOIPTQlS7UZC4ehaydS
RN9yXEtEJlYB8FKNSkhGAN8nAMvp+TRWbG934fz6iTWMae71le99KEqDGwSog+uoMucnVSRizVZg
Lm61UGCQk7ftU7CdyW/4WFJo0GQLw6uFygn7b8Dpv6yCK4C9swCdRCh9a2DB1DLeF1csqJGu9luT
gDMAWEX9sMJPR8caKGsTh1SZ4qR92roeDDVrEJCQhQzD6AhawPMBFcUM7QIkEBsKXl+q7nk1C2AP
dIiHdQZCcHLAKsjK6Mpc6pX68jM/kxtXmawdb1Z194IFlpwwzqO+T9e6ldYKIBJIjg/DFICK6Dk0
z3TSJ4SttB7LuwsTAqduQpVFR5E4joSEQlw39qzlOhC9eGkcPwD51YtbOmVxRJA8Ki4THKKTb6kf
rgLqGzuKJPW1TWYuhJzHTIXLSaTu0fCjtHLVFuJ3fxSrGlZLbO3Lbz1VtYXt1kFh2i8/0xgYuJwJ
e1pcG/Q4m8PJBCGfTkio0s9Is1G82aYz85Tc2JlVsDUGz6LlSA+S48GTlF/13GEMUWdq0AbzBMQa
yFkVA5I1ImazcyeKS2XqNyDhSDuzuol6FwS4J/gDk4i1DBlsbPTOMrGTd3fv/j3kOrJjtRE3+8lr
FNLp4P8nxJKGu9qZFc5xjF53/zwOdvXjzERFSETmrW7XAY9g0xyFaX9ENwZY8ySix18yi4LhVcoc
9xMg+3nogEAUNaCnmE9MbSV/vhzodM2H6TdDA23tuA8lnS2dz9NQIzxyxnphd00cGrw+nDTEnbdI
BigV/a0DBt9qujebetJxhP8zIKQtBB26V8tA77uZOwbWOY7oTKelENdJ60Mk/30DK3wufOCKBfV8
fpx2BDTdwtSE0R0TTK8tqZrc9hKssvSBPL61s58wUfQe9XE1ATt+clnZDckwmjsCn2BMgGoq3YCd
ZHgbZOCBQfGkaZgEkGg0Lrc1GfoO4N/Vay/YvWCT86c7n376vJ0bWzLryN55FIZubBjd/GAtspgw
UWg7NKcfvP1Ud1ovQZ3SeXQTcopTSWYFtkzmMWS1ECIVyNUTUbldCCS3tyZlcT7/hH30eQ4Ow3TU
9BxxUsX1qbdMN2hvoklsBdOaHpaMVJylKlXD9lrP5ZBF/T6GeE6id2bw6oHBL9KiPJgt8wNBIvA4
umeFGgPjdfY8cly4Y+Flc5zAXSMQw55s5DYKTOHrWJolSAdNI/pb7tqupL8Cie8Z0dQ3MmjVq48t
3rjAN8i3ykIZGgyr4YqkBFaDKU35u87QyRgng/pqvGhskRFEV28RzyGVTJ9l8zGSqJkcXQOElDeI
THdqsdOVZ/n6Upt0jzeS7tRlCk3Iu/8cxNcxNNsHurQ6FundrnEvSNPeWAHFjE+tnBpQ1DMAiB3n
YRImkRDZUEyn5hAfZUYCaxs2tWugkKVnBP87Agzs89mLHvOEjBLO3cIUeNgi54JWkSjd5qcn31VC
yEWFMztA5Th6EtJ2wdV2yVKydv6hjevjTMK1p3sYHuAjv+IM364L+x4koId0BqYWbIj0zEPrcliV
R7G/nZjV+bqqU9/4jg1I/UwWV9ZV9ni8v5tQs5B7dQYNW80z755KSTNnXTMROykl57PHRdHYBXkl
LNiDgMAk9be1tZdCWX9FNcGir8phLzpcC6EjV1pDNaxQ+S0cSqX8XVdJXI7aQnW5wQuA4GV1dTuS
3kqBtlagJIApGCoCfPk16ISDCWDGbGTEeUo4ouyQ7oHgHE9yXTss72bIuk9CYOJOOxEagRX9TWhW
CJBpoqpmMxqP4jlQG9uvab0/Rd3EELI4tI0L4x5K+cGtnA4aQU60PlD8iAbH6XxMtjA965hITSTq
VNvrosbvqY4CUvYyLXUzcR2ZXJGujY6RcNH3aOlUFfVXCsEPIKrgu+eT6BFIHqej3lotpLE7MhoV
DzzEtuHDnKx8GQmsRjlv5XPFfEiRNI1sQ3mYiMkUvX6fw9h4gqgHq1ppKVEaYSG1/++1f9wz4kH0
jCtQmjNyc/5CBk84YQFdBsfYn9fL027L7gKGQLIS8vHRP690c3GA7gJmV7PnoWckhDykwq6ID8zX
xWKAxZrDr8e8dYOG7STC1Q/kbv8vqF056mVOME1xLyo9isqDR5VZ+hKBTPXeJkmwPKWOzeAObXyI
S9s0TrPgaPtRX5qKnBe+srLIe/g7334L4iCfllurB6hRPCgmCvQp/A36xbSlxb5eOmHvZH5zNEI1
5urHlm78BmOz9ADwjEXPk1kaCKSFri1hGcmLa4kpTkuemgPoVfhcI52IunP0b8/VJxeXVeXp7Rxn
6PWSRBRgpirM6iWwTOcKj+CZPAO65q7VvzU+vUOIJWaDU9bx68+I7Z7H84y8lSM5oL2WnJOnlTrh
Rs0T39xUMZg5Fo7JPAFW+SLn/WczbN15qcpS8cqUs33a6PHQ8u54+JoUWxPs/zxZTbYZMBgRFtCB
wA3ZEx6dwDz4ef42+DZk8cGBMnBSA26KWVpG+lJSrxqI5gCQe53ojjT5NfNTi2ha7xXOdzcvs0EU
PTqk7yoTzG7+7684+GYKRodlp5EdEEUawUuh8XFxHrk3s8PrVH5sFU9zzc4/xmKLWge98DcEQHUA
KS6NtghIgq/hp/09/g3R1GggEZ52YTMsSn3ILj6yj7fPH22W2I7AH08+WHXwl1f3VZj0eIuKQSeh
Mt4d/jcvl1pMoh+X5stda3oGH+rm9FQJbqGG/ULCAqCi4pIpEsM/4GO6HboACCwrNFGS1GjSvuxm
OyEIVAF/j9L55hybRCe0quwfKTH/Bb2QdxhCVbBm30Hn0TWxDICozokH7Wc9nTUEL1U4996YSxOh
0qFOzWfWOuWy5JBrNQ8v46tCgMgsrNlbqvUBujObcXdOlCGnUQiZZ5PQbHl3wUbafnQdWCzLyJI2
zDazhOAl6uchGQXB95UtEubQ84SBtqvo2qAtp2VDlKuondnQ+7k7vJy4bNN+UFSYeHSF4ZuDS/vj
HT9iBdLl0kA1scIi6p+o2h/kLK5cK6xAbnuD8Rz7GreMWBufQ1gd1JcydX94bjM2OZ2SpZz6k9d2
55X6QE3AzL5HEMnv6XlfWf/qp+hCPCLGTokyjW+RbeZhVkJzdCS9R8fL6Dqb33OSkykc2G/lSEWW
LN1Y01JyZDoGIxEq1mPtEx239DT1/vWZTe7gMh7M6vnYOmLb//F5BTwWOqQl9VXX6d4tuQBxW6rs
57YqqiAwEUoM7SLU+zGKRlHzfT17TM3vTB1coWaRSNUU0TtUB32IfLkdFQpJA3dMJXJr+4ogg3zw
9aJJRr10eMUTjQXwfIjUMzyy7N4ik6zttA2bUhjddU7AjOeU0JmeKIvFd6GaXVWYFSQ+O3vg0no0
yH9V19z1XOzWdBCIxWAaMO/q/y7riMRVkjYR9ZE5LCMPvAwcNu9e5OJFnk6dE7odvFiazCIthgPR
H/b0uaZpkeHBsD4HRS9/VYPsScka0OW+IAf5ZLyMqmPfHiPvKo8vvesVRGqDkuAwz7GNDVV17JYx
m0m0DoQPfiqA6okxvmCceTlps6hepA3KvYOhzNblGpSOu5FWSol8KJGh+DPPVmOf3bLFaW4auoXB
YSsMd8/i2cayRfK899rkIliF5KPAHHawH3VBRyTzqi/VfVKPEANlSveqSVH11gIuxZjmGdjbO0Cv
YiyWGKMTfvGJ+OUD77KiXUFfnNmsZNVn9n/xmu+08b7TZRkEC+d4FrGn1RjSJEMH636vXeQAyjvy
2Nzslof94iwMlguTX26FTlD25wLd6RQyUPLXG2CRFgfFUdJe9kX75MQPk6SCxplO49n68iKBNwlk
N95xojDq67Sdnv5Cy61yi8SjCIzqA7OH+b+hqrdMZxxjoXGr/oOwUKvnstBiUmE5B7aD4H3iT55c
caLKppRVOrW8GBp55yPsiX1q4Sb8Q7MbjxH3qVIe+hWlcbL/pFWATyghRdfRzbtPcb2eKb6ft172
IxVIzLNx7pZBStGAxwDLRg+QyTjCkapldFwLquH+H8HDwLmHYLh3FgGojJw4mlFmFax6UAzYON2w
wpffK9dzODCwd6TjC2eP2pRWCBF+VRGkhTodC4n+rHGsvW7kKiNfudLEgbROZQuc+RWlYJbW5x1O
Wgnu9j197dVXncw+9ECRdubfqDKLbLc083eDyAZUUsWCeWFmVJaYZLt8ofqj3oMgCeSE6US+aupf
HFhJfeOKm1T+0uzeblsy8Veb0KBkCOMB6236PyQo13LDRfhHn11N/MgbgW3lwLgijObR5kGx099O
8+mtOX0oEXHeTZ5RkMuQ10bsquqhN/AtY60zBCbXHamDMfDDFjCkazbAume3vmFTDf1ImmmdnjdW
Tlxot7tt4MfMzNGY+kyhZl7pct/NSjIXh38zQ8M0hLpLPFvYvutS9flWTfOwQrNgJmdcJTu32eUz
MfX935st9xNPPrFkBsr6NK5eeeZgyelciP9s32tbnEp7Jdlagtx8ssH9gI+XQWVrh0up8+Wo7vDu
oaLItTYu3NcRcR1gVvFcUgpYIqRGol8o/+toD6tUlgGDKAfTeYs+SjjTaMdRtLVpbc2PtTpQOIsA
X3reV+ob0YdUuPImFNyp1JZ650s2OevBCNS3gqlQGEbE7FmP8B5gtOG0ZQVXvJWba79Rnw2ytJXU
kHCrbie89bgOJRb7CHMm06gTvDP9nDDZ1wJo59o7yg0C3M4rSIvNwPtsz90lKb4eIGsgccGYsLuA
eraFF0rkuY/4xiCVw89SYv1URe/zfgzvlSB4Evz9VsJil15oCCybrbkcgtFD6cuV5dHHUd+eBuFr
bu3fGUHgiGQCuYUKimQiDlEZ+N96iCqWl1g+NspKEx61Wo8LtwxsZBwBZ71qzFx06w1TYZt4SlqY
CfKonbenB1AaSPKaeEeGy49C4k7DOevUXo8eVvKjNPNAGqyMVgDW5DV1/2bU57siwUDj9kHVn2cf
YJlNZlyIeZnEZ7V3Nk2v4+16teEVbz7LDltYFzfF/9wKH6FggsCB/vy0kxkY2AVUDxQMqVCQEIDB
SuvIYMOY0dZMjcsLw4KqvxoctMObReHGNjsnzAn86rGHJfBN9cGCo4MCAX1lE5S623GJcQA03pqr
uZkVkygmfR2uMuNr3Aq0Ns609Hqp+dZHcc4NeKOdeW8iM9aCeTozV+PTtrr6k7le3JhXsMiiEvDn
Sohv+LW2P4/DJAiyKLiwQz38HGdEHH72CovLfp1kPHFNrlRP1Z9m8pbB4ZW5/PLXgkCTVwnPQO0H
rqNHUtBV+Cyvc8uww4whUgPG3dJ0kmVyA8lR8Qmof9L9rpUN2KdUCaGlGh+7SOR4HO/LnOps267R
UupSE2odBX9TtDfD5BvyKgybfnkW+TmAnX5MmlU5/Ao7v/q8b3GYpUJj+UTi72hfodT9IwiN+PtX
6qZWlxTiTJZeFKOfPaxiVfZMWxITaNIkySjhyFgABz9qw8Z6ZJQAAgBaPcifhq2UHq5hcmX9CASX
9bQiY2v+EK4QIsyNv8RRrWnEa7tkN40jmvgDOApbmI0EQ3m7AMJvzUp/Q4J5E+Ca7qiatXNV66lA
Qo7GIwNvTdjYA1uI8Yv9fKI4xnBEF0o5YqwatHIP1fYBkGR5biAvbv7LAZ3ip/Ko89JXL02fGtL8
rR8k3LhIgjESzQHeLrxig1P+fUOYEZCxMH5nNnKplMpIjU5n3Meu0GKoMWlhn3GMqN3g1ctW/fZU
HSJskPLhdWUGn699jrv0QpBfVCfTbw3pL9xiHs/1q48ffkytxK0WJojwbBoE0+fnOE+8nHO+14sZ
/Nfajap4G/vOUSy0VnSRFa6lk3UPkDFY2bJ5bvEGulMKDwAAIrooYDdtBXixx00qw/+iM1IG4Avx
a8i1LTGzz4LMA4N9F8oWh0dyvU4Gj8C/2Y3o64znjyQCQzuK7Urb3njFyKq2JPYRkKzf8xXvcHz8
FWaxI96N0qLQJeT9/8xh5/7Ti3TwuKRHNfcgOWviiig3a3NZHYSQOEHgJG0QU32e6cc1NoZXLULv
77Ry6ZQvGD8IPiuRjPN+sG6F9OVXld5xo6dpu71mC/AXEpQbqO0j5tn2eiL2PrcEfhyM/Hz+tpq4
8apXqA7rkG+S11cP+jSHyHwM/f/FOAYLMQkhJHhRh5g7P60a+olxolO5CVmrqWtxA8ZBkI1zdXeW
WdyP9tKcHEjNMZsH1Hejxp6WJwqSpeZKfxcDFfwmrQfCIuksj5lqup8rM2hRECbTpBXY7Fll+tB3
VtvSh3CukalBSJ/PXh7bNr/DP8gGpzCA59qcNfz4n0HuI4SG2iGjnquDzLCQ57sveSAipO/Oj8RU
HNmj2gQuWVSk5jI10C+h4433Thv3zNeE3bho5Sg2yHpzsJAxRHy7NHanIrm1IvyoAmLXU1LeX/fF
WsK38DT+zvwDkCA/UPgeDZM4V8FpUHgx7zxSRxi0rGb3cxRjvBEf6reVd+mhRhbQWHTB/a4gbbpE
a02xtC6+rGvjuVy7UXlTRd0Wjv9qOv0C41apVxdVBCi5oGljsdUSX3t8xw5hRY6MNr8O33rvqve0
m8Z7mgOpic8sntOp03sPEL3JepaSPIgDAilSbqCiZ+L13WYYkN0MbhhrOyBTtcyJ/z6q2IqZsYBw
wIjxFNNotNn+cVP47ugkSwtEAYjvxZzclWW3Fzizbjje9J8TNCudCZcEx94E0tHxSzK1AfoO7GVR
NwW/jByoFOHS/NAKQ0SDBJxY5lmvFRYt2NCKVxwSPxzcOX1JLUbscVNvc/820IcbnOsQgeUhFJV4
DGK15ZukcH49rMyteUBGxGVFLZqkXuwwRmIhU/D8h7s7kF6BSvsuqPb+h2B6icb43q+k3NVc6rcg
fb+PSVH1J1Su16d8CAlKSMceTa3GT6aUPjiCWJ1L7ThJoPDYJotNmHcE06XIn6n0IJCvZfYedvJ1
1UuFGJyLy7WY0v4TG/kRgO/9as+cdbVzsgYc0N/u6eKpzcLyCHnCImBJ80qqaWl7wUZvb67Rcjwd
MFWb0ooPo9hXSv641T79zFXuo/AkJ1kH+M+mWFEG8riIOEiqWUH6Xi3wbf+nsxacWJBfNPHHgyck
bYXcAt9f1iPlx/aVHkjgFbsNkjjMBTRGTJp+Tgzwm5TpEweXkwhUKe2/VUtP5nwfduUTPQt2G9dy
IoSjF7d2pmlBUosb0cgTyVh+fScDGCtXj5lKUpNQAeQnrATQ3bb673q6HjShfvYcYjcgvEhKhWmH
fxLqgAx3FIMeLxEvfLQdj06w184cNdyhEI8M4kLGkF0uHdmFrFsAsMXF2XgwR1OAyLv6tz8OKMfG
mLDWaLchMQ2tBdKhTWUNOVl+3r/+fk6VKUOplWxVH+kqJlTbalZHOByIDFMQqQibIa4oNRPEwkJQ
DAQdp0su0aLJkF9iBVF/3kZiWF/aqpWyNtl2oij7HEPJQrzDOVFvzuYU8aKanSPMXw4MEWhS9ONK
x/81fGxc6JallgGgoWdSrEJ0VnP75dFnzHCdIgkcrSgyXFaVJsBYZuNTpJbQ3ilP93pWZsrLDq/p
Wzvh8JYul1+fuJgfHs2Gu7jU7n3lyL4fJpHsBvAHgwKlVHMNo80ZGAqCprrnxLVzjEhgpLANGKe9
7qWF1vwA1zVyhjZT/+2V4Kn4IRNdnVKaA1eiE73rIvoCtctOEhmOuIDmj1n/QMQ5AktwZVV79fcq
VFr5WOV3ILzNRcStq0T6CZG2qkWhicNLyCYR46rEdxph28+R++7KFaJD6AcISB/jaSFI1E6Mb6w4
L6FGPWUZuLM7gfDgLKpsLG327dSbrIjbuZIK/KTo+e21o7V2lVWgb/nFE2J/iCu0n1Di3cyHGPQI
yCj/X77+b/vZvGzfekHjA6eqrceltnSLNCiuoaeaAbnFjK5UXyJqLbr9Du4/gOoSXSGpCE4GEk4w
QbVBzC3FVcrnS8DN5aXq+aPFrknGHQbsOLx0l2cziMZfoT3+qbJL6U6nn4aWKD32GITHXzR+hIVP
g1daB5p2UJVIlAepDrQAEldDyb7QN5VC3ttnyBw3GCE6j0tNuJTljfpWSLk2KWB5ZnU5bgg2Yq6k
NY7eqMUt41Meb6YuxBIsLyfAfD9WugXggDUOu8MZ/rIq7ODJRtTjmmX4XIBIcY1H8uTd14rp1ZzS
7+slUWo8/D4a1/TW5Yf9ZT/AuaFflK4uJFT5pFdgjWmh1fqyLpPpFjpVZQoeoOzK51CofnZjgX9e
ZfheeO0qsemD330eOUtatVeDnPjBVNX5y1XIS17GeIJXAZ11Rw2WcGcncIClvADFBbIPhyEKwP51
xZRV/pbH6MS1HveG/3Ggari4EahAWttQtMk5T8cxJb9N48WgLGEXXuyjvBZ7HjNp65HWSr4ReY8o
kfPRe+dF8+IQaQI/eum2Mbt1nwgwN232Mejtw7aiZ+IlYwtmD0YSutLExhcXNoU9Eq4Myq2VXR0O
UNPLQP+MFzx7KNo8vSu5sCjfTgfVHxAkGrxxR9QbvSaiNhN25G9tkJR3HSjXPFpdeKl/8QjeXiPS
tkk2glU9/p7+Sq83i+J7VTHr0jKgLJduIGgjl7pCpOTV0A2E1rNTWZTgJo/uyoxog8NenPcvwVOY
HbZMcswbxCThtlvWdUJwIKzCjqgYzmJFC3RpD6NhbBiabqQjb+qa38AX4F9eQSHGbnLEYPq8/WmZ
24i6bh++CpVVYNqCDdmK07KlpTG/hoaHz/i1Ql/iSIaq3Rx/FfYpDFO5cKSjJsxlgFbI/H+NMjsi
sPTfYr3PlQ8d/r7sAuEyG6ftN30NDZF7PF3xplOmyZwi767s9y8YoPPeoqJ6EekWvqfPgUJjx4mo
aL92f4ij6RfPo9gBQcPrbueTFxjcD5xs1QyO50U9ZdFAiSQqHmqXthM0Qp/9f2WTdgg0nASI+kCu
Eavke9VA7wJBGQWhN1RpXo1TVZJ/8xnBRZ6OU3b3ckfQs0MKFtEYwUT0N9i/rRypjTnc4ACYTpC3
soLdy8oK5E3jQKTlET8m7U8CuI88GsM3SEpq3mhAGJaLCj1c3GA25r+3cJbD7RuZmfkOeBR8F0/b
hJMMdniGs4tD+zk2O4ZS2IVdxQvkvbMwRwArHun70QdZLCZjgfqqHSYit+Mflh7lb1Tz0F+0GQCp
hO68PnLijVVeJNJe+FC0LQS/BNk0/eWV7UZVrTjqufEcqAEqxAhUpkrVp218299tz7FTptQa3XKO
ETQrL3Vo3MU8e52mlP/oGDhXdPqOS97UGA6xSl/CO3K276KEfS/A+xQEAWluR1KAFXnDoT2Y5MIm
fBPtAXA6XXzxeo0rfKT1sHfEfiOf9eDHYRhNjwTEdGgUP3xmvw47xiEbKBFLzXlVRq6bKTGX2QY0
lQEBJFuzQ780jDBCDr7mlW0yyhRHeKNh4d1BLmrFWq0qO1+gjDu1JAeP54S1eUTEH9ndu/Lme0Tp
MnJIiMInTXYflPHTbH0BOayxoEU918oLcpI/O48/H1N5eQZ8q+X6o4jKq3GPeOsLlo7yH9vtVZ70
wvZJbY58jtPqtJLb3PGsfxog0eYAKeh+S4JPuMkRzVaEjuBRJ7vRDltGmDBMvat5wEQEVS6FLG2o
efuWGm3FTRSNmoU89GmPrPTmIAoYvfOg3fPjvSTOq3HelP2oLRaR3vzSHGaUSpIk+ovLyVKS+QyC
KoIOaw1N/ZcT618VYVkbtQe6fiUIgE/1GVa8rLAFJeU7vTa4NogjX7jIEweyCEGz23l9QpZxp7ML
MOkAHOJTBoF+e1VCVXIT7Tqi2BOE2npEmE2oDgfw2kfMhyTdJ0Y7aWFv2o5sn3YPCXFSZW9o9b1f
tSemNR0H0yX9K4GlKgdvyTDDAVDXk57zwEwI8RnRmvaLGIUqakZMmQQx73Co+Jao/C2bP185bLOu
TLjq+B6tL5tJUzXRmFwnDcrl2dVP9SqHhnNnq6cQfIDdc6fXj9dONSbLlgvYeCrREbcflhrXyxnw
+6pHxgEIWbrr+gVtWAogKEX6VDlP4vWvkHF7tbirbxLgwfpRblXTsdT36cdeE9ExZUHKyVCk3cNY
q01e3LXAknpUgpkT0VHn3+4pykk4Uz7opfM7GvzX82bfIjNHIUWS51V58MJqaXYZF2zEI1PMbKfP
rc+q+IXAe3lSsIL/2dB9ZYyHXYXCPkS0rDRPOOQ0vR4AN2SihFamWtOPzz1h1wvP6jQxHhXNK0FA
MTxxaLTkyQCw/XtidKCkI74SSlnwZt6WVcxWpev9r5PyrufWlq9X5csYrWscN0xbaZUVr9sDR8Ix
MVk9n7Ljq9k4VCl/lsEnlSlIpHLEKdDyU38FhdAw2urcw4YgQcwMYxzbY1Yw725ciHZ7RFlCYXPI
pQ522Gf49Jw1Vyyx1o5q6krfn++Ok40Lbykt/kKRkhoyNXnNhshhKSu+PuLu83yDiRzpNroxqxOR
Vu/+RdP01JSCZzujKaHy5l45vZHJ1VhmquBPZLdd4nOwVYflzjSkHtTiXMZXt99PBE1Gdn0pU7bl
TUrX/Xqj/Un5vVzgCuqik8JEHrHqZOe3sIEz+PyfH9BgIJM70JwU8AMYuVwbpDhitSQwxbWz9SgV
jjkkJCq4JnEFY0OORa6AeZit+iYcHTt7KdYApezteW/5kz4RrJlqYE5pLgUB3scK91FLZ+ITYsqF
qMpJ8bElRBoww36mv7uE+J9EAY9z5CEHeDHTkt5pFFeu2029v4F1hh7vPJXrwufAt2OMuhSpkHyz
GvLiLQf9eG+nJDPcht2b0+pp13zLjvr6syi2CIfLCxtTPWcQ0rajPuiV1joCeURmEKNnjQzr29CP
RiZl4yp6LRKUbW1tgSBr/VB6dqcM18R/Udj0NxZolRCCjOR/9sJAA0jiQxHVmZ9umIOV/ZWRt9HT
7Lp4r6q99PIDAM5RukbtgH2YXpf5XcjWROdgABTDICU9Wlx0b+Us9lsJcrTxzEr0nkZmMyfWhdGq
pbRKYTAzHL3zYiP/icX+QV+sb1lwsF9zOcy5GRsHAeOGjaxjInrQhSY6+RUTmmZaKKoWGp1keTOk
hyx8Vc0QDVESXcEb7DDA9avgCUuiGUhqa/ybl18vhK7wHOXw9/drT5e3Y+kkpt3bgQTSnE8kDzkN
IDoPghrT2KKES7wr2AFYsYWdBW2yE164C1Wb0wa23dRVdHz1tA60KBHmQCl6L4PdyROhXVs6X7n5
DBGMfPQmvrrpTgctsGu7CBotyYlV+Dc8BXXU1YIND6LtPzS2SCYH32N/RLYrrQ0+Qsp6rEdILYM6
Nl9MnA13v8qckEYzCK0bYGXWf5d86H9jnMjKNhjZjUtPy7sF3FhRwYO2ifzCJGIvjOWzHtBM+NJY
xppAFr5nIal4jRujthEX17F5rni+fWJ6B+sPZVox2fOq2GlNndfeFXMIARXRO0v8vcdcLdhZWAvp
BZp7JuiaJSjd06bQZZitqhW39/zEqKv7VfB98KFjEpFEBKcconprXF/z+7No//RLcfeNSoqAuHuX
Vh9553OXBeChg2kq3bNAUxMMfmFEO3QJz2ZpnNqgG7c+ESA/xIY8voHP/sikT9woexKkzXb0L/7X
D8p0aKYm8Bz4ZK8xf2TMt3/b+OiuLqkv0Gs6G326Ecd0tb/1cXw7TEZLvZmwudQ+iM6umtOWGJiA
11zYEWIMdC/yk2n1b39KnFkc/IYb/0wmERJgtOJbmnFBK1lFV9CO8Pi6Pg7tUcEnNLHJ6qglGqk8
/B5iUoJo+4GWLCcCGEowpVOtwr/C6/U8QKRMOXvwX4Z7zGxRp3/q7MQIgQVhOX2tjA9iVG5ksQ5e
GdO555nCmyuuAGGQrykMSo6/p0AOKAlYtN1AdxhIsMS3IIt83lWfnxl71jfYe8Q78OkjNNkI9CXp
i3y9Jvyq9EexV8tp6mj+FQdTokociNlJ97op4HgcGu/XZtEYf8yFkZ79LJ8qLRH1Elm300UZ2IrN
gYq8AJ/ks/HWIb4oHhTtX4LDQ/EPaLPrPByscPVj3fwtsr0uhvrStgdOqzVaWOy2JOlXu9N7nfxj
s/QX605iioWyfJ/OAB21nW6FjxbOnCjnX3m9/yUwkGTGJLMo2urnE2MKWcyiqORGnGNWuhaAkxZB
vo48g7zChX36F2WpxeLitoYQeJtOpMEnmOysv45pUx6ieCtD7KS5VJXGP9LezIDBxrjA/LHCwJGM
H3A+px6oRcuAMhpdTGZJjcmkLta//EwhmBcGSZEQ3vMle/xk/uDsAKqW1B+BFgT9hsd8i2zVuoWI
MTtu+JtKroO9wQ/5ddsbxLWz1tiBLLavoDWSJnTbNBLlcfNCpMyArIpwzsUE9jNS+UpNarfRMuEV
U7Sde4Xx1tOGV5H42skmgVF68d0r+ddW3zbBydeNUIxh1H4fjnyUo7/MD8PVb+jYGTfWJw3q3zNf
/zTI8ayb7mC8h/9sOHNRhNbmpcESW8NHROq0auL7Ps5pd3QvYMqtPmn38aYTfWPpOwEqSSIfz8PC
M62hd2HbAUfKRm1w079g6sFztQ+b9ntcJA1UHE1PoqI6S3MYaXvx/iBZIgev6wjgzK7KjiW6zotE
5nX0WOFyfWoDL2P8wZ00DdYRgGvRp5fOkYQU8qz4tedVUkwZeZ3bsxaJKPHBU7jk7mR0b+s7Zx7/
aAMBZ0Ajd2HmZ89wAVZ2siMw8Kw4nCgQf59czpq4++XbelKYeZUPKEp2q1qA9JUr41DrctxMzHVe
uaatChB2z1tkGvMMzdtBqVHrLAZaq9C8SBw29AhHltgkU3D7xgu0IIDiziwdUGSTU4/G+3N3tIN1
zzgNDE40dFw1o+AR4odjXpQeaLLX0NftpvdlVwfU9dV9qUZqe98sKeqaGgbDxIDg1j0g6AyaUETN
uXd1Lo46HrKIeQ/4hMLUs/r4aoHBd8bwlxLASsVjDKlM/QAJZHFYe8W6M8nGj1Y33p6euGLxx1w2
Y92h1EZAwx6SC3bj/DK7mvd1/VSaMOcL3hi8TmSbaF468wUh7qhhCDOnoqLcjrnhKvXndX1G79QZ
fpqIc1eEcB+k/R1Fc9XZNz1bEgpBGkd463opm9hOmv8tDOihk9fUiAyBkCVsr3RuOX4w6iLHpxqQ
MjBvB/BHZdBE2JWFRxFrUKEB7w1jqf6Ca6UyYVkxWtSJym2fNrNt6tlNJpMpatjDJMPDJS9zV/lk
5XHgl4cqF2TQYZdx7X3vwDN/+1eiEG3qfYHAxuQ6ck7B7UIiGLqrEZHSmdEVklSR17fyCfltbKrp
0XMot2QzdU8FwGQwPT8kVXQDYNCrzrHgjMWsDvM773jl90X54BKxcVYgqp9Nm4gHZZC0Ol+gcmRd
8pUW4fIf8yef7+1/XMHT5c44k0JGUwuO40gduM32mxu9emJWHh6pJoQPnUSyc3L4E795kTuLbg6Q
N+z6aasEuGuiRyNeG10tZHl9yJqsRj9nDPpiNsbghOMqPWdJawbXWUKF+Ij8+gzl9W5/6QS6Peak
Bjck1DPZPC8XZaoU+Bb7q6oGNc19v9bIrQ4f366t7+I3YLz7gcpJmUi0z1wqgx+X9r93+xlQz/BW
CnSnSGrPWQhoBTRlqWOSE1bP7EubQNK7ARPpo1/DLBJOHxieXY9YWkigqCX1mDmZUXwkvOzC8AYf
hcO0dZdbKjAkmAeDJ76CV3ueQAzFD9AuH6LEhgOxThmVXmTm6SP3g4YvakzpnKLQAlzfAyW2oMap
qROcixNsc8r5Hk/o77W5teEgK3D716biMnALwpb+DiYb3Tyq76nL94DkWY25DOVNtHGCT3xufi0V
eXOXF1ykEU84iDxAiv6v0bE8YR5H74qAO7pYy0jAGC4KyfOLgcuF5VJYEt3NbBrH5fMlyYlHo3Qu
Z1K7ThcfuECgDireCDUlI/H2EbANtaqzAsl9lM/HQGmf/1q738aGxVg8AP0ooYW0Dy20Ae8v/4yW
xcYkkEUfK0FHyvdft88Buk7xnWmxqOyewc9nnUfmDwoQi+k0U6pnnJqCRf8l3nhwXsJV3RLnVSK7
V2xI4Ajn8sv8hgtlOPCCMx4kDP8nv9jJs837HNGzDvd+hxYuCCAQ7QT9qbkigt2SN9neLBAF3dSX
0AHNW4BKDDLwMaYaBUTYkowRSKF+G2wCgl7kNNsqkwtZLX3GHCXzvXQGh6xdMtT9daBbJhb8QX2Q
TWpr2pg+/Fc7tD76thPxCAwd22QALseWc2U1wGD73d+JGcu6RBpQTzN5P9VoPgqqz7HPJ2epenIW
mLE0uRguPiQDXAUrQa8eLb7YBRM+E7M636gj7oHHYBCOn/SWK5fFzWjGkhgd6kXKEwglEiqe2ErE
SEUmZ5PoewXtBHVWD91MQwnjzpFnEYU+CknQdAWWAaUNmtgxet0QzGNE2dwQDurOVkrkql/iexdu
MbF4XhXL6SCk86Sj225iTX26Q8E+ZTcq2CG5MeFnLibcXTggdDvcpxEwrq5uEAKxms3P0ch3eYn4
pMk3T3PbYulGTfQnyflpQbfB6NxbqFpBpK9g1HBkkU7qGmGTK7c/EQknAPxviZjUvqlFoL+rqJfs
RgJwvEHuSMqFc3jmrrP/SFccVNRGMfx0OW32klRnsrMZh5x05/fxqm5Usdbz2BjgH2j2fkT+/cEz
d0NLFKEOx/gYhWpndCoFGUlp2hzEDJrGUwIL8W5THmcrsFoMQkW2DTVDp+d3dRIU7FdD6Z/30W0f
9GX3KBQRCJw9OLvG0guvLlp2QYF1jIk+XQ23P3oUFJjxYWBPVqYp1DdeqYdosMF34PDECmdn1WPS
paErWSsPEa077QqeMqGk6ISE0v+wLrJSSdCC8mYTGlLdWE8OQCFFk4iia/wk/wMk9YV4KWEPKVW1
+5kb8lZ8H/z14i27EajA5w+eg6KhiVfNaJcybMScaYGzQdZFlo8zOVdTYAsgb19VktwboIqw5f5r
9X696JyobMvC6MJVmL6eEsoHsL94wrtPlduTr4uDtvCM/ZVMpe4t1O4a924KpZJoV1JTbrlxy/GZ
BuOf63Wckl4YuygT++GMG5WMyFOHI9Hb+rV0ug6IwGAi+VmC0S82tKO0bIb5RrPceE3Y2DZvAx6v
0a0yAZDgvMygmDc5c4l4twhzcIfXZv2wsx2Cy/UroTIkA+W42DKUIQ8MfBxdyDwO9JJbwgSqWk8M
vJIAjgINhLOcdvn5yK8vhy8g1NzInB5bgwFIvmNCuViOIrjh1lu9ap/j+zmtMCeI5HJVo7CxmHhi
mctgbZgy2RSpXr+108oiNApnn9bIZmKqU/OjsyXbQyWLnnzvKMWRFYfQPCpYQGEaiq3virsfVxEx
H8U3BdfljJk2DHI4Qf28pEQxhRrDIBQMyu+KXuTP/HVUe/NpmKM9wf+EwtHkOyutNY4uIZQrRPie
6A/Y8ehN3thYF8WtrB6gRHqHvYQikhPIn64afkgP5ypC5mEPGnsqfioNoWgAXOeF6sLzFCXmfK94
dJOx8SnkKWGR8f8n/9P1zvSKJ3mF45SAsnIB2xjWNcKrsbPJY/Bm384OoV8kcCFBzSTgXRo5um18
STvS87pjAgI31fmJIpnQKqaiRrdkJRXBROjxa34CdThc4t0MZS4onWrLPU/dnMt6aHwodK29R3pM
uo5kQob6GwfElPQ8EmLcpgQy1NLghOeFoCmgNNDVsL63PbvMVG1XjhpMUeXogRoZCAGW1qKh2t2w
qcKn/dm/UkV/Qg1gKDQjm1kz3lPG9v94U1WLS6/pfe7Tl8yDqEyTNCyif4hg9JT7GwH/+mFp7Kxp
fmGTmC9svGvO+EC7yBugfKPGlMHf4VR1aZzpLNIOrwpBTX+ocjkKvn5ZMuqCCdCMNR50tOoNzewl
+p5+67WE+UNieeYK66eHExNsH0iN0dndwuBebH3kBw1jel7isW0ZVBajXPBAGac58xmw3ghUFzZU
2wjgh81zFRLtKc0NEvcyg9TeiqKC1j7G8gqDuvs9gpr1JusjO84yTStY6A4841hNTv2xSBI8cooh
esQK51agRj/+Q7IS3hi+gUN51SQPzzQ1dXUuODM+JT/w2XeVE4ihbF6+j85B2CYuylPzAKgldYB/
FF7+Lzv1Lz84hhY2XMv5EgS231lJQqtPHV/X0xsefX31NvH4UjnPMcVLKp9Atc2PYlkliz4qDG04
HH5Mo0LL5gXWEP/zEFf2y8G7rOpr6yI9zTHIUuQzlrsV+IXIUaO0693JjMNFEHGbNRyz9cOL39Bq
iV/qLBsoqfnlW41fKkLuqDPQ63+Vwhczh71wTJmZIdFwivUH3vLzQZ6J45QHRUADW4WBP43hFfJG
6h4masjRSpYQ7NYd2D+yR6RCo/xcRPggrHbRSnU55SFOFkhAQjbEDRfhTZd5tHhLjGVUHbVz3Se5
WdCAGD2x6O0Mm5U46XGoE9TDegQU4buIMaaJzX6D3kdx0hCP/v0BqhSs+KTbAh0QGdCI7JO5xaSb
5MZdiDnyPVO2MwXeRdX8/tdgdKhj+29a/HJfKVVCTMJaqXTOOceysuKHO+H0gE+jyltmeP26MaUA
JJp0JNxBoUKoRZSG/NaW5I8cnWLi22dpbVaECrORzWcIlSsQNvm5H7bXzQADfS7YZAM47QMtfMkI
by+3/dBcz3y2D2q1mFZ2TFnqVvCt1uNb+5WcfcmAMFHgyFHAVO7oMFsWb9qU649xDeKmDCyRaLPc
jZUTVZAz5PMAONqIg6SJMqyGJAj8KmAfaoLKA57cgN7oN8TsW16BbEkn2C5Lbl9hg4ui+W0bWPyP
KIYW45ktZuPtG2k5v2tZx7vKY3oFKs713m1lFOeXrcEa1XWzM8kZaO0115kiTQPrxtVhqBs+Aa7w
o3hyMbLd2rweULh2Zsc5hxWtZZkxQ8UTh/V9XYqz3Kgd8jM1gWLp2pACnK7HVM7hru2z1hBjoTZF
kBCiwtfi5b8uhYSFSoEBJKwSYaWSVtqNdclSt5UpGhw3acm90193Rq4M09GzTtjoO9/rUlLH82bQ
cH2DMFNN5CqZU0uIyiGKXBZKiMHQFKCMpRiX+Z9pflNBukoXnQQnaIFiIgDfXHBbJnaEKTxRHqLz
GYNGGvpOcYzqC5T74B5KLZdqYx9kCx3BxQzgBrTyj6bKVr19gcZKicqrKrKiIaGhghaOA6jyP/eQ
pydcH6cSiJns8d9uvQcJSYkfezlxesseybYTQHclHgT3YxoSFRO43/vVjn3SmOYD0Dp+I15UcK9g
UPFIZpfK+eivfKXThQdKrjA9vTHWUlv13J4vJbSBr6PfrHVbA4iH74NVas8Ma1ZJlp9dTow6jiz+
VA0UJjXRsqaHI+BLqxrg6d5wFkleN6LONv+q/lSVokp+i1A01fjO2p2pQgElLDD6UMa9xj4JXCf4
fSCq7KCWhjIic2JSnhFhLNnozQb1sq+ZlC1vRi3sTcL6qDKd1U3MHhrw311u+3edpfpEsJwwzzCV
zYAOSo1R090ZlHY14H4qCanrs4RZg12cihnD+6hVx9bSKsugSb/0ehturoR3IV/J3KRPz/JiNuy3
3HSYisxWIqvN7o3VP8RISi2NUWYFaEYO1DRkaC3jS9v87aLAW9EngzzIoI0s32hdNBqUr+81+kc9
PZash4bCwiVIaH/kqLvpZXSnccadNsUgOLSlHGkt5AlLmDdz85FTgbBkLWpmFs5fS1vxGlnCMki/
NJBfQpfTuRgKgqDeFoFb731rx2i/DgxLVd/+6No1pmlKN1szkOWkns4q0G5qApjKF6cw/fNH2cme
s1UsVJnyezXip6Cih9pQGnU8KS5QJxKSdILfRl9R65SEutPkp8CLsePVNqZdlh6neb+algaveXCP
AL0Hhd/hqdmw3GldJuVSEodQkYq/CD10UHh01yohrKra3qwY6uX00DhS0EApkdRUBcW0GjH5dSb7
95OQvkLAcTB/xv75UAWl1NWZmVhcH1yhH3WB5CObyAX/REWB1rodJ/OePvZdyxRNUAmzdB6ZW6yH
rGLCVjPv0qqJ5ckyfCgE2NO5iJ+bc09Q/bfmMBUCpiRrkwgHPniRwLo+0tV4wr2HpZPAnwGKqE3P
f0P7vPZdrLaF2GvVQfgxf2uCVrBZaNLYggu+wrFkK/sggJuAmfrkwnIPnKZjZqnhKyJB06gGsJox
qv4i+qHDD+dwObBRBoa381fr2gC+Jv0tV0NQL/K4rul7SbwH92AlSpWEi6z0yGH/MePCYu7Y9wan
0O5zbe9wMrmfb2pKJOKYOS1LSUCHMes9etYtlSb+cNwAt5QAd+OifXAugJvKWeMNjzw2JMBuHWv3
mHeIeuxvR8CF7tALqL8YdNdsmNcHr+eoH57XYU+jgu2mbfhnqZbUZGs4yG+PBdYJoEnFegsvMJSm
mX1YL2e6BwwZB7tttsN49s+XaNn95+sxqJsHIkQHKJsNvixTthUNZG/JbILhItbsEat4nQWw9ZK+
l7ikrJL7brNHJm6yeJaslpixecdVVSYWF0CV4WTB6rtqnWKgqtIk0x1wRJTxi5b/TEZGf0oSTVl1
Nob0ixBOZ+ULDIEKKvHW4pLMV2jTNwhkm3adRqmDxjbrZAFRt8bd4DwjJgtgZZPTE9CiQFJrtcdA
xBkujHC1UMkKllhXGH7oQWWDO7jRk59bKMd2Qmg0mTtp/4G6rtJk32ew/F+IbmYORRzAuwvPoT8V
XRwQubpco+ndYd6SSDUnb6BAnrr+PPvETrcxCNf+RaL6+iDxK3g4n70j93wOC2bOXDn2DMjww6YD
OWjcJ2vr2kYFfAP/MsUhmVhlUEkMNz+suE7RXUyftKcO4/QPcDOuy0uhfRmHpucfE1c627JzD2T2
3OJl6hgQxA77rawOVlQItUXHh4zGjx3g9671wu3bh3RdHoLHsC9CNPOPzMh7LoarFVuvGZWOYDiE
md0jF2pqKj+v6w4MApcJblZ9sZQ/9J3ETLMkOawzGKm+4eBGkR/oj3uS27UWaZ8JviVHBb/OKSl2
gm1Q8vblL4Zv3biNhys6LUvBPybhbErtwMnulVF/ieHdKikQhhGCrZZq+POf1W3ycwuadpQMPxIj
X6/DLzPVQBGCIepHyZBJWW6KRcAI2TJBSDexC1+xT8DbUZj2SuhQnq4A0SpwFBgT2uOXpr5Av7bQ
b9TpClVAsLF4ST8JdDtf/LIUy0rfDUfaVc/KdhTxAiKZucwb4+nvEw0jPeXbkqKcAN6AvwrLHgC9
eeHuAAKncnEF3w0YhX+XLyVe2SnxsUjJ6Z2wrtAOW/xLyZxHs32XhkWUcu5yjyPn1PkIn7+YQf28
UYKlY7NwxqubxGkWCsg/kESsLW2nGduaMQXOrmG57YsGomnRIty07Mj4y8wRaIQehwB32IKqS7a7
LbXiBGpsSQRrGoHsrmaKvfl2RAc0ISXXIjhn/pdN/CJ51+Oe92Qt1D3EZG3gIft+BXtm6DfyGCOs
aLXp+NSUcdQ8L+gXi69qlRZOGfB+OptlORbUD5frtLSFIBEAE9imbMTPRWH3Bjcv4PegM2EH/36T
pG070c/gs+P+FnD0HGQdw0RqcaGObHVTYL/p0w2qUi6svtPDgeV37sZVjLGL0wa+eQBRlDQblRvh
2pLOKAhC301q1ZL/20xvY3vRpwhc1104Kx/Y/HNZh2jFROq6SEbpxxPS4v0w/U3S4DV35ob3gOh7
1/RSyA143SlLIJAKrVtT4eF93+4RHb86pnSvJ88J2taAqCL7Vm4xTP5z72cdWSdC+NH9ZMEG2KLo
F1ozTmPOWn7FcBgHYSP6QqAeWEcC1M4JH1inQHbbqOWCDqtWWG1TCBcHQpFF5yh0gEhypz5Bx9V4
H1OqIQwL+tOeiAWMGfVzhN9FBAZD87O7GZGEcfj3Gp8gDYidXMEijGe8EZaDIaNDBY9AzoU/G4ou
NcpJ++sDREXS7+4NYzLZPAUe5MyAUKG+93OL88yGYjxKRaTHn590E2O2qJ65Q8bFYQsvsuEuK63c
908nTqC1n/J/luwvhLGMbWUpagwPEVHCQ1vrxrnfAcohscLtlLgRlWNEN2Bok9S18wgHlNKtGad6
juDG5yVsZsLVruh74aDRCbq19J2appjyXryKtAznukBcapyT2XRP6Mf/a3GuRscMvODDvFAGUDJ8
D+6WVW/48rxfPvnkQu6n41uvkX/gWfar2qSCrBUHBIuOl4dFvJRGdWSxKg/o/+PJbnGAch0En0Is
Iohq6DPoaa3kGaYy9s6Yc/GMyfkVmiKll+oC/S5TcY1WNKSK6jA9cxJW+I4U9aG5FYT3gM75cQ7m
PULyI25qqmxwui/Cbtv8N3c93SgrJ2on4sDrzSnlOAWYDfG534LI6I8gLpabp50ILTb+aQbHYRTm
m5TRMIwx0oRK/pSiAwprsjHZYP9URgDp0bOFIS6EHQNDUhI1vq8XyCi8drXVWOuz4Srjvahc5QQN
PSHw4+iE/xItpDnsP+BTg/zWbV2T6iDklnLkFShfY1AtLAL8MRSbipktv4DXv8Oytn5LTAWYznm6
R+VuAMBSVTag+F7y54xaXt9fMtzdUmB3sxxXEZzdTBGDrkoFGjB9mzEmGXJQRtI6VB2uKDurKjzL
vPZyjWcszCwsg05W8ru0MSBfAqw53OwsaZYX86Sn7r6HMNEZh/HlU9JOjZBUH3AeB1RfHDwb+YR6
JNc9iD9cgXLWVnMjJDOL4FrDqAJIwBwtr15TUJl1I/3bRuWFk6dnsaLlTI/aeAiN1g+edU62h0n0
TvivCKRHMZRNQ1ZKq9UE4YUq4Z407pbwurzVndwtzl9hE4lPQDhmLYkuhm9PSA68L/KutRPoPw5E
56qYgpGB4vHaKyfU5At90AEUUxA/VmJ0psgFMGSZpp8o7qX/Hpe9GdNG+bNZG/nKaZ4PA890LEZ9
AO9lAgKOoesk2jfaTWfhoWD0vPTn9xUzAOvpnvpQ70PJvwHzfZP/t5NIPKRHZxNiVtaT4nvUIEI4
Ki1ciiIkow1w3h5l3Q863VKUN57o4LnivekUK2/MVuQUZUxAW9XyV+qoIwAIzy9QMOT+XvYihfPK
FzNVxWyNZex+g/BdAA32v0UVRB3mpG1GZ8Ij0rQsARITidvai2UlHBdr5ufBGUBGLx/6ELrwjURE
I7600INe/h5Dmecy1yRm2RpvtHMs42wBzxCSvQXetPOTwMxd1vEBc9Zik8nTAeFMMjdMjz8NQqR+
ABldFZS/1F5NjX/GfoeQRGdaoPVQvOLrpmYaDv4UzoYdAg5oNla6PGhjzVh0UbnKQlYAp9lOFXd9
Ib8MWu7rZ2Z2FIn50o/Xxlkk7nO7iVAero/K4AcTvkZAIehZAc3sSdxJtUlk4Su+IEd2/Gj/Qwhm
ncveK/Vtugk2hCh2h5tgrBqHPLa929X/Jm6KzR4xd0ghzPThMjYSmTLDvOsf7IMySGPWGXIOmC2h
2xeui2LQSqkjWZs+O3PmbZzlLSR+4wsLCnrhQcOjDCRkEv6Y7RdksJB3QaKibrwqDBcrloTFNMvG
CiPcZu1HJ7z/8vShWoUhPmPNzjdVCyAEtwp8pNXPZjX00hKkDUxgMCV0qRIt4yot46pGsylB+0ql
0ibVmKUXPjQXxPkV3W5i7LHGYvXcQ5qF8Jmh/cv+EnoTJlDkQk3m0krcENa4MYLzeh8VExafTuAz
6f3MOB80CGiqe8uEbWDHa4wvMPB+vvHgtJwDte4tjqV5zv3y/34inLVRRoZWal8wQVLviuYxquFI
fU2P+IlbEz41wfgpIzaYFhPtbe46KZjj5U+VlD+BFfzyeiQFRhj8xdsPqgMr36v9w0G0qVzVJetP
+WNsl4qmMU2rBPApUYpEAfqOJ7sJFJ/h4a9JFgmUeYW+Al6y/u2HXe44EE3d56i2zG8TRKQRtcTB
AjBWEvu0riWFxZ1B9OizhXHv7u1jpiW1cG/9At1BNCg5VrgvTZlFIYdPCbib7K5wI13wQqJLofk7
ClZ28r73EjO9McyvSZL3L/Zg87eVvWgDCeHtQUjlwX3jOHigBrXAvGANFLqIsuhMZL9c2kWMUWfn
adS5uhvP9dYC7siWhQ2RhZ/P7wOnZ/ppfxb6/qZwW0EGH5nCAQiWyz1gsxR9rRV1VIbc+in0K/WZ
J9G3Dhy3FWrpKNvsTC050tgrG7BY3RHKdIqPKcJ4pthv0jxeehmGfCS7PAPkxWubPRGq1LJWUYFt
Cf0veOoXK7c5c5EFIfo1ulaZYItfIqwMHRtSBlm6+shQKy3Ql+FCNInNUQjldx9wSd8pEUn+4NSu
rudZXci0/FmICO3NpSLFSxaKolGyLe49E625Kg3Bdsn74LRXIBRm1luXgZW09rSSZuBmA/jRJdv+
HK96YOkTWXODE+LRXCVuBP45a0oj3zrYx+lki1wB299YPsewgO21GjoXSeQciRKBDV6tHvbG85sp
jwQ5RV87ZDgQYT0PVq2H3trvk1+V6PyzAETR+FXVdN8O94vW3GAIeqwjyWeIg/PbjuZuj/gUdONm
jx1kVvfpbxQEAkWRM3BYOGVTJh/w357kBhKp1EniPepQ4BW4G5wtEW1S6ZBHOmsJM7vRr/zUJjrF
SC6KhC45j8ULjOSFGE2+m5Zd4hJ66xn8c9DMTY3lPLyp0nDmozNiuj12ahqbkvmgyF5v8JOTiliF
l4D1ImjGX1OUI+BjpClJQfq4uZbm7PiZHhog3RPoQpym4S9MIBIB/LebhTutj3en6576oUAvDAgj
dyMkZnmdiOZ4nRhgqXm77jGndN18CytPXy+i1q9ZYDul8Bv1sHzxCsmAM8z5LYZnP82FaJmM9GUV
FsSNm+QRYZGI10Afwnc47/tZNRGlTh0OBxDU2EbKeOIEuQQRvBRoVXqiizoI86LymNUQHTTpVXP9
ZqeXIjwJpJ5ZHeVE+/bK31eu+tq/DI95rsjvIIcex7yj1B2Tjb79iVbsdxuk8XlUemuCwWXQGFDW
asBm7hCxAACxticXZb2BY5/n2eK+sXYMkg8vBzxjqerizOZRnavqRHnueh0DRxslJNIqulQWQxbe
kyQ5uDrVphjmFWj9tVaG4sx+23FymctjZOjAyqx/hzI49rLQ5tB0KhX9NQ/82/FI4IY9ajynvI7V
e+db+VW1D77PxqJPColtMG627r3BuGYBJiUIIhAQgNExq6yRupeU59x/9lP4DrsBEecqkWH3LvLy
4j6S4qB+gHQBFgQ+uRdQLogynK6W9PTqGTuNvhTbgxCaRPga/1ILcUraaWdeWMeqinE4gmR5UMW+
JTdlmsgAjniEAwpB01Pj6Ga07t3ow8fqEnUV7dQFbjR0VJDyeBM1kZ2QkTILaMtX0QlBp5R+Pu+F
NrkxwD1J9UQH32QGz3YOtfqCFgkXsTOWXOPS/SuGtX5knnCTUaqD/n0TQHgowcELaIpQqpXs+/GE
TKhkJvXKHV7DJ9vaYoKaB4pj9GeT9ylLnIrFKcaBhYwmYcd9uss6QtYeZn+EFBdL/bBhQmrul3e/
oxU5fEs7xDbMVtK6pcsSOR6A4DCvBAN9TL8QZh5Zyzadfyjzfxg2ySyGiQij9rqExQ1n45mf395e
JttfaCmjMel43xa3SNgSPn+6afnJjykVlWqo3GeuQze0f4O/ep0WcMIU5n9RA37GzJMdhRRRxBKX
r5kwovbVQXE6hjYyItAUu+bZtBqJU22kvMJ6H4WbuMmOpysMqcUNjW1ibqWf0SNgP9yk7yP6yoMY
DFRZKFmSe1Hvq4RAQR5JB6McEe7vclGHJEEgQLT/omDPuopZXK59OB01ku//daD5YbhyqFFZxgRM
KxW10f6/VFmM3Hbynx+j8iP3Gvf4mEnUMzxrvrmXdGYKSjTq0zWswvtjzP2h3RC63lYce+LD417Q
1Vpk3pGPFd5B5PLI+9Eco4L4dpAfioJAJVk6aCpJ7J3XYiHTv4+toUPVkh8zCYPORIkm/EnsMWon
uEdili839BCi7rKrQmd372cAiW46m5iOEUB4jowrZOrD3gzPLAXP1JFypySvddriHTsmihfA0oOL
B9DwClvYbHMaagdwxbB5AttDnzrvcRNp8V7as+WJClhrWFoO20UX/h25zNfJgOAnaWeMC3eor2Qo
zf8YioOJvUGbv91JJwZI4iF6+68+0q/h4/UcSesh014ix90SEbGVWSPmJ8wET7Xu41mcK21ulgpN
/bLn1bFrS+0pBdBaRnIu9Z0DgH1ifSKnBjK/86/PCom/gcKpLODfEyKfwmsFf+TUdriV8qTYzZ0T
R1dcst58RYNpTnaa7EnwLYf3TjAH3D4z1h7WXNSwXbMUZg8Ru2C+ISaGBPya8yRZti99gI6OuNVG
s6Fam9IJ7sRcy02E4jQfeDsalo/E0Zukrti6YGiP71aAtU2H/KIpvDhmmXAPHiATPeo0BylzobPu
bqlCrcDFKhzvRT0SbKar2sNLE3XE6ZUQG4LRn35eF7VlqshXade+ZPkadW2eZBhq4QVv5gIXJFe4
+cNr35Yd+GadbJLRRj6sj0ecKtOO9RPXd9/VYhJR8XISrCia73LghP81H7g3jt5CkBPs+516KAQ9
X3J1qzhiglHxpQeeUTis7rmWERkiw8Z79/GKn2EFL3msnvmb1hI4QwqaZdN230ADpDat2e4OllBo
j51Jm4dJ5bsiWeXEcsd0PPDPz7Jlzxmg8x733qKqMyGkeV2WOhGYZlPWbmGuaPeyyrjRazJfMBdC
59IK6qsnEDg5SIhmm27mys99577KJt+xxOEQjRzN0Csu0+A3Jn0PdwaFQ5jY/JdZCUjjJ4C8k+Dp
dH65aKRv7Di4U5h97UwlxywyGEeiIOURkmKS2OOsiimvvNMHTnSuVmY+/1mwa+iEuURfIN9vfbkl
FK0YH+vUXRLAVXc0vKWRc9jBgXC9ULsQcHPTDD/SSMnEkBJ1lr6JDMX1RgzyGImR+ybjxhlol1bi
d3hkU3PGEdefp42AZZxfhPOxuCFRE+J95GVvfkaB589rtZ1YQ4Nlcsphi15SAIYrDAhG4U2iq+C7
jqKZcLi+bl4Nyh21JBDIO857jE7wOmQ5YrQJMmXQFX2B07SCmIcrBlfiThww51TcsbjM/LvWEV9T
ENh3Kt4HnPlyZBQibcf+bSuvgAX/zH8/Gn4IBS2XJWe9zDPhO3jmYTmLfH/jWHsAr57Ns1pbsSyp
LU8+IWKYJ/hsuQc8uHg9++sFdjuNNr1aPuFXLu93lsNWeXYVgArmiier69cZ3u57nQntmspYrZen
sy24JOYzksVoUsgrOx/AxticVBIESksahn4hRz9sZx3G/9Qf/43qdJNdZ24+dZKrnlKabWXcm1HE
ZBjdnQM0YCr0PXrgmcpC+b4a/7/jjAlLLG6FOvXnQxQH0nptqiHpLxVb3RL1Vy69XRY+6P6vEyvk
ccQHdHUzZnZWwA7A7GDcmGwV4EPKNtGj7y/48uCzGB3kUMBnI27WUGD+6KGCMuzqZD9JofHWPydB
APcPTTxWjsx4+VfBcSvu9/Pv1+A9oHI1hwR+dmu5/hXTLd256nIWlDfZHkFT2B1X/4F65pzoGdjy
J2oEMoyDVyb2jNECPukvbvnZQaoioxXWZ1v+RTpQ+rbB5D7BgKBvS+sEjMhcgCMLfiAOTCxTz/dV
9TY93AYI7aDyAJeEmqZrlOvtpH3Zg1+pK7X7BJCcCogBq3lmuNNrdsWmfTRsAp8lGaViJqYX+Ht6
aByugHAC3++WfmLAz9Do5s43nGjXC5LQy8+nJwymBmA/tDPSLU8pthLgmMAi11bgSx9sLshO8/67
tVw2EkCtXySktZKzOSz5MLK5rzrLrN+sSH5wV70oU7/vyhl73IsaZbcmcjOQCx+0SSAru/YAEzdX
8/EJs+vMIz8kE5hdyddU4uk34iOGTysu8UDMhuRlnlQCxMcabGZ3oUEPtOlAsxw6weQiYpB6rHyw
0kbJaYc1sUaHc2H1dI/ypa/ioP6P1303JulYiu+b3/J06o7FPLO+uDVXFBAXOL1tBNhEIV2J5dOZ
xC0udW5eSWSWTfwHy7UxHmXaQnFRiOqPeNr9rNgPNVl6aAV0UwRKXP4uItKM53ath6gqnpYE2wXd
U+GA+NOuTQWenQiYTBRE7ivlBePVS+yLzq7FCpF1LY9OY6iQxcGCenEoWbtzwc29mIqwEE3DF1Tl
yNZahtQMyNdSoYlrMFTGK4/yrcc/xzeJOxAybJ8Zbe4UMPBraZdB40Lz+tlhzsh5HSHwy8q1K0dC
BJqGBpY8w2ECve5nhMXcLL2zHoGPmwyOXzIptSU1avoFzdNWXQyYvSdM3d8N1np/J2ycvdmOKVuV
PXoNFjoKA//M6cykL3MkNmc8plRnOpdZxpE1ZO94yI6pVOjw46XcdIXH96cHcLKxVOewh4Avwjc4
x0rc5RP0yU2uuSwt21x+pIn11ZYO+6mOmxOc7/y8Z1Sa3Mxkebw1I6V4DYMBNAJP8iaVt6OO59y7
2w5xcN3wN//YFFcnqySsePmlHpDkNxH3vOQrKBfAMV8P5eXr8tSxpw9CxYhNMBAjTBu5F9PjZzkV
FJqSxnuqE0p9okI0AO6BLR8/ST263dl7wckYpJP6Y++XF7ZQTumV4iCJE90s8xHzkNJrj44VuNpn
zXCH/mFK2zaR4+k6gn/BykjSDI9lTc75qu9YhriKgWHCLvLYhxjS4VI8yAY7OuAF4tdYRu5xhLp4
8IWdtrNWUSyFlqWjJVZALoExby/tEfq+fpwHAs6gHnlyvCTy0ARn8J+sGTEpFPr3OVhOjxL/Z39V
aorgq5GMl3Z03YKRLK7WDqfi/XmhuEsSYORSfwnpWkfzuE9/xxnSOiaHEyG7D/YW91KIxpEdOZxM
+PtF8a/Akk19IOz1bNVV7RfbDnwmv59VCfeQL0nXuscKkF5IPCbnF6CUg5bbDHMdni6yJZIrDfR1
YeHXkwVanuL65sXPSoAPGP8usR7/wu9jlfG8HnU8vs15qaWSvw+TyKqb995h/jLGm47xQDfSZPsK
MyfZr6dFesTTW2FEBKN8ke4DP50tYWNMd9ij4hmGlyM/uYG7YjgY7i6oEfuVD5xvdsKdbX1TirfI
xVpWCbun5LsdHQYzkYVNq+5B1oy/JtY7lKBhXCaeunIOAg2iohRQKAQLYnaS4PWZEBVl5NyQipoi
A1ltoNczE0jmQR2Em3oFzlOYrdNamLBCh2JpXRknJrWlzQjKgN559x45J/AcLW1x6i72Cf2sTevM
n1QR5unuASfBr8+tP7XnRwDMuxccei1AamqaQBS6RkOzhgTaU0XTaKMXGSOmSXgrEhpuXuT9L8gg
/Ia9H+pxOTMuTVO+i5xE5d9GnDVsIogAgxLvOfD1BgTA1BKV9ZETDOoWvfVYI9JutupPmQtatlx0
atDB/8b1099ogLTn3cPurwPNm4Y1yuTOcki3DuqvKkI6qipfOmqRzAyXe+HdBDUBGwsRbhxAYKtj
U+4+AVIaIc6J3nOKQEZh8KpFUAlTACFFfXbi4O1Ifwv5LWCMspwZEL9wKxvC8tjHDJ3ZPSZRH3vw
KhDbXksQoIqGo+melCbbUynyS3VR2a/yyCyodBFSAfayoNXlh975IcMHdxqH0QWTqc91YaFsb9bi
7AAlHO9iYTTX7tt4xdHopWWXZ2yHCGTDLiWaPG6YkWBYFFXTiE5ZPcR8IWNtyUiEvHLK5UaSQd/u
WcH8zJqbOVhY4jmTNimR5Svt1CIRlo9qEQmg73Giy6oitx59El027jbO1Iecre00b4mmRBVRYNgG
C7LuR+4HsXWTkhtanm8Ps/WhGeu5qPx94mkQJKFzJH3dWJTmLnZAP3z8lj+t9p7pASCfhHjiBNoe
XLWi8S3itIKIsHLYIEZXvN+jf60sm5uiSkdjamwFnzBN+RpjEmQTPa0GKJedt6JpRdmzvb1xS16R
MGbaPSaG3Cx8Ip5tKW7iCao2P/cE18x5SCmvqgdxwqXwZtWmeZnxWHAeDxCN3odJ6v5BsfsX3j7P
NQbFXwd8FD0p1DlptNvaeqrrC4I+frSvI9PviU6Q45I+6miyTNpL/jB8ccO5Q4U76T9Nv7o0enY5
knSREUbURF5h5VJKwE+XwP5yB5yb5LtC9LfWy9vfeo+J5WbwgomalUgTRM6h2OdMLQi713sRz1Nt
fIYqkIVpXyJQv0fmk+ICy8XjFFfjkWKCkiwFHfhFgUMzRBi6dqs3Ji4B2cw2UoO0BNtbwE3HVLqm
gE9qp/DGoT++TD154XP08VrXdpG+UF4YGcFZc+BljFPPwn0GiDAaxe/Mk5h+8HfXZ91/bNedmd3e
UqTw38i7fa/CS4KPTUDNQ9H1dgf4VoBNwiCmkrMz+rgPE+6ajxN0FCyR/wRzNXiY9WABks5eftL0
5522E5MCXWvMmOADkckFk3P11HFJdp5EGl3VAcOxQR1zfhh0hrPX4iektLctOuLvY/8X8sUUkB1Y
Ge0xGrRx0KWuUZaCdEDLadpIOgwH4STwqGybZbyNsUOVNQpxK+AbLrGZPPGOH9/YIlJ9UTGoTBDa
mRetN5+cz/iJME3O+k3Tt2C7rozr985v5mOiI06VkPIJUqcaKFuWN+OeapWOxHQX2R7LkL+6oBMO
ZdyDhAYTRjmsD59rS/Y4wxEBtZmqbiHyWzxCiRiAH/jLY9uIftdzz1QYIthVXkDhBTbKCEzazbhl
wW6xs6B/cNQ0kd9N9Mph9tPXamo6X6+qmgtCRc+7te1YtLgkNEF4j/z7igM9XwmB7U6nixoxUSDu
6ZN3pPkjg/jvQBeUrqnRxaNgg2u+/I6Nx//3w7cQfnp0axLC8IC9ZC31XeUNl1ht1YPM9s31V0XV
IYeUCqManx5jNTV9PLPkxqiYhhu9nSCnNQhBH982VXHZ63c6QBoqEUFapkTpV9ZBHmAFqSwwqgiB
Ezrk3T0wU08YLgl2SXklL7Hnl23NiWE/w/0ZtMj29JUMCgipDV0wQUGrGQJTAwAL2J0RbXwbqWPF
x0r3QQNsX4WdAnINg3hOuClyM3IU6FVFetajpA9beZimep8Zf2kxdw4HgMzxKXCz72VoNzLFHFuX
4weh/WuVjYresBaPBAqhzjOcewTvr2teovAoUyguFnp2nZlBzrS8qLoSRuLS9tmrXSHSTmucO9XE
nAKJN8eaIkUKDhYTW7X6Eq1tGR+VJd6YOC5G71O6/asJivvrfD2/bQclWTUQUSS78sNKxh6huTcs
skmnM425YEKrT9AL5mc9SkKsPlS0UN47qwOneq2PixlTM0Uv/6mtZJHwHrjefX2MNtUM4knkGR9e
TLTQedQblvoDLEteFy88l6PrhuRT6Nwui1q5teJ7avQUy44R/QI1idk/Wue9yu2PtVehs+HAb54c
1rc43OuZGdW8EfZpfXv08ibNH/LYLpRWpx9gQlHE5a1+B4RkEx0vABsaUBpjZmZbDDydE0AM9LT4
eL22UEFaETS3uTRllOSMy04uAYf7zFk6vFw6o198S9EI4O9d5k1+EBHmM4C5aBV1gXRtVi2w1SyF
slP8038JAmgLSXZiLp2RgvXz7Zqop+6UCc80veqc4ISeuFbydmcK0UMra1cxXn8fWfM3r0T8lSTV
a1tO4kkXwONaVH0/qUfYm91s0pRUWcwAwNChOX+FPqZ3tn0MyNbM7zqtbenKomsO+BPPIt8LM5YO
k8/41oJIzQMA0GGUO+C9VJw6F2VhE44Ks1Z4NUFPwT0EN+J1+Bgyi0JK2NUNM8W+T62dzRWe8HuB
euNjFzyVXAwQhGh2MwrWzAooqsElkpoCAymq3tEtuXaZp+bAPjvqYDrU4ZpG1isT8i8aeUkT/hN5
rD5Ym54PbyOZ+39o+xpgNT/MaGoL+Sfj0rMwjGG2AVG1q5ANdRFOI+rIEy/y7Xxyx+O5XA0lklj8
SRYYZVHBXXCGnNsd4p9PTBUamBBpgCixamgmmeLzO46sYLWzqgNbjkHRKrB97Z4MT4O7q/ZI0ySk
O7CcEbD+v6XJBL8771O2aL/NoQJoznMPuJJT+bV0uEcQMiTNo0aoZdVykP/fZPLbVcBxh5gpvj0v
ENq2qvz/Ozy5/tudlWMhVZKYJduZbC7oVXlBQ/IhzK3eoq7nZ34bYZqrkRnJ8hACoJn/A3tvwwOh
jdSCyO0RujA0ZMnaIxWEr98IhbWVVYM0ddxj0/OphKjdK7xQnPXmPugj7c+U8cSERoKb5jlF3pTS
sZetFF8Cg03zaa/8gWyKpYVY/igecqlpIzXtX3+GPdN+8xFd6ZBEkrf86Z3VVyUjXMkavy4gir7U
tmQUApFND0stW88XrGLYEkQKWE2iZBsbZ2PzR3T2xxSNhh0SsCZWDOFvqYAyZbJ4sTVyYzwS5+oP
+YQdqHT/rIta8zxyiQkWnNCecSJ7qLSUeIFSbI+v1aMEtTIISWl6WdUDvDLn2FzbIzBAyPi3R6ko
gs6ZBe9+B9tuifSM4NsU6HzFvqcW5ALmQg1okwEMVF3y4xLTtCYegxKG+CUBKM9YjLlAVMqLvhDW
QymHn7G8/+UanravY0yNJz+54tQHx5AzlMZQhIPaNgSBHrFeNznj92oK6bU0NxVHyW6gD7URsRJK
ImzlWid0u9uafegxn6IzNkcccOXKX1YnXZFV9NYcEF9yK2fSLJ9r5iryvAxcuFRut5ak8HKH8bLu
gS3j9lzmpS6FghAib8tBZFVEroUp0EBbwS3aMy9U7N0FagZfLts/YI9CeM65EYR1enrDSfYzc5o1
j4lWUdZ2WPQYJten7kIVpzlRCLlo2phwG/zlms6muomkWv2Xk/g87/gW537zP50pp0M44CAozwv+
e4CzSaL2ziixRKXml8Bevv5/fYkMYPptb9Orm6DA0OOiWhqSOhTaMdbRkmIqke8gG4fV9ELkLr2L
KvEccElK3hRdTQ4/9XZpRtx611/znjgwvFQaCG0dGxMBmosG6RhMWLE9S3Gb56ryW4rgeDUT41WG
kprrOESJpBk4+zlzvB+1LNgQdxO1wTZKiIvQaDpegBAv++7Tym2XSSgXyY3xeRSZWPThiwZtiowk
s2SgnCRLHJrGOJYAFZkIQSzIFgj6jNj0nw7bVZwwMYrpt3XykmIyJaNm4HDDDz/A0y8ctU4p3rgL
OpaoJQoTicdBXdxgkEQcPoA445KrEhuiFcJqOdrYO/szawWWAzHvfkKMeErYob8AI5fZ8UCE9Bau
vwimKsfgcOUMID6TY3oe+lDgxE1pIvSVv9CQ+QHJcSXcadS5waoVHvN+wMIGqN3sN3wMAdOKEOC9
uBHqil2bHSnyMBnpgP9uSnxu3H6ynW/o2HHFELyR0PPFtGUs1uuntb8mNOyvRQ+M9lnofNLWHN0C
dHnpiVRQcVW3fFiE76phmSZQSLWRlsjPhJOCYsxiHDAAzNpzb53siMPrOrieUcGPTHDHqlsHj/K6
AEqyGB1UYtMkWS0EUeEJ0HXf0jKaUb30GMNeZe9WN0l1o0oL4wAqTDe2wcAEAbKHd1aRsghCprZs
tj8o6bboTOWUCvy0jWthnOtB+4/weDDdmQ93cGtRIWobF66LPt19BgL4etRdR+Al3twJih5Gu/JG
Th0U8kgpG1UJOix5/WiykPK9CsaOqcPaKuHIoXJCGOQP7igSwFoK0Ad459L9mlUwnFRcM4S+SkMB
mC+foDGBopuMgWTnnYkClGJXcOYtipfNRfiKA0bpvYnb8nsW6VF20kMuiwTS3fEKWT1261DlTWdp
9t99S2/jeIfHZ6UCiFOvF3X8yvDddIe1u3e+MP0CJDVfYkjDmEPgDU2DyeZBXKHesfiUTOsP/kxm
ojzsF3AZLzSO+rx8u65M4bbd1XqDp5Xs0cKn/KoP9jxGmujiOJNh9NNcUryBsVUj9kl+zVmB9tmm
AoeFDkikb82f+Plgvh7MLJ3+UcLdSjuVTk355RGceeQ9pjpaJR4WVeFy2G4+kvFfCTTHkuV2khFr
6MRVMvE759Vj6xBu71w0Tn8cbEPeCMbdvpF2GNma44hB7PnhXHkiwq6bZ3wCQumnNbWjI0j/SFx6
mma2znlcAHVAGmDodtx8YjB6A2TZQMR4MDACllYuZj8vCDpiXn9jpMXSgtAe1ix1TgqU/2zOAH4F
My3YQBkgXBEpI+vWQNQStolQlFw37G1Mk3BTQ+xjH4y/Hf8ond9WQdNVVighIRCUCpAyjg0pJbgn
e31y2VdESyRY4K8PsvmcPi/R8EuxJcs4RfPaN8yw+6MuYg+pUcsHs8XQDWAWqfkZzE8TW5WZlLs7
QRFULaobqMYUoamoHRZgGmAuIX79erO8njppIJ4df0v/GUzRND95jNg4nxDdHTkC07hPe+T2ppoX
olpLHSVr+rNAYPqhfyet00Vo6O6bLRIStEJilbiA7oq7yop1jlzpHAanAJHiMp60QQ3I7M0KPWII
i8R0xaBLhYIBAI4RGm0Q1w2qdn39pYhf7KgglshBJ5A69z4Hr1zY2BhGbPGeTgjJfwxZtz8nIem8
N7pSV2NvsFYI3DcDYUOOr52Ptu6/fGAmP9miV8YeLnjTrGgO5lMpcgUOvFTwcacdQ4dZ+rexPwXU
dFLzkNFkyzG8VM/Z0G5jFQubTMVj1KHoLGfAxFpa9SPIy6kaBfWiHC0MQa9Hy+dMEx22jskDdY4v
Kepo9PmtvCNzsyTiZGbRcnpfSHGLk3bQ7L6ZhEIJISfhz44KzQgcaH1O9aKB+2EWBBzi7FGKKhU0
fnoTBaTf01+nWlShll4YzTOQC5urhvxLjnbjDpTxM7diPZAMcpyme2ozKLGX0GcVU5TXtVT+oCzd
TJMr6MKqyWUtWk2t8OQkAZGA+3t/7bUGW8NeUtm2dKhU0Unnhm9Vd/j7ZXVqVvc67cKDAriB3GRy
NDNfOCz0XijtSq9vGuWOWe0VINDhsAaXnD1V4q8RdUS5Yypzw2fRBkkCqmrokEUZ5U5ZBO0Dgn2o
Kb9N0LQ4L6eKwEfCLv88RyoVLXOiXwbGh9UtEBL4rIG5QMv0T3loXXoJcSrjU+laQ/h7DuGWW0aL
HVuuVGptAeG2tlJzly8mgnMXnZdlPEOBhE69MZz3+Q1tQum5XJrq7UfE3dCGOeo5KcXxwbFo87wt
OVzEIoWFr5TGNTHdnP9MLDB80uvn3ko6r5J+HDxj8UHntQAZ4Gbbsa/4zbbes+ywkqH7mXKxrlSQ
48rjdIcXcPeH5bn4QHyE7d+jhsrETR+cl/mGkhUl6R/I4Vho0dq6FTKqed9DK0On5BxUkqWZSz6y
+bXFpX1J1PS5uyP0LOIRTT28BXD+KFLwKyI8wdU7LCuD+x956vH84JdnSKqfsB4Qr5AcNDoRKQ+g
h/Kp0J/s0na9CWpJovreW8mBLkumWgw4zYsWBdUc6wuHJaHktK6yZeyl+CndSWjqiEXu61w8nYgD
K+T8zbxRYIQHSm6kQEEpwVwL9ukslnKbKHpLFOyosJUrz2IMF1WKpqGjzq+0Z27M9jj1RzNJWqjh
OddGkNwz7fvPtT3ayXVgFelGrHbEci8tjSeLxU396UPTdZxpU6xdeiHPsa2moP6YsMfXKrFTlcOp
eOZHvsL79rfivVO8YTg/XVqZFUDI4QurUbUPdEwxUyAkPWhbe3tp+FT6Jfx5237UW3Z3yEOqqN9e
3V5p7x+9jqCKUo1jEH7sMFBxU9iaB0MtEA9pFxblGpcUEpIkWJ3dKFcw5BJcNvke/UqmpYPLjz5k
OYfk74cTveS3nPx0t+PG1o9Yqze93G690uXaaYbeparv3ukcxbDynJrM8FizozHlaX2PJq0vBeVb
VzAwwWAlJsS5my/mSObohnc+d+8chzY3YIeog71dZseADTE3uTqv8B4jqkvjRJgrU0rG5yMR4fNK
95keP0oe2PEyOyTOKovY/sfGRuZJb+pcdAIZeF2AxGVQf8QqqZfP5I/olSlG8SPZlJaQig1uqNWm
4AOsdJFs9MZtGf5PEW7Rh29y/7gIXRPIsOf7m/qtF4SwPUBVEGNmWpti1qDsyOvyCWtjaLly1czY
HqxmeyO9HqPOi7hTBkLTZTvRDie3D7BUW7ijLPwRsFyVsVpSCACguuFblEsh8EJYs29WFn1qC5bP
SqELF6F28WpcxNF6/lcpsT0/oSZPiySl1nV7EF8JJTFkuGaY4q9tVmKGJSNIQo/LHP11WvjKdC5J
CfQ3/LZE6+MplaqUhXAIC4vLtprVVb+IFKfXk08DvKe4hBHjz+Nxm7p5HdtpCQc0c9OZz23Gc2t3
6I2AYV7AD+fKPPFi9F2G29Mz9eGKGAEeyzvpOQ0rHjcTTWTjTe2RvgHmyhr3N60c2lUzYxBy5RcA
h4qe5wK/tkeqrq6YEgPy3EAqcf27iTa02WJFSfSR6eaa0mDv2SjOmr6I8jogwqi4qsBBGgu8Myby
DSK3UXkH5dp1oYWYMqb1eoXVnOrFKLpIQdgrzsdhxr0lrDXDNuJrGNDtIDYV3cH4Jj8FtMXZ2zlE
7eDiAuExTmkcSIJS7pL/nHh3SnGVBf4ywwae0xnOpwb2nReRlVYeEhGZF6qTFXF+U+BK/95wPsc8
Iz0o05gvnhxYGYV4KZYJ/GtRyI82ki/sq1VUsk8TdzcpnEgA/LaJYiIP88cj4qtG7szG1TBFhm6d
SkYXwnTrqYKMrn04CJGmSPYxow8RQzjup1cA91mYapamVCZ2K3tzUFNpUxa/jl8jYnSehCET2iOJ
p08sG+IIBVPK1Sn7jvifEZ4DUiIUieYxRGIATCHj6N8ED6Qy5DzUZf1x4BEnmPbz7bkoABYT0nqj
NdeoV3p+7WN+h2rIyh8f0I8YTRwh76SJ6QVN8zRrwbJBD7vITE2tcwvOCmtxSutf9yhyyp4ms1Uf
aMcqGWYsS/jkZKXxetrv5nEaVEYLSXjf4HyhpFA31wucmjXNnqepRCdUI8R3tX6o9CBWTTQL1hhL
F707L5Jo6OnAxmZYk6N3A6VZRYXqUPt3zEW9r5Y4licQSrv5KXd+ptWKwuddIt0myyjYSKcpOVL8
yTcS/+QFx/UHwAvE5ELF7oMr41nm4paB9Xm0n9riLmLCmnLgFQySJPv4W2zC6DU/wneWyttyORGP
cQ2zKnG5Doxk7gsihGxP0iMnti977YWqV2MP3jHbHSjGBUAgdTilIPOR665RLCJokdVuntR/agCg
5BXZuwYvihPQO5p4H3wAiIjAbRnmyBbPLSh9nbM3X9ZcoxGFKG3+latOIeH/QXBuv8inKxnOp3Ho
QzZPp2bIA2qSZDNXhM7uT5BfWmUx2wyBgvZ6fu8rN9fF+RSnaIvnhyo+uIHWJJe6GmLx4cJiIgCV
fTn7nKgKveYLt4FVyhJBe834q2ueEJ1oyBgN1WFpOE3BajK6/IREoNQfaI2SD4slzIh1o0wor4C4
emyeIeai7fEU3oLz1xwZMcYo4rxixPwE8b7wfgH4U8E3XnBGrkiu8Bk1gOnmKkhNOp9/B5YTcEz1
SZA6hnfp3Nlj+DrR7D1dlyQwpA9D3c5w+yBnqpOX1CQNBml+28/gclW8wAry7TmrfRPBSGz2OhMi
GdW/8ZIuOhBurIUFZcvHsmZW8jpzFjfokD3jVhNOQ5vnAXENRuNItNoOGMTKEtREmGic0szn0wAB
RVsTNFd6bJIOdn7bbYsoLOtpaNue1DtVaz6qkAS1sc8SrhupElvRIiruKD7Q4BwxRE951P14g7uB
5mmCJv9R/kShsVcpLIixOPYMu1r6lZeryBlcQ6DUasnLHmonkiQkIPLFiLS/qDGPbX+VuljXE4f+
YO6RbRK7sUASFyMJeL3HsVldtNgR6UMRQzm3D4hPFExZaMQ1sjDe3sjrldMOvwzp5JeMu4H4BcAB
K+WLEIs8ioyeRWYnryAPzTEHhJ8Q+QVkzU/OUO4XFN6UocrC91Jlf3Oz0Y2o1JKdq+DXtH3KJBN9
ES2vQvIfuzCg45nIRxgNiWgD9yyaEeMH7XsyQeWmW07prnOW5SH+z3IJtPfrS4U+TBnasPELNGUI
7cIK1AcZb9X3L2M6Y7nXNzh5nKquXfsawKPjcBSA5zLoQ/9B2k9lMMdKNIpzik7bi9I2/g0AtZWK
cWVtqX3PGla9goMlG09uwFzQ9U6c0LRQKxy8x4GTSOiV6lkE/EKb8w0yvnYb0dF7WYmkYbEAFKU1
tMu/X+ktExrorJ30jZfreuKxkHO/86zp+Zc8gInxGqaEiVO+v99Bc7Ij4y/MLS5Dak0nV+sWra3+
/oG2v586sjrh4d7Md5OjMPvQqFnCy0pV32BZ7FZandlrMNSh6P/0P6oAjOyg2gprpXj4bWCa1oS8
WDaNo96HyYVmFd1fV9ErH155J+x1ldqrsO2jQUBPP5IwlqJcQBFxwlkm0ssF5vYWiJQxhkXWMjjY
0O0Ib7M6Tcs3Jaa+fnjO5bDQp/JYITnGnpUa7Zut/YyOuPnMr7rx3272ocJTJdVvzC6pnzNH9p3O
VWP0oWvdldt2eEk9foAD3YGEUp4/mD5Cq3Nz4CFL5n9nMN4elXtJc8aYEg5ZMtFAjHRXEQ9cyA63
gCzjRjEnA6CrbeH224v1oJbtZMarFS+LH47XkPVALQQdrQwxvhU23XxZnZXEhK42zMb+Y5lHF6ya
UVDduoGW66PfFQOBF0AWv7mkQIILW4A4lOLrtOuqwYrFPeqztEfKLUPPK47Y3xMFIB8l+eLjv7B9
HNPMWEpiOgP7SCTfZGQOKmoOdheLuYp8IYRmhc9B/fCz+pajE0a9aST0pH1CSPa1DcPsl+z3W8+T
Q32qi/ZKSjfobCWpIPykWr9NNRdbCDzwyE5j1UPTb5ZW3BuRZbEgpLJirNajn5O8Ma2USt7wKEen
iyOjtPZZWxrzT/eRTyPR2hvvjw5Fh6uCJjtlx+9WaWdOo1xyzfOqVSqm42Vpblp2nEiUfk3IRf9a
UQkaIdhEH6O4g0TDaXcEqROLNeVCGB6Lb31Q7IHmMt2loZy65NM+7lxBMd1sIz8g3xRXOL/UMLTE
DrY4WhPwD37b1i4s0BQCxvYy6YtiXXiSKmDzVNqvSxWeqXdRML9g6p25Q+YcpxHwtEgHoi2fQTy9
hdfDEavQSK9B1vAwXu4oN315XpNj2Guj5R3WvRc/oWgUUjqtHEK2hkDu2Ezdu9MEhCuQXjMxbyxe
/0JSI6nOLXa1viLdFZN8b4f8q188PbPblY9oAAApEFaDu/jg1lhLDqUrEtte/kyYz/81ferXzw43
KPRgSnhQvJLtZEWZDdURXbu2+06vxmQcC6FDHoAz8Fd9zjxn8UA6grWpunaj+frPi+1BLT/1wMxN
r8DJjgj6xlG/FU80zRssOY+nmUmtxyPgx7yxsQ0RqVr8SY77GrpGykT+3FsB22nxO3pRv4HhnU0F
R2OyPZMbvZcqg7x5vltUuVx01ovsxFsBr9EVhmk1kjv76WuaLhzFoi3Xbe4q2yAueKa1diJC81Wd
H8B0cf+r+sl839cRCBlFdIg/mhWP0yuKiv3QohCB5jOIk6B/Aj/3ywRY3iWJ/jc3KDF6Tv1qfnvu
J3/3Yrl5PfqGHdjpUtS0FjprAg3Shi85nS9H8YvQ9hACGS7WaEbFoDUxjY96JtlZZd3v0lwOkKV1
MBP/aKxTXQF7wai7TRW7pJm+gLFCOgErBh5YS5SiODcQqRErrqJmRUqY0Ntu0oMhVAWiug1k5KG/
+nDAcFH/y2r7uz2tQXbpLsk5RlQmojUqfPk0TSCyHLxg6p9Nkg3ZjbtzfbLaTJ0SFl/duh1QbOkO
lFfoeARw0AMdGDWPKnRzzoKNXPqCXNhDyVmIfNDkGYFl+5NZd1pntREHPygxmon6KCkBYEFKh5Nb
x1D8Gi+aj05J8q6H6Ou8bO3/Cq3XPM2ojv/XpRbGR/ZMOSM5IBjYWigAkJ8fwRasXkNi0MRzGkSK
mVhwbS1MR2QaHVesHByP07Hg6E6i4r75zwtGzcCqqbLhcJwcxXZWWYFk9JqDexXlpxObKa2Gb0RV
9iBib1GtlUmbs7WUIbiD+H5rEKY8njCkGedFdCPSTh2Q4/LsypTHcVeNQMG3FNFBvxiAAnjciocE
0bvVZEZTTs1MEPcbrJjHstWlU3PgD9J8NVUpcKZUwfXaOIR8XnHVbFKO1ejlpRYdlXwA8/k/kGNi
NZqYhit4/I76aOWfpKLAW65ncNTJwi8PQlXUubNiWnsIeE8dUHAr+U0jXEBdOLK9gF6Ov8ykYauQ
ROrYTBO3/KdRhso9zOPzZ6SGhHOxot3FTiijbAS5oP3SxLO8UKBxdOKwNXkPsO9Nc2t9q+bswsvw
QshNwFf9vBOgSs4kS/1XJfnty9wzgKygKc21SxnBY42EfbFWnQEXrDl7G69lZ1vECoImDzWFcRZb
lyPs626Ix3hWxOcUQMKha3YPdeWYe3yIvSVDhvM6sUsNVVGR+j9dLP1QfJCs6l5GTzB3D+GyxyU6
mXfbBw7IBJo1GKda8jL4biFH1lJl5maHVvo+0xofMEDqgj8x4i1JLSX+NnP7CNRKsOX2XaNNypVq
56WFmfGdhEXXiyHBPeEh5h7jdKVbtWT8y5+Bn+xB/xx6AH28Hg54e7pGTds9mku/UKn0cvVgbWzW
rtKKtEHh3vR0JexCUy7+ACs5PLE8JhlMsOVeKStN8KNMabxD18lCL4XOxglbSNPPQLtM8FxFmnmp
oG+5XXMWTRAr7hZtHA/EootcI7z5N9G+Y8jm9+KW8Q8AVpeHdo07WW5PU/x9q7/GkXBM4Xryn5Ig
pKPYkNuSGYr6RRK4YhaZ2LbgrP/h3IdHGrxPQymFonBP/dnoBBFB7UYT3tYP01+dnp4ygideZX+H
/5ioymoz6E5DzMjf0cGBFaAPBmb05NjffEkbq3pW/YmXZ5Ti9vU2bAe23I2X1yZV42DtKgQ/RsSE
M5RKP+ALzksKtYLApWtx1fXRg9VEOb/9VzJC11de/jiQwI8OjBhy9+z8ito4q8YjmUw0Nr5hJKsS
6BaPN0xhSwiTsMq2R8SuKQ/zkhv/BzD/cL9ahL/6IdbGgwLADLcUoJnyasm1dfeRK1tpIm8SvnEI
OkeHjTdGWSlMTEWJdcFzO1w+Ll6M7iqjyRYiuAx4u3CfJytCb+jF6oqnDhdK9EQ8/YOh7QxmhljJ
W6n6WRMJY3rmXMBl/EM/WYvDWtX59o+XeRCQ/NkKwsOw+5rDxZdGoqnZIq1hi3WsFOMxaF46p8dd
i+KAeoT889/2wUEBXMstT97Ko4J5WHsS6elLwnug1YP+aCzGzjga45vcGQ1hJB1Hx5CzH8eOMc9X
ttRqj/E3WqlnrMdK7EvzrGWXtC8ymGAm+V2whICwgtEgUdAyqht0t8MobKDsP8EQLXYrCjPr/L33
9K6vddTdfTYdz4IQgNmMwPNr4F/M4MFVwCRHrIIi/88E28DoGDD9Otf+5IaHPDKlefyhR8BozoLY
Z1ymMyCsyi1NX/bDYWGtNR3oO4NHYZVIWuG0JisrLOU4Ili5m6EshTPOwoBcVPKRvTcxejqLBv15
UAOSMa223HoZK7Zi8pzqPyzx3gLHYIiSk3SF7D2d05ZsCkT+0RYG7uIbVRDrdpLR+2P9u90Fmm7W
1ksMbC1qpB6ZGUjsTxrsHZVcqIdClQwnkO9ogyQWqG0crPkEuagj19dfWE91Pyzgije+1fBLx2n+
hV/36fxlONH8yy7kZIaxhmTs9WEtDimX10v1g0bk/cr0YhEV5e39wyZZw89xZsWwglQkyIrhBjMo
6iOIp9/FLJXoRTTfjyoErsF7fwFITTHxtDxlrUk/N43UK3GWXFT0cDqIe1zNWBrNZfPmFhaAZbLX
mR8TD7v6Eq0gVnH0Mcjbi1dsGBa9AI88wSxHm2AAXL3pXLSbM1X0z8XjsFwAIqzRd06lWPqRerLV
hh/gOzgOXJkn7jt2iUjh8aGUuYhM2XqQwF253Yj/je2hc3X7apue6Omm3ayETuitxsIGv0HrCpTq
hsOnCMT7LzombY7+yMRjzz7KpurakALJ+QvUSQgb87XUO5M5HTu3BllUwMNb4CBI6xC96Em+8Yw1
366bH3fBlArdoqWw6Z0+KW35edq5QlzNIKO/IAoY8FCTLEu8KaMxj5Oit6luDkcouP6NVBtCIpU6
D9oRqJBuqeckO3bXboxpcoIm3Ypqgd7rz/NNQNhSGS406bS2Z2Zk5OpORKcpbULGtuY07N8lhQ1x
3JEzZ5ecwYvMErXNAoylawGr0EirHcTaVGlrnmO8hI+tHn5A6sOXBYt/xKFkk0iRgbVa6R+Zv1MI
DO1P+Unw7eYKWDHv9q6bDe1OhC/+PeCHeoT7yHgj/Z0hAr83GmC4KPOJZQz1CO+kJ49hV4OuJco1
upJn3gOgR+B7fS/qL0HTf0/T4BYbqAhFfuSr9gkgggvZgHe7ku3cvXs1qZCgzdu9u2IB5du4/NgB
8oDyzAuitg02D9Myiu/z2rm0hCFEBpU46IXqvqmON9NrITYftKLIJukyuymMmcb4Me1XKeBkeizO
igmfVtpqm2SdTx8ZK2YR3dstKxR2nxWHMr+M9BmWJe3zuodAGuB3UMECdEq50epfgKCZ0HpNCbq/
Pt12Ph9uqRPifUoz1fA8M4vNVoEtz+GL9R0vNlikRlbTGr+UYyCHEgPL5POTVsx61cH+3VPfg9jR
QKuwCu/1dJqxw8ANAi60PyUQSRh2il1i5NdlqcBo+0/YXJ5x1Ls5TF3bn0pH1caRZ7OlbiWrj1Re
T6RpI0n0AAQSjwiiyVePej7OWPitploh3c4OF79BTo60qnFkqX2DM1vBtTELdoX+oRZgpCMsUcAq
oxX0F6AfOLOeCnjp/f8KB7UvNoHVhqj5RlB68pkf6lSkNoxHBUE02MH6cfjQ3fmgo4qwoITRwcqf
MqjJBq0O+rbFiNIvKIKTOu+v3WJDcCbzlnJzfgA7h1ZL5STiAEtBhgc7vmKdVXgk2IgXq+8w6CqM
/yeaLeE/kLQzyQZDcHA95mYhhHkl3WZXAIIItKt6Cl+BREv50q4T6MAMc83p0alwPpTva2GvzUFk
DzlWCt0vw53HmyRDK89l/3XRHQTozGWgOFoO71AUNyTwNsX2+IkG5pyh56mKrhPs1FJQcOO1uyiw
Nzc+vtxmdpoE6AcGtC1AZfeDeGQhlTDtXDxw0u90I9FVNGB3qBYLza/Lo89knENaBILPXsV9MueU
Pi4XYhJsFhcOUbIR7TdurWvZiR8YtRLyQXhR7+FCh23ic8W56nFmJKuSeR7UyKW/jUozo8txpnO3
r64r8XUseffHzPouQrsGwThWsD9IRO8M+T1+bAX7gWgGXuGwBLqRafyU0zHD64o+KeIiJ+EKpAZB
MQp6tnEDEBFZbiYSLxEeG/mbBNJhjPVw5hThd72+pxtotpjidAuN0tvhLEFwzHhY5tfIdR6biVHK
ZbZnEpKSuHoEi2k3GW8CJ3PlnYhcurhrOUOQEThs6jGxh13LXz175DvUu+sxwBy2TTAAAHM8+drt
TEy4hiZ8IOKXbexwGQrdCurfbrFaXn0+ScnLGLunt1gt7BdvB20G33CLtS8y5w4emg0iAZBI1Gd0
TWaetLscB1Xnk20R8a0kw9Yh/G59tXH/LBpqBnmtR3pa2o35luQXKQ5c5Fc4bgxlK8tmxrk/O9Jn
ttYCOxeA0ZnhBhdYrOm05y767DlivUivw31oxje4m0aIhi0ZzG4GBaZuAKYbqSVfEGOpR8uo8M5N
QOVisp2F958vi5ZrtR6k4mbyznCnXktbCRBv6b1Se0tejX9kIZfE1s1JeMNdjpcN1u0YsSwYWGBn
/VFKYpiVu4v8M6AWZlg4tD+Em/IOcBNRMbOL7pCsPv9htMqj27LIkZwPlRdsLiH4ufcOb0yzuiBO
flRCiYTQ/BPJNMF96b/rWOtnJRNTSBGdfzcs5zsknJAznQU79WAii4Aultott/mdM7DPvc/YhGmA
bEKc2LcwV/wH3xSpUPmLI6j7Dju4jRFyTb2eVfLmHdPdKZVzPgYtzkEqiUXYIs+MMzfb/AmxqwMc
zqQAjiqRGLQBB/LZNA314Vr2rvm//p+64dvGH2qp3J+1kQ6ZlD8kcyWJAt8Xqxp+GMPzOOZNCWtK
s9zwuKOhycT9Y98s5raXGDLgcnTzvRvGwKg3iW3wlPt4IR8jN/rGz36bpb83/PCY02o3JNePuIAW
SshTCUfUOQZ6ZwgbqGBmY8gIewGFNhen3rpUlx+l0eVgLG0YeOvcVQueLQt74i+IziP2Enh2QLoJ
Rc5zlzlevKaQEP3d16PE9OfyZZlBIFqatNcgD0mkF5aTOh/Us67TjwvW+VfQYgYSW10vzYjsaSF/
QBwjOcY3IAZPGrgHdP3cSzbSntf8D4CREy1ulPvmTL/RGvmwfZflBsWnfv6MkiWsa3dQ8HJ0GTjj
5izihJmdmclBPvZ46l9Zx9FlzOajOrTUSnCLSScJyJoqTTqh9FmjF9SeVZ+FKuuSYaeeHPkzTc53
2rkrR7XiCu27jodKX+NlOakEeYejtvkmLDWyNtny2EV4fE+mXXyT4vXUGcRDYRwF6E5+CG3bpX90
QwhbMBZtdoaMsJEj41xi2iVi3dMTquG0Kn0kueWNkPXU1seUdHCRkWdjT++h3Vxv7zjntvSF1JGF
ooFJKMuEieqojS2lN5SR8cVfyLth665DJC7uRyrqAuAW+OznnbiIckH6TatH2OmOeGCq6k7S1+iD
FsJfgV/vSGJDYiPfulJgkFGLVquHTUhvpHcynkPLdyftMxcUgpK8vhO/ooGC69ZOkNh+F97yFUIa
Y/irYGBnbhjAws1pqORGCxDvz+8yA7I8vQBrGmcUzb4bNQ7+gkWLInVNY2/Edbni6Z6oiiLbdzDc
DH8ikG+NHmaxe4FDYNimozsjiUBI182Fm+KSoAXhVj+xZph8919BG3pA/+zlQs6J/NfR2HUslbYy
eUcBtoHE1Vx6+4g5r1JRz6XDntmO+mn/BfcCm0c2qgFIT6SSUGrvpbtK6g8FW3a0Q0t3fOfvrAmR
MjH5pJ1PAs+3yeFTta8/Yk20nSZWFNVZTE/LP+rGEXGu8yswmLw1vHzmhvrpnusGtmvu5YfvA/qV
41G4endXhNvOZldTqC9xTf32HYt4LGXWf8TQrf/OBNCJKzn8PWU1XxAezIkTTUBMXWPn5eNgNS/F
WrSnSoVJgNjwS6cWNokm4GLX6zK9hKzGP0UCn5oT3DhhIskKQEVSyJ9dfhYgVtDfkvmMf08hsS3Y
8v9YEf284H6eYoTPQCoxumnIQ4lODtMvsm/TtE7d22hP0bVSq1fgL+bQ2DyXc0CKPj0/6q7ordHP
F7aY8o8An2VOSRITO3vPyjPt7nK5PlI0tOaLn0mJYgHrUF4WK9bjcwhLDgO9VdA2fUzMha67keQU
owzWCF2FYLUWUXmLOd4bqHG2xqR2xeB6rNcKeQ5JGDb/O1ZTO4X/D2oJxOhGhssnnECmvCym1j2W
moqZJ7lHK7JVe4npCONQ8cS7LDv+f0pTSOvdFs13glvtVDuMw9lA/LqTQ4R5jYlYFYMcCLXpIHVz
xfIvwJIg70tiKAKyG6DD/snPWREnL/YlIe5lMAQPPYKtrXsn36PQFwzZ2qJVasLMp806urmylzAU
KRGO3LhYSdKR1KSnbVt89sGRP65rADOUpjQI3JAnlterxKO7QkDPFGaBufGQNlFu+KVBplpmYvv+
BGivb0T51VaHy17HcEKZoTYDhk1pUdsJli9sT+lBJ9PAgVd3pOUpdRvxhMaP0r9u+CXFn0wX6xtQ
SQ2Ev+F+4nHSHyycGXUW2lz4pT6RTIqr0TbmzvkkccTtTOzti4B6hqQsRrsmcdal+iCZMsiG22e/
Ca2f1FUdZXGqbdBNVb02O4QWjzx/A8CQ8bOsm2S6svnHgQ5EMwVTlvu5h+H9Gq5KhDPTUJxH7qGK
zOsH2Gk3F/5RpatubMohkJPXpH4a6wvlIOxy2iu4BbZx79UUcCLtv/lJs2SgluuBQYNknQd3F01h
zRSYmur9xnqZNdnZimS6nx28xhXBDwTOK/5en+A+jmWRfnr2N/IcXr8RMgPEjUTVQC7HulfLpbDr
OWGOnv7Re2oC/lkAUtBI3SQLbTViWR1+ctsl93TNZkAo9VUNbFYGOtCWQvKNapXmWjMSgWH5d6zN
AFBwLV5cWIpgILjC516OxSDxYSez960bZESzsAZscig05WVlq/d5qx2IVjBFWZgbzPwBIdn2XPEs
jJ/S3gdk8UXUcIque6vekHzQT83hh+Q93Kxs0+G8gHWp45IcAENlBzj+KFoXwb8MK+3/wCBjletS
plMadMhW0akcPYMFj9etjXe/9TMPQfVNNdd+DYRiHQJJySBLGUlFcjSXBGkCVK34r/1rzIc76Opk
u0OYyNkDo06+0S/bWAZ8nYuz4RbNEKFsyum357Tp8H5AYxiRLh//YTYKBvHwglXGpt+h7vdIeALq
pgL9C+A/rZPLu6VVLYzObuP6zNY9MTYpqUl+Xm3gOny00+XJZcIKpbpy8nAUpgO+BQgbV3RD3s1u
u9m4OGn5qjlUAbC8Ipbe/o2RPZYq6X1ZVSvPWvYTiy60qF5i1WcbVg+wzc+uFp8hiPwH7Iq5ULij
N6DR4Hwg4xrz6E2TWcuEVuEUdhVKwDOWR7fxxSVjoPNq6qxCFfPHJ3RnAlIczZ7tZYXJWa5VBOeR
0AyQcIx+vRlTLtgQ8PXTO0CgzeYCtE/id51nlnF2/wKmnRQQ9qqm9Rvt76CiRCrIWpEUnydL+jno
XWAYMrai/8WvJuE/hcs0R97Lo2OoiGMmKUY+jsGxJmAAd5xjqsjrXp0eAyz80zz4o4MtLmXBKjcR
Hqg87H2WCIqGvqMc2aLcJvNSObrpB54KOj67dwr9SxiSkeTu7JbU9q3eFIsfq5nY+DZb+QLO+dKz
42A2cvSCM8ShJ11r/WulGkLxItsefwzYKj/kCeX2k2lZMeQM7OEh6U1Nu726hCu8U1H+pjGLDxQ2
6G8DynzuAUgadOp6FxjM94vYnPK2601xOrs8Y/9C+KS2/XzVBAKyhB4PHwKN7k5FAVtFJzFFPa7e
ODAMkj/ZDEDUQrzhasVcdV+l+R4i1+XjUOqQXiAYjjx2gINLggT6zfs6sZdiWOUpsUySUviFgziK
BVSdx2IAw+8s4YtcyKvSizL14PLK/hRPTaufJsw5wXPpBvQtv+2OBNLxyF5tFnEvi9KLFwAXIUsS
xUzOd6ekL5N/9xJ15Euut3M22tJAZ8TcC7PshNGiFWaYUtKvWiCpr51b8bSgCLnaYd9BmhWVgOLE
G2J85nGSpSN3IkzNIzx7liAW4IMkfVIlSh7+p5/LB2XEcJfzhD6MhHTXpJTBdAHRwZODy5PTLWeZ
DrXgJlkRKC06TImG6m6tKFEP2v3uxsXj9WnN7de9xxy8N71aCAMHk68M+oprypogaGirbs6NwmpB
yn+49CcS9djhkVCQ5RVUTIwMMfU9xIM5M5G2pgy4TRDukopBtyFwttU8Ka+zi8kGW8ehJkDlYcXQ
YZAigpkEKiwQ9/KSoADAaCMhUr3JEBuzcIfyy/Y4GwztXuLx2ZoYDNVHGrSyWlPXuortIxhasjhp
8RyT4jdRYm0jmZuuLJKICoy3kY9KpeAoKlpyHQDiSyjn57tYVMp4juYAzTEC0lP2UIlY24K52YwD
gnl5/Kvy5QKIuCZM3U4dI9POSrJeF7ax8rwj4KJj2oKhfQ5UPQxtTgYLOM2Lt8n+v0SySTYJiPS5
BzjW3ibR7Bnlnm7giPxrRFzn5W4RrlU0m7ec+oIJToyV2EnZa2NA8WTVQbjuw98bEX76T3OENtCI
4awazdqursaJLAThQ2dbjxRm8aThONH0LvH4vg3Wq3mosNNHez/5uAwnGRc1ghSD0O132jzynUYX
aTM+2ut2izVoqi+4lr88G/XBlbsjUsK0eADfsxyDk/srIhSFK8KvgUiJ+u7j7bHBT6zosIH5GfOd
tk1g0BR2R4Jj2u8V6sKxP8k77+7lWI+1nU1G+Zr6fTUDPxx3DAUrWKXheyVjFXcFqHR6m52m2JYn
c5hbi3o1eGhTadai1n0yVyLZhYS7nvag2+BASWexYTyGG9mRfT37AxI51Zc6prg14Yg+HAhMZxXj
9BA58jvz74NQJSqZUW8IGa/xePPCd8fAbnaKSS1wJjd3RiAI1WZsovBNRxr+qYMRie7owLN16SFw
NolmAXMeL1K+C0x50s12YBjZ9Fpfqowt44XB7+MpGYqJeKGcDtLCvw7XPW6b3c43SdNk54xUECMG
d7GXdl7hDLsXchZVkhctjuhCRikLXnx0yBUu5RbkIavHmUYNk60Du3VhMMeBjUAyBJ17YWJqVw37
Qqifcx2JjkXnsHfwZROAFu9qd3Wz4p8NNbJLJD98a7K/Fv6uUsDm5guibnOWk/PGtMjxLjQ0FRsU
f88Hq9bnmHb2PAFEKob0DexLnfX9UPEJRge/lKqI7uP72pWFvh6PaKdCOznfGVQZ5R+z59DXJx0A
en56M7sVhmHd67G09FoUjHdRTF/tBJviNmd79Oh0/DGAc96FLh+v1mjJJM+hFEwk7st31L1Gjgg0
qeKZj9YXPesHHkyuv6v0uTJORnEVtu4BRVVivXifAwgV+FheQwI0KUhXnTcMZCrG7ZPjsj2YVtO7
44rtI6zshOtxnkiArDvEe9L/1Sz+zb0Sy81g1L94ptV8B7fyRlWb7RmxoRDth+rStbZ5WXbt/E9+
7j+8TplSE2MJ9o4HgoFrFop/vq4G8bWib3l/XuwPnGJ7Bp2peD/FExKztfDhutPYe3kzBdNfqRI7
QZXiQbDj0i1VwJzZNzvky4M1ZVtG9+FEWj8Ned601DBbsT3f1O4Mt1jci22nRws/Rq0peqOEPm/x
0uuIZ/6VRQ3dqkgls4FtqChsz5Wm6LC9FUbpzuRQiOy30/sU4oQS2iQlBLB4euZuUm7READnJbSH
W50dZQ3ALNxbVhbY+z0XJYHNWO5/EPL29mJIihoJwsUrUL64bWeP8BUv573PCeDZiloKFYJD1awE
iBXCO2QciIVvoNX72AYRoZOQY7SHOwRoAzuBu5rnoy8MCN5IuRcsLlF2qcJU3pX/PcnOtaSwyvy3
pfgU10iEQq6DhxS/Wd/Sh8Rc1pTCd/m+eY7yp3ftskh0r4cer48s0lz3SILsodBYxE66fnkp33dB
lZ+a0ajUB4zX1L5/V2VSg9zCGWf8MjbA4P7Q2rY5kU1WHYvwUAmxKo1xYUhgiOXIs9Uy9HD59a/i
R3Lv9WpZjlDNNYvltH7S+NPD63BrPxgxLwvsb+cSKz7gDpPF9emiOLEfLis/82AXgJXHSCIsQ/Fh
vsnJ4P96u2Z05OuFhDz60nHZMFWghmWbsLKpjQ5K7IclaaV64/TIIekaYZYHMDW0yBw82KpoZXMi
1Bk/0+UVDtR6KGMTlZkSNrtH/pkR6lvMtdZQhJ2V7eyDI+KdCJgzKEwn/J8TSHVvi3Q1x68RMqUF
XIuIu5WnZ3O52gPfjOqtZlsLFjJuWzKdLGnsCSoff4Z9U7ti5HKpsjU/Ls1o11pGD+U+KU9kLWfN
eUx7uYMx+WO1us5K3+VKnW5Nq6YIQct+RKX2lVj2/MUOiSAxkz83UWLIbC/YXh/CdLnkBPsk1oMH
mc4HrS+x6+oU3IBYDiYds1473RBBoNG4Fwk2Mu1m15zxeKwroxWZinnWWWc9p55jW6wGeRqskSx9
pwA3MB+B4RyvvCqgxkbM2vUP+sEHh9epzcZolXk69DlUPnQNGAqm0wBZOIP26NmaqhsJPbQmqZD4
vE+MmccL2hGwDOMlbspeJyfjI9CGtDoRB5vRZ+MiQdjKltkqCyzIqJUKCcRXBWyqQvANuRnszkKm
i3PLxMPIYH+wGnTqPH/ox52bevqjfn9WlAmCY8X9RC6lj1ZfP9ss23f37COtlewm8c5yhWXPrWGX
rVShe5Ga9st1e/2aPrLl2VR0GuSkpX4CHWZhH02okWXMGtpfCgnrMpqXUriPQbSiUiILm/elZxVQ
GmK5RZkMCaers6G8KmeSLJKvDw3lSFGT8xjRovtkd5f/0qMTkndO+dyokBZOiLfz/TPuBkqjxM8A
Lfdux3gbm0xQideT+Tvx9nW7DecX8tP8DlvjpIRwbbWFzn0e7kw/ZbkO/qHPxzevox69lL0oOHAx
Xc19XaoUVtGDVKXlXIF5TiAWiOqeyHE1347tmfm6M3u9ZFvxcVv3Qk7bf7Y2zaHEgAy2fnq2gwnr
ZGwOaMZibHSrsDkzNwnQZCtABqVHZLdBlvYf81Zfr+Wp0DJpX9oOJQj6oGzogtfEqXErEU81phcT
mTZnO6+XDzFPzJG2rxFlqlhkHLtfWWb3zJpDutAzsT+ePvbli6h+8yaOkw+xLycqgvISNgTN2uzx
06uOkjpGJtUM34RGFountqEsjK5nX/Syp8sOsd4/g+UZcP2r9dQiP7VBXLZ3lZOFujqtHFGsPb8R
PaOv8omWIuP6Zjrqkx7fMqvWKha5cSnWhHbBnpJ5qzFjnPcbw4bPTZ26rv9EsCimH3+R7jw9YqTh
k2pzn/nisVmjLol97kCQTr4LaDYtIRWOnl1Lb6pS6KkBxw/SNYMmMuxIsqB/+eHluYAek4XUqZoY
DLu26MjjQmalq5VnG8BMGTz97AqtogbB+hQs7Ds0RXYwwE8crYrd25erXHd4pKM1nuopwvp0zCUc
XTAyw7Vus4qW8HNNvisyzijCxBTPOdIntQGuGMZUmmvuxSdXJjWtTJcR3gmbL93Aprih7LngwX/v
uDSkmocjr5YJ2g0lwjf6EmRa2Qa7IeLkw/Q5nmVgMIbEpG9q/E5VjFqY460t/pwmVTy1qtYmvbh4
3Rq7ZBrEBGAtRpz/c0azRywpCz+Bo+YkqjZoYkGZHGlzVxuTRFu/pvwTbeYeVB1hojcEPJTJS1Fg
RPIIZjTBDDr4ZhslAGgwPRXPJE5dvNrBJDRg43nwmlDT6uh2E6iMG6Ym8a3RV3N4zcrBreUIZsI1
y7Fr4zRBZtuDIjqvANZ0poQj6ENveeIQ1RFAMhtvBmTAHHMGAbmky4XWXHpzvw3kXTNlcmVjKD0I
uejHBaiX4nqjaFENs+7tP//rSEvyMiJ+0cz2G4JB0N/nFNdOioEAboN6WuhZu+r/qu2CdSIcxS1J
XWneZxgKS56lpvTAhSOvym525uoiNVgstPIFXPv1MqitG4ffMcQkpeFgb0r9vu8Ls2TqOYzHH4+8
T8vEiSS+On8N+LrHUSdjOY7xf3a0PcToD1XMDGBM252sfSSqP36fM3TMYXAKemu5gpISH8u7XrwA
+ods/yVmNzVK6gUy78bxgI0eL/njNUzHLdQQFQ4xUHdBiWWrfU9oAT7nK7GET9QDOyOsLJ/Bu7NJ
oOc5b2qcvKHuI/Q3Ds577NdDcj4qIrmY56AmuBGooqQb29ZN4i7FPDKyeQ9CCEiYPaEpeb6Ebuh/
uNhVAeELGue6Fgbkv46bkMvZWrCySl4RJWIiWH8xFRKq3GUBCYuGGksC/PvmV5Oa83KlDJN1tzYB
ESW1BCRJ+215EvZlgQGNqxtbOqN2q7HF6Ti82fqVg+c/RBMH/aT7S5GT+EUVTDJYYPl3A7j/5+iG
G0/HC0BgDn7gH2Cv9PKLYRrxas8/VjZGMOQSLrXwCnDefR84H+R6MCmmeInP6gxNgFfBj9HKRVcS
SlZ1DCLIjThbNrVn2eiGdB+rD5grlSQUP6+7QfQ+Bvycajqsw36byIttmb/daSsSs7Z0J2Lr0WW/
v7iv96X1bbeAlY7ziMmFpK5NKeG7Bru1iqOsNOxjvrzl7YQs1xxKMExOPHmxnFinlGecKpY+fwCF
1+Q2AMVBeiY9igjoZoq9wxdE3g6EXZsXR+TObqyHNkbB9iAT9CGHkqGFKOLQEu9DxpybAOvNkC25
3afac3gaACiyVWGw40BgFxVi21196wSNh10YZsBfHcmmWkg/PAGEUwywmzknwshNXefffeqR7ZF3
HusM5Hd39NKoRcIQvorxBlsk9cF168XSOIIx0XcC7rL2Tll5LQj2vAmIJKQpNDCtrQxJhtLcdbsz
WrcZhBMsh+YK6UgGejHW5GH9KtV3uXrHMCYD433DBKo61J1121cE9RvHTejvYUzpMzm3cnuSM0C9
P2nA50hm5iFtcX/NBm7ZzR87fxVGwqcqKhtO5W0UXy5XBsvao8yGRPjTlDWy7oEC7yg10eudN+aP
PBvT68MBvvOCd7MkQnQ4cJnkquc5PojTut/U4nZdCfJ6zUolheYUC4awuFVas6oKrfRjXXBuckY4
L+YtoX0n8uLEs+3R5JBVzF4AmDfgXs4u3BGrMYrcjxJmbXXcFKAGLAemEZYu+auUlJT0dnIxFmzR
AKlFvpHgN0SHwc6No/mQFqp4Al493QABckYyoGwstM0fKFOaawffKZGfk2OAqC/7yt2frqeuTdfK
xbm29vTrC1AJE/4F/PvH8iqRaaF+CVdV7+LG81n9gRL8A7UXsL1ECssK88YLhhoIfFP4sEVT95l7
UTvhVgIbeHqS6256e3+Y3Mayh8r8tt2tEowCrNiacPQFY/Qc8VwyxcOahGUvx4JmlpvH8qheA+vQ
LmL4SLb/xVbVXGhoOWz+wL1gImxZln079lmHAOYEi/j67WOsjNPYMbK4CMnS6J96PGLFiHA0ypwa
vmMhQcrK2DMaJgJac2+wzXPvCMBsN2YHxjCnrw930KIVif/4lxt1uq3DF4mdrRLlLwuDoCAUP623
kgDQ3o7YrlZCXWiJxsCVkfRFwq1A3VtcAxGYAkhxDAUhviVecJ0JVX4nacqiVrX3pboXZxkSFWD+
MiLBNbyQlFz1YlPAkVmiJDQ6e/7RVj50gkuJZL6V8YNZ/Yk6UBR/MFFEht5EbhNWoPJZQrkJdXV2
4coqQ8ABVOcXB/eCt/h+a4eFq5jUo1rlX+y3vcP/G/Km1J4siiavbEk9XGiAy6PbcT5+BDsuR9TJ
YUEqmuO/xffRCayDKRdqgWRHBYO5b2eW4GePBQDDpRpoRyv/I7OMkPiCgcVzH01SLcSckv7WXVpW
1UnbZS5wMDLd9u6YoraF5pUO6cHIOkUxg+9rdeMlDLmAgfPOeAl8zHmy4ns1xv00Dphz3PR3swGc
YnOB5+lDPu+BIKmnB77l+ffnFkejqVkCTNdBXVEHYtfjsld5v9q0vZVr7fAQRsdD7TMF2iymcCnM
rztSCdfcl3WGh87YKBfpZqkbuqiuF1RFg+dEij80wjyt9WU/wd/aUfvLxkatsXDi0T1mcFgjB+Nv
mJfDBtfchJZhMe/XiQJdVI9nyz+WeG5p6jPfdQ49kE8+04UBCjXqpU/S++JRzA6vyQwFZWNsYjXm
wEHkD4CFPXFIa1RcAqVp2u1lGjJOd3UjHMXTASgatZpwCY2CoQiv0e21RN4ppHu4xgJumWeUBGDd
jZDSD8Yi12QicCVP13s1NIr1QiRwUk0r+IEctEoooEz7x4H1H6sngIXGMQNFoWDZ3NshZqggEQqK
X9LgrZJEIw5/xeIkKMuj3c+kDCdOFhPOb/5tI8DqI1NiS449CRRnjCN1QLwOCKJEmaf58Fu1oByn
yoPdyJh6Dk36VcyY6hgT5sDjco6Rumrjn5jq7U94x+wnwsIYxCp/Pr0wl5GGABd/5hTEfvt3cMdS
h8/Gm6RPaZpfpKz8woRxzDtggBVL2OT31weQBzrPhKiAiOd4v3GYsaqWOWLhxNhzt99EfDj32d46
ThN6m/ESu27iGiqB9eZPIV6pp5k8h7/FyhAkAFANOnq4m17aOucxeQBHbmS97Of4eNf5HLosdEG2
ReSRWzI5ryO0ZqLICDmnZOWD2xbUsLkmrJakMgY02dLCI4/JVjtu/ZfFo0oW1KMULDPEyiZQo2KV
aj1jtlxwboJ+2tlSWeX/TcipVSj4xiSgmEJbgcqF3o6Bv07NVni4uXdjTaz1beX0okvmdtpjK0e2
nQwl9CcggpiVrxlrpVj8qCnd3ytSOsTFgwMgMp2Gv2VP+sdOJF7SLuv5sCALl/o+VKo8LATp49Lm
eeDW01+BiFDQp+zXCVsoYiQ9O4LvCY/Esmr3IWFmetl9mDfygVUmqD2E5zQKAmxf7v1+29SxWyQA
59eD+piqus7J24oWPaB9rFmQqzp9DHfmXOPsXbOKZyt5VUx2dY1fQvTeIjzgYnohUGf+BRuuqfiO
DfM3iGQlgAHwQkuNPIU1POFmf7GEhumWIArzqNwqkD5U219Xe6Pei8s8zPQzJ5eowXEuVzIliZZ/
RzNUpyOI1mDf857DQup2wWx2VW85wbnVzucKwZafCyP19zwC0QBiLn4Wbkn+d/h9PYAC4Faw08tW
mkpac5oFZYUPMsW2USESG6ts+Ij3zxoKeEtLGb03SG34XWzVtrQiQtDMK4hed3jho64ruBS1E2Ou
IouY2qthFCcFy/sGY+g2kXKs1flGUBv+CO7P+h03udVeJdYT1DOidSYaLCnjC6ZBO7FD1s+ORadr
65EM/7Neoiaem4P5Y99HnI9NADBcqZzXiIB/2bsz0datGdZzNSBtoP2wE0civYL72PuwJfuryR6x
nQAFamMhWS/P8CNzAAFbXT6F4q9TR67oIt27/lUCTNXUk67nhEBrFK6FMj/JeLgYDlyOmOeoPRLv
Hp29AO9DEpkGY5XzBdq2fa2/0QwrT83xskcrDMWX3BNISLXzKY39KlhcThQMDeajn6QHYHrlTGka
33ri5eP6pvLnkPE6+7yed9UL3JSt3eLotLrcQ4Epz6oIEM2YdJ/vYnvgeY/6WhhSLAXNRG62kmg6
Ebx9BbkFXYslRHACwhHfdWX7UQHPS0YXAwNbswkdQdwmAuHPSQkHLAmkdx0K6Xb88EnZLPHuVMWm
mw/qmNDRDxxnXo6RygPmTXhSrIaSud5t3NkasdTjP7SyOpNGlVdSm2IU1WfQawlzT3OVY2Jq2sQc
HPXCLmlpNnOrDLc3YL4joIyFz5aMz67hU6PZVD1hCcHlbzGgaDKOQwDuHe6qvZsDNtxoWtNSIXx5
ZK1fH1KU5XQ3tqgnf3/sbClwIZNtAPUQIxF6/hN3DCrCG0cn5aUzweXURrXcP+hXoIoW5QrE2N+M
Hu0ULQxHaqEloNux7QxSFUiHm2hDd0/HJzhhjNwdnLlwprb/GD9agyCo4xdfnSNkulYK1p1pQ8e8
Mpxl8AJOH+2rIuQLbsG0Bw13EDaIVFQKObYunLjukjrpTKAtqfp3k9JbOdFWOGCwylvMQBb0ZzgQ
ZcJ6bWwPjlayc2iIOa1ACNrGqecEm5w+gK1RyRvqr59hOVH/DBhRBjUP7uOc1C/7sNX5pJIqxd46
/bieeBJ0UDW6MGAAgB6K6jUPTNSOb6ZlxDeSZxs0F2KYXaeZ3JPNcUukwZJ5nf3o2U/n4VWmj1jN
PykIUnprrXliw++vY96JCBTosK7krkcDRXl5/zKoZlXzEVz5G0g/bW19nt2qcNkN2ODzAQTQjG5x
rg0PLAy2XVnSI+6yS6uOKYGJcsNQzIMjy2tF4uWdYk4EuwbKs+lqIXmPhgpXupW1cQK6lzMTPaF1
+f8tBz89fvwh3heRfuLRVx/bkC+S1vKW+26F6sV1E6i8iOygFke7SJYq/hfM5B9YQy4d9uKma5jW
BBkyV7p2cJxMP+LdO50j2d4sKHjJUzzGJOlxa6gfhShNc9Z9f9ZQQr3n5YC1RMQckgFbQyYhn+o0
lKZrKeAEb5JkZeQT6Z6uQNt6ZlPjUE7Esqac9B34KwLRZUldHcCZMp6YrObM3EPYsZUazVVkzeYd
ml77mK3tzyMM1R+r0FVONJZlrImng7Y4pn+Z3Ho0skUfyZlJ4Xj3ldXwQoL+rGbOH9wvDrfcoXXj
A50zSIXzxxas6eDVF9RZAWvagcNLu4ro5Ix5doAdxXfWCD1EHo4vZshB3WF66hT2rJqNHdFJA7rK
L7g1TI+zEucFVcQFcD94/W6F8lfw6yXVKiVE5LR/14qf83I9p6pOgJ6tOCdbMgMExjF29esrIBWW
kb4Wk7Z5bD1tmUHC0VD/yDj65M1JBNdVfZj8e2FWFtuDxqHof/DORMNZBVGECnvCm/PRxVzS1qvH
xgMrICUAuT76uIdfHtCx0z7XGP7LEIU0aeLZ6q1/usep+P+z8TjezrkGcHm2q8wlNdjexcuUcZBv
ouRCJHXXDBcitLKs+oio6TU0Htofoz+qmiPR8qguvnVU7XfWj+AvAffVXVzs44DIoTFk1Bd29we+
JO1VnPTARrI2d92gqutq4izeb0f8CCpxqDHK8Ug42nsI0xXsJMYJFgU5lUj8vLJzWQverrWd2pZ6
kU6a0CmqZ4ggzVGHYvWgJipPbnCm7pEo+Tjb9iyCg+5U2tSF3PtPrlX0YUlat5Ss2TTUsacvRrzA
6gn+LdqlMYzO5w6rquQLTEI5qIRRlfkEE1lKXqENC8w1tR1lN3UDiE76aKWJ40ep8TzucWeyDgW7
eFdnM+8uezvdoE+RTJx3knNK3kABSGvUOU/x+SgAwjq64lE4fNJE0Ul1k+EE9f6JbkRG+CCvrIkd
bu8N9nYjgic415g7XyiQW9C5qHTx3kTUqDbxXgwHd5FWtUTGzWY7Zs6JCJVl2y+lxuA24QD7ND3B
Vbw16h3VDtG4/6NmgIWU+1iXt2gHZ8t7jbokXJnDdwKoyOJ+raewCrlm7IQe5p+XDAydP7PrPfoD
a/pI5dnhPk3tfsqyKQPR2xImxjoJH9atVnTJ6ijBVHuckXlMZ85M0svAMeC3J+X19G6pc5lbyP+O
/XeU8qEkLv+UMv2ByxHqo3XgjVTkTTKJlcaBdEtD7YEVkONazyXRmjlri6gtMkvGJug5NnFxSzUS
EyO9PxPCJyE5etPjjZ6AvYclY5tYSUo8/sxc0prmBKm0TZgrvOgcFgrg5JaHPhg1toyNm404mXob
e5Tho2zdMi74vJb32xQZB0s+8Bch3WgyiRbo93LM1nfP2v9qcAk1Gvx2KvkaQU1Timxe+J8YTnB2
EschwjJ45HL4IiWes2EY0tpzMVZqK3h00oCLv0dmBArbZMyVbrP2bbqhcGjspd3ioC5WDXOXSvL3
o5rPxBYUekj3ocNK6gtIw4BXJvI4acnOu4QhEeNHkARLC10vgjpbNJ2RXayoMupRadBJkYW15ywy
+/03OnflC7DoedEMrsFETTjL7cHWG74Ec+W+dPZwjW1y2T6/G48DyhmC5jArNrvpaW186p0BFTz1
dC5a/e5/XBYAUFEHfACGoQlEt4j/uC+yKUUuvgY3ZJOo5y1tUA0KXM/eD0b0sDmxJWEcZrwuvqyk
Fv7DpFmIukTTjRyrrnqLqAMEBgfhX5ImHhMl3IuzDRwBh740wYsVulWxffGmmiMhg1JbvevNh+/4
ug1rzSuf456lcBzkWbxJ5wbZ6+4spW92CdYPtT52UF7//2Q3S9wwpxOjaq0egxTkDUp4VG+p1Xh7
4MvQq47w6FGkkhTmAk2QLjosJunMbUMV8o9XrUqrcff1JbMFiI27j+0MORuhNr/m9AWxtnT5h6lS
/FPUOjtumsUNjCViqLtP7/+BBu2GOomwUqw8es+enV92G26N0WyrMcAgrwsyHOSlDMiF7SwV7hkk
PLdqgDEPQakGFga+NP49K59O85I9/17wucya4//XoDGHBOLCc/NBarzsVhraV/ZTLseRTfp2DKZ5
+6SloyOWxSRuRD8hVVUQu4GyKtPOzppyyigBH+p46oG90AHE8iNqo5meaYaDkJkaH67Pk54Lv8h4
5a6P2GdVL/TWi89r8ivwNp3IaDKMn+gNN/rwiIocXOdHZR7JNpzLFKzWM/UWicsc+XT1SvdbLWin
ITudOPNHpPumcnI+sF8GHsXnYzHWY19zLdqGfzxmQNRY9bJdGv4kcdd05IU8/WhPs6a5IcwG8TeN
wIE1gxXMpJFNUCESKoxDYcT1Gfef9mrmNYDTWG6epGxYzt3Px3Nds/Qduqw+5AjnrlwC5J/P/Nrr
nQNLCMRfwgSPTBWtCn7uj4dbQy+Jif474eTM9iNYR6s0bcgKxKUfMf5LlvhPFO3zVqW0ho8JSmMr
lUOB/HynOFWmvciTzhkNa9BHHfhk1kQ05wgmy2RcfnWfRfWFfw12CfBGNbJxnjh2uFbcq7GqcKXs
OKZ9jIcPFDjMiHSlL+8RU0yPBCMDcN49IG3GtVBYYimK8eo05nt4V6xYl9vsP/D0ciImJBxqdPfA
k1GWGkPfHAX0vFAiKNO1Z8DiC1VAJxE+KCTVMMs4SUxtBG5/YEwQFbY8nYIPHwkk8hGCEUuUy5Al
hYg6i7093/k3J3iHsBBEMOwZiV7hMbpSq0b4T/rsQLpfBvQH15+aFjtQBhNeAhy/mMx8W1I8QrdL
I9C/G25lxfYSqDXNQGKsRcAC6HlLHeYG3CQsqSlsGNdlp2s3YDRe1dK3tzupUXoYI0lzv77HicQY
emvsG7WmpmF3mpEf2BiHS4ce7bnJ705r5sJIzfnA2Vn3Ci7jn7s4BOMit/Cbst+k11dFEpIN2TL9
mwX6/ZnybnuKNyamQoRk5vvtujRGXvgJDR5a+cPtxrFdr+1Wkj+dCfwk/ZvUQOT2SV9JcbVl7jPc
uG68qlFczWZhRj6kAMCmD620d2qpsJSxs3rJom6Nn1mvuX0xidpQTybDUqs+Md9mrM+AtVCjj2bD
o36EGp8vviRly60wcm30r0a993mAdrscmqJZG3IHz0HLQo8I3f05C46S+68HK8ETA11HbQrkZ6d7
1KbSIMWuLC/0zFXD2lxPhoCo6zEiYUPLXTSGWCUdce/nC5CKASMwgg2PjBlAc7ItfWxumU+ndhRu
URnu4N5I+Y2G6LzwSJQZQ4iV2JfOqdtDtMsQlKfppRhdu6gIKT5Rz+bv82Pnld8Nh8nMJ7o/qH8k
bQ6Vv66X59dfsy1keTi3zuPNRtvMMiPpCZRIfRT18sl4JUMhSrsBIboP7Ite+Wy+N/wPU/FGStHM
tjuQkFrTlpqFxF11z2lvnnvMByGA+Bu5JCWP5hmrqTZ+BpJKl/bf1iUSqbSzFd0028OcYU3H/EDu
nltoMbivp1pcGqdPL0DfnsZqh3ypcz6KIMcpmFr91foEySMnozHapkI70GfyveTlAHiPPGH08lxt
SMpheImqoWon8Dc0AwTQ52RlleY2O61HFslm9ITO1q+3fcXPo4bu4VCrjFgN1cJWkKOvnkD/xLBR
GrsyNQd1rcZM+qxfLO6cbYlSUNuy0CagsQjY4s3LdJZXGFAt9CaK+l/kBfKVVKtOTsuhZ7Cwh0yy
iHoqUQXSqPmXNqtRbKfBZziDmoDXX3NwoikzmvMSNaOiNMkAn5hN0iWFEePqOOrw0uIEPr10e6Q8
qw2Yp+qBPC8pEXkMmI6ORO/oEmDRX550692x6DcBXSZFMT665Si8Tp0VErePczXdilxDh3huwqmY
odklPrUBqv4rmnRI8pUFnyloymBHfk0Zop6jKBYfKAP+JaN5Q9jq160lD/K27VYts5Pz9B4vVH17
avjJly0bRQLSdvEtne5An0TsYbacoeZT3vEkp2lLefyqAnXCIOHeIsQXrelDKp8hu6dhGA9u9DZ7
UpTNy4a/pgf4Casx4q+KcHHHfRJvYDqvHBbuhGtprWB1vKNKbhwRDKLJJgeaweMOBhrFRMd/+KNE
vVIym2VxX/SX+x3HpWzR/RGYdh1jrpXylsefk8fvD1E6Ha/fxII92mdEOMTNgUEkgmW0oimfjBn5
dJB9GjOkgAYHXrJh5QxgUSuvfaKAqT5zpaW0bjMfedVdfPY85P+3PIRNtOLvwuX7nl7JIlG/TNn2
1QHGOoFK72m0Ui0t5HbP92vqIKpqrT2TbG8sECBcqNL56H4eFLxcahDr0PUXP1kiKbK3woMzm6wH
64SfIl7leI8gsNCpzqvewByg1/ijQ2f9qCJfgB4sx9gJjByh7Oe8SGUN7Jz5imkClLYQ9hJsX3vA
chvwgmAaZvhWbcFBSaPni0T+eCZlsu52+njP2eCAsG1GkIiS7kKJnvmgXL9TrY0IcrjK2sQ5FQ2o
BdJtD8FWkrGunruAX/cx8kfuhzvKgKK5oTIgruvt5sDWA4xSGoi5Bf8r0VdjV3dAQxDWItBSCQCB
Iv2yYbVOM+e5PY2zEcJLdvT0sSrwqCkUJ0F5UYf2JZrZx/WP7EhmWkqbXQDIIEC3dBSlzU83sJ8P
7JKrHTmrPm47dnuBPf/MLgI5+gaKWMzu+ocXLmtM/hx3BEdR29mIqtq4ESPZZgqna0STQhTjhCMN
8TdLfEYjJtsj6wR48lDrQQvnTOXGQGS7qZPuflSLfBx1tYGTI+X1ObwZkvKsClOXeDWlNyN81Nuf
/uqzq7A7dDnKnN0pkGhw+YTZmd+spVpxGtGgvOX4kfLxZeU2NMeTL5zNmioHjxyIxpnd5LNCwySh
YnVXWp6bOsOYv2kr/mWHi2TCsiDrx5tOassYpE3jXbX3k0iY9vtc/EEzAnTeIAi+0Zo3tToFkWmc
oRMnpmFsOutUm6jBpnKnZKFLrVTTUvrqpUwiamHYprTUuZ8p668Cvrpgm21M3Jg6ka3uC4WY3qAt
iNGCq5LmENnG0SSmP9XWhJyrRxSwczehO77fhyUg2/h2jCLewAmwio0OAE6XWS+7woOw2F7oU4Bp
g+9h46iUDwrUbHA4bZ8aQglLSi/QltWSJn6VXdrxeT3dbQP4+UXeBieC+kueGMHP6rSy0VETUdPp
2l863hsByBSJCuDyKtihy8z9LL2/OHYAaxJSxv/3PjNVCGB/CKaRKGdLgVE5H2P5lvJNSxlU0s1L
rLlEZuS519dzkenrHkjktjVpMDAWxQTp9/D+HEp0oXPf3dk7AktXsUhi3g4YT/PTK1qRYjOVmLa0
CU2D+I4rwoLW5Wq1/cPeHlMkRr4ZU7G1ZRdLT2+IwZmSEyI3xsFsIMIBvKm2XLZPhynSYOEhMJs1
bXo//q3hZGS0Fr0GT97R4/0u5ljX5I9mHoZKZjQRxXHLz4sGHGcaO95KR6oDTZzjhfi/YeqQnaX9
7VGL9gKLN2NpQezJaSHxiSYntg21xGLF8bgyMcvOS2/Q6ncdSoHnm/IHboucUAWKvz0yg76NiJJO
DNzX9BK7Mmz5wilVEJe3zjwdR0wahDr9uWaAp1WLqwfqzndQhL6dZ2uE9to5GREXUTx0RIMPOZj5
WKlEwAKH7xUi0eSEfGeSOpRVzsvbJFQnLFQ2LzDfqDWFBrJ29F4WCY4bN49nsGOp29kgcZaZboUz
XNDrzytNddJwRoZKMWwUilnJ5blgHC2dy53OjQUSORSBVJ9osDcNVfsnU3lisC5bAiLapxt8wxW9
J1B/oU5hpX8U+eOLM8lrHyXrhfqI7MRmwBp9nokbcvFwQzWAi0GZ4DDK7tJNjHXw7LLCwv+tDNo2
lJpiCk4gJrXXdtgtdQMJ1e7/brSwbT1haWPbY7rotKv5haJCe37nRV8i6aY/Sk9KwNYZEqBdZDP1
lsy1JiZW3tsymRsTmJdNBCm/+g30cup/c9rN4BLyWFbbHX+46JMZyGzIXuFLWxUK0+cC+t8h4HtS
V8yAggQiyCt5hLU2KnqGzvsBX/sJmlBmRZQ7uOt5669eicuBI13z9ZyFbk3iMyRHIxZGYn5IZg5n
vL0+qkVxHCQSGPHunNSr1YR+CxZkx8jRU+jGN2yEt9zO3UagXf7jr9D8tihxzmVQ34WWJPljhil4
q62TJZgidScJFjWsURrhx1yp7kdi62Ir6gunDh+NrZX07VEfTOqD45f1D5jccIh55+JV/508RC40
xWEOsLMlWX2HtlBK9LBKrUAjPyFeENOPIvwCay3aQ2+e3ALpEE6UyUH3HQ5ZcbtNcDkWR6mbchM9
Y/2MSr/oH3SxM549u6pOG/L/NGasijIxUQga+oxVUij3tAeUq3lcfuN1KCKdv061UG54A2UegHh+
29UZvkaKqEcavXdOTxc0M4LJ81OMcwJxZlZ4yvwt7qm4q7d2RBTBX1mtdXRXCQbxbp8XCvP4d6u0
R4exQSRg/8Y5sWUXZh4JdagvvuavXLBl8iQl3P2H7GmR5IJURNDOq2caQilyByvueLiXzIq8oSav
e1mNXTc1WNWOaQm6kw81/O3WtgvLVU+A0d4SG0Ps0qctZuvHvu0e7T1z4x6hzJ5XEwsqW/bB0/Yd
UOSaAEdiTtgf+GeUgvULqlllze/SB6Xy8Ws3/5GDX4MV0I3DF7XeeEGTuQfkDu7VrNA+LmnBdNQh
Ticet65l64H7w1uAXXAvc+vEp9N6pQImSh8h1FgxSQwJXLrdRrjJGzL4rEN3gfoOQ3gUAD6hxnQn
BcNvSG1UqSLywYQCwD2yq1P8HcJvsxZ4s/kaL0Jjcv9XDkJPdiOLIdWHzGPO4Xvo2YL2pLwndgPj
304C6PGEqONO565U6Kxrvy3uPBw6kYH3c3wgTGpOZzRjJvAu1WgT6EEmO9fB3ENue9H+WjB8pwhc
t74iD61zq5zvSsJgjY+JJS1gxDFPJjVWThYCka31gyRG5zg4hQkYjemUbrc80ANP8fM6zLvhuMmV
eIR50UQA6HEc43Qk0HuXiLRyehJ182W2Mmol3hAa1Ct7cs+oLKVwzUhCRQtK2IdRuF9ANYnACfQ4
KERrRwbRyhtqSp6yHfSCTptKbdwgUSZ0oyHu65pqM2blVtELzuj405+Uavd3/1ku2sCtDY5nn6S1
OoOZ7LOBendUBk2oAbEn91zjPXF0/7Hw/Pwv4IikNlOF3AeyJT4Hi2+cS8zwi6Hg1hxPSDtfPfvZ
eu57K7TcQcBSvtpBfi0QljiMowWbpb7GH7dFavzXTozySOfsohjqeXpfAhphM7G3fPqcTCUdaamA
j1Hh6pM/GIpZdDGSNaExNZakgZ7WuLbaQHXNhBY/onKgAW8lMwJiwGvqIKJtwbVT0IwsRRaF/FXI
HgjIzx4MuUu0w0B4JbuAqlb20CFbRMVapSQgq7xxWY/9tvRZNAptqY5oeFIyLnS9qV0ECBBuCheo
xJEcHUqeq4WxcjEO+7BZA6qnE4YpT3Nie/POXx10WAEAJYXy6s/iE7h0eKMHBFN8GnVhXOLM/Xx2
FU63KF3BrU9xh9ZytfsJkaC0qBXD2rSZA/MPO/jRaT4ic8M0Dq+3smQt+rj9SzIP1KzTjTytaD6W
ftO4qUuHyobBK3nIjnYFkLg1K6v8efzMCQd9DVmkY1OZZOVNCBu5D7h6IGBYtxdNS4qp5LmJsB+q
LlQMDEmbGx8MxFeBdDZ3KVW5hZl7TKjh9nKIGUDS4myBfPvlK3CpxoQ4MNdfB5fuarfDhDc1ed0s
xntGlinuFkaqk9p7+6864HyT/TbxCUYUctuubzcA0a5Ma8EY+de3bdzssWvMCB3av8M/a6nyEWVF
XzyE/27xrmPYoAYRlCxLgn7dOPRvVvrddQrdnIKzU/+OOix32wvx/V1TnvUOhIwO5el6MvGcNFzA
0BuIR5zgSSs/eB6bTTuiPux8bHb8K+kJLFgzPrfIhNwpKqHKdg4m8RQwjXts9yDdfnJ9l0yAmH4i
BS4m3D1zSr6Xm0rHu7qJYcg67OQbANLTcecDFpMVaFEgqXN2xLzg4UrCj9SMG4Dvyfck2tCV4rDE
3aM63XCecMbL0itKA9KKFirtvmTvg1WP4TQ4tLFQFkiFdHi00dO3EXWxSjqQXI2OLLe1+pfliI/r
Ma4Kysn9tu8wzxb80y1zM3m7G8n9IKwivLA6vLVlCQJ3CqLkyY7yWmdYtRViA8PIc/+HnC3Grz02
RSpNeAXiqRl/OEXTeB/hTsDdFCzFKqp/Ro1btHUZqzFK3jRLNH62GXaO/SvJSHx7lCS8pF3GOlGL
ygbABcPpgZsfZAot7L+loubPBtV5eB54qS+EE0m9ZB5Cza7m6BL5g/wAqF/8dpPWYvR7nVhk+5Ux
QodZqiW2Lo5e+Tp2gRB0zutCd5epfIOuJRz+0x0+ntCxr/sbWwqVDI7ldLvIlPMOFfG6iK9Efmg3
AAkju5MM/lw0l0TTTvb4v5NvGzMltEgp8YPq9DZhGf25iMiO7NcXyN9/m67Fagsvgz9wKFvRA0Cm
Q3TOvpUeoQ+AUBpEu/DOvjtH3Axq99r9nWIqLdtGkniFdWiBf+LMIGzwcbt7aQ9qjsKZPwSbwirr
0AzDbO+/Uo4ZxJ3LrPvvTsMIODa90nV5HZBW2MmY3MmXw+S15PQJROanbd8kUM83jtBb4QZYcCLY
YVl8a/YRn245588+sPwtezvzlhbVkzH0ZyNL13WxSd6j1ZNruT2kBuR7/YuaqmXyHL1sS7UaobpG
j+XaEeFZoy7HH+ywDyz6jRMGm6oXkHgl6kh0lj1T4TckVxYeGzV5rrd8CROMlN+mvnU8RiXFO6HE
b2tEAHDRgPuXVBpG2JiThy6MrYkdHeQVhJJl66Snm/DEV7/DJjF5uF95jc+g83aN9wQhWi4ZvmsS
wQouSmFN0xJfFFfc8xo0BZs1xXN5RLoILcyIRufK0ir7/zdmcN7atCj+M0DJPqEAiBL7LlnZmo0G
dIidgqhUyVfPIoX3PS5FIDl7T40BHyhV+9Heo/f0ARkGQ6GSWw0QF6xVaVbzbnf6Gnth1jlw6hvi
bR+IwO0CxRyXUrXEzYZP7FtLT9ID3I5jgKEcIaRPEjWREbWXEdtTwhfYHE75N93ehD/URISvruCg
u1aDhghfppJJF3nWRo3kPkxAYHXdGKr2TvRQCopxvzm9K7JN+C6m+6va5mW7z6ls+D6INOPldqcP
blBIJN7+l+6J48ntE3hxvH9z6ZuEp0SL94HX49Z6eR7DPK4B+hTIz1wBIJNxNeNHPp7fj07vLtE/
r9RLBP+eXCDqc0GUSnLptCbHhELdB9+Oqazzduy/RpyG4LMdG0oln6h+SCEvCnySGy9goGwRPw5t
sNAWJGhsqO2M7/wQ7KwAcaPAG4FkwQeoAyHt0b65yNpICwDCWh48v920BTwmy4ZRNB2MauXxoAZB
hWsLiq6uxsYw8J6+1lkPYHO4ftiaxqT5orshhN/WMNnwZ7AROoH0RFCzGiVtvjOv0Y7NCLErjNdS
T3dZa2BGjzLY5I3mPF7F3xXyKpx6mrX29d/hAtQDJpxioHi13xgDXjBBMQmoUia/7XVjLb6Owlkm
Qbj8AlCdwg+8gFPhGSRVcE8yU5j9kproNXVyAMdbEC6CbiD7KmVKniylUmqYD5a7SVWWhIoLq4ei
ImH544Ollx5nq+hHEwwdH0ALHg+XcuzDOMQH/UwgGzbRzV9r/9RdtNY6XxmPtuc4PtLk7mEdCOGo
jEeKhy4MTNuAYEQcBf3eW0DKdv2edBCKxKY68Ce7ephug1taBE9oxgDGqG0QqNPvqOsP1uPlQwq9
DWBg21d3tluoLR51YnQ/ZabvK8aNhgETefSfD03SKNLrm9/hLfapBwbz/Tb7ZMQyLYbqJ+WzWPPy
/A3QAVBr+51Mh9joD1OHetsmF/vZNgWMFYoy8t8rkqC83a21KKmKIlAHwE+sgzDQzQe9pMdNdZgl
R40EIfX8HqMArGiEfKW3G8Lfz9va8v5UP0gN0wvy8gzpdWCTzZMc+1xUnVYi/ISQSxqUdVApSLaa
iRz3jWGNjZMT3CqTrRJXKXRWL6Lf69jT2Wpf5Oh/Q3K1FQM2f3RLQBVW/5SBJ2maiF/n3VR2QBaU
vi5GTU2+KYprQeaC4BFFBdq5nhDR1Or6j3We05d+N4q1HrN2UqAMw/iGcPnFd0KdTXY/gcbgnFq6
hmk9qF8R2Volrn+IRnSQu6n0M3qPanyj2bcwLCWIhDGvqHpwrG6NeV9ciU7nAMd0tTgT/XhvPWH+
nrAxg0a9yCZpW3nSZLPdVOAR6zvaWOzBs1QH/uh+BzwC716Jg+lN3/uGFS0QJy6iZrMV/cyNfJcL
LMX7ZhZ7p+x/U2FiCX5E6/31ECKCpQTi/Yseri/WKyMyCKSxAkFOAIvY9bxv0+zdRaiB30Zsy5c4
jaQdM1wttTYix2drkC0xQi3bcQocKKyWyzzVseQz5DobGi+KmfpUAgPby3WSx9DDdSADEKzPcBYc
syxRC8sIQi/Y7u481wZ/H9sAyWsxKUpLkXaG4BRuW72E6y13cpGlCfQRkdmf8QPD2yUwbP6yGqM7
iSgMx9ftx5waqcBkHsU0GZ0PK9lHJdCvvHmffsNQrI0G5wJPDfhCm/E2K7U8rKGgvbpDC0gHG39w
x9YRs2WGXVLCh6Tulgf+mr/lgN5CXH9MSZS2+YHqJnsF9XR99FpIKGA6kWN0bffAU3COeLYedhyx
ufj94JhpgUKBcPKU3lBMgcLAaGaoEQprRcAzIk8cq4diQvQrKAhq6LP17UyO2/KjoFZGGQz3XM2V
bOm7ClGGnZ/PKv6VwnuCUVm5NNAfnuskUoSavda1wNJGFUZ37FHF8+jgtcPXONnYzO3KqKS4E1g6
XZ43no5jU2/DOUboljNpbR/EQSnMZiUfcfKSimR68VVueFCAB9Evu1hL0T1pvpT2eqj+Fvg8JnJQ
MBJjT1Z+NG1nb5YPPp1iT6rPxkVlGdZ3ohMbsYoQ4Mdo3JFYKuqONf36z5cgNQ77+3NI1SqW54Dt
jUkQYp24LJwWdx5OsY6s7kxUiRecqtgl57ZEYXlnf4ItA/RaLXoFCs9qIZdyCySLKRfwfx7dgSVQ
NdvOIHvwSBO5pr/esA2cpiB6rdBqsZJPZN5Tf96gsOmgeVE60yKg+SZt/H+mohZBLlyfC11eM9wF
1fe5kJ8DkukDm+9aErS29TPwGUpu7PlEQ0LpLugDTA1Sn9hHckOlZdvYgseqseUWfjC7v+zDdY3O
i4hiuu2pkhCIhwEMBIMTrXsiv04kpCWA3aPYZr8CILTMoQbK329U//mtZ1D/aDs934H9WqGQUVRA
CT6qkjCaqY7/nVrnqRefmEFtmVfeLIn9sRkssyrRt0ud7+B0tBrVRb4UkhSAHyDSHEJpH/JzotCk
LojQIOgT61wjYWotoX+WzZhGNannMI7OiJ7FJwPnfOBSm/Jxtk3cEX53KpuESSyFrXX1g1g0PZW6
GNq7ycmpT6gpAxlAyptTld6g6OiWBkQikUyBa49u5x3U7wgAnlKJ3iHVLiW5fKS+iSaFQ07rt7/p
Qzeo5dPsU3qk2YFWMFEfubCfFYa9T7XMl4nmvLOXaZcmfaTFxo0wQ5AHWIypqYQH0Rz50qY99/PH
8ijULqUTdZf+fOuMBz+ByfiAajiP7YfA3mJvzIObcPkJE69tH4RmHoNHjkNDmGf2Vn1T3SEq6owZ
LfC0R5HjVx2IzmU+15un+mOut/3btDb6jDZ346QnM2WBNXPmU7gYq+fmFC7Ak3zZLz+r4KnHo1/m
75L0nSXaREgD3hVgMBPtBivtbBWvHNjJJTzVsD4YQBZmkNBPuCWTxJFDQ4N6/Rd/h+i8N/ngyIlF
VEqNb+h4ITDrfOB3XZ4w1RYrUeTxw/gOhtQnyc9hX74q7TkCxi6RfcFwz1Bw71fVloU5+isZseEI
iM2oBrwwsInKR6qZvhSz92Ygeng/4X4CdobNMFLiZ3JKjLBeG73+2bGW1Tp5aF0I2g69KTZUiPtE
dNNmQrp69jkfAIZugxrubEIXrglAO9MkRr10UOnA2Smw+SB0SEFgLJiv3+cYgqojwXe1SLuZXnBK
f3JwfoGcXzNhx9APyEiDo6ktlpMOIqC/OhwWPSr2+GS27L9zlfSQu9QrteHzfvHHcXuxmBw1eEX/
zKjWXncA0WLGDTpH5fYVG0MLXSYrrX81IloVrQ0oc/GHP0Pe24+EF99Z7Ww1ifEYszfJsDow6mbe
TbECXEcoYonjWvTjg5XbFJCV8J6EPM2v3TPrlaLxjumwA6cL2jdEiq71u2brzs5+7gkSR/wuCTSi
nOZTuV5xOWYKGx9XHpfsd6HrG11xIO+AP6qpPDxwRSae8bnBWXT07l0NvBRa8f2ClhZMkUL9ICdT
gjdJ5KyXom6vPrULgmp2a9h0xtdikmCTMXPIrqmMEimQ8dYsxVAhvAvnox1RoQCMueHCLlKKnOYn
WhZM8APZJdUFeGP8ZTPvKLjTd3M8403sgdMoN4Tx9YmYxLMt9efg3lFqgc+/+i3QyWTioaKx8ONv
De4+O+qtR6wGmR25lZqPqEKqKTwpKoojITMxk9LBu1KSH6x1dKL41IK0+2yV3TdsxXD5L1Ba0YnG
VDx6Pa/PCbCvcPDH+hEAgx40CRQVjYu54mfNZ3k9z6uqidnYPcohEc8aIUWQVp63LkhV12zwWa93
8Vf58wUlvj2HypH7HnlKFejwRlrZ6WBot504r4JMaxTaMP5S43UrcErU15JIIKNE/sLS84aQyALM
EA8kr0MvDhKnZR69ZQoeKcMpCY0RA+66QTPybIm1Moiq0X1H6VjoKfzAshnvJTwa0rqdlBVQwFGv
B1beBMDgwS6ZXMHjttXtgFcA/sNkxTMZ0c+ssn28cXAtnNp861egoJw5v5Ivqybdg8sYZfRrJ6FD
eEKMhIdBSu3SDU9QRob8cHDXPVUp5U8OmbutERO88CpX4dBoA9t8x3df26WuS2Rybxc4fnF3YUBv
5+HKUwQV7fLZEFSG5c4bx317CntueMkvaSDP/dbHOpcq8WSjyIAOXoWqcqcV+cETh1QRup8aHkBy
M/1VlQ5wZ3bAgNOjHwEG0PbQH0UnxTOIZMDWMXb/sXfQLWuXy/tf0EdF9bLxNnPdX8f+4US4iNH8
lw7Y0xlCHAzt9BUCJiQgDWt/ATENOXn/xnw4HbZ0SWv2u68i4QUPJgNekwfS408NHuIGWe2G6Ua+
vuhnnP/Q156tUVq3jwpMQIpgt3VxmNaJKwkgPZTRyxP0dvGo8gOkFG9wAdYY5bhFMf5eC5JmCFy0
iD0y1arGhmHbO+g+YJlC3po5jDZN5gVmO+ZJRx15B6DJ1mkdwl82MsFAN0zO/z6EutcX0k5fEiDH
nRRm4IOoyxbUmt3WGhzQCghUi+i7My/NKThhk8XPYz+zDN5XYcpv7KgMEDvWntwWbzfiP132IllK
1yJ0L1yeWMJ+vNo44EC5Jv+hCNKRjHFcKXl/t7fWhXtMbHGh6HnPkVoodglGiWJdK9tYhfuQLBDb
yUvQrl9KQDQA/Ld1kLQUz43hoVpgE57+PX/Bwp1r+WbTbzlYDluTNofE19gEzm0XbBko2jo0u6wa
16WlTgYb3iV+MDiWgzX43iOtMbWmb9/udUh9ZBGa8My8ORLZhI8gve71lUPF2GpsXcBbn4caHdnx
ZAAjOustTNEGgwIvVUWVHYypjflgBdSfJPI16BVLxAmhSWZ6A0xCLAZT5sLxkiYG4+1a499uo5zM
OXVuZ/zw2FS1yOFsIuQn+mey4XLjFNI4ymlvV0iFHXS66R51Dw4jI8GK+7h1uphdUgLYEZFWDtbQ
wk+zvf1debuFYOua3jcw211A5XYyZ6Tg3PKBdql6cpznnAPYCWOxvLlMfBRyg14YJ7V3571YSwZ0
eUFwEEzuG+thzNLjnhN+KR2ZmG0gRlPxGyPV1N/EcbNq5F4cjhDqVL+eJnez3DivX22d3ISicMiw
FF5IkNC1I1MdNj8RFkBah7yI1K4bMQ0oo4a1IIjnA1tjnAvwVCg98drRkW9alRD0qGziuXv+Sg/p
GfRay9LqgU0FuPa2w5aLC8dczjVh1wYfjPMf02qRuPIMWeYvHSQzbRXyy4Q2zZGRnJ3zb7dKtB3y
QqiENokG3u3HPnYe5xZytbuuK3wXYxOBSwz9sbeMcx57tufj+xgQr7Pd1a0NGqyisby0nSf5ASYf
U0mxI+MfzWmJ+ERcuSLzmx9C9leWbXUU72NCKY7pbRmwbAYLzIPlpLo7Gv3hIvPU/MFF6e3hTtWs
jagT+apjs/Epk6lAJfCoXrqmPJML7BlJTi4jGE9Lyf7uK/o8AyOnLYf9hPn45SHYLXYQgVDipjMK
qOMy6/nL5j5ZHfymok9iq/int7gfMk25IrgBG8ugNCLKCddYiKO5X+kPnhLllheOE3GUIGj6QUml
+UnG1ugSxFDvDufy/F7i2sLkpab6pmAOwZ4d5bXpFrauQ59KKTNf48glEpTWCe0em7YW/qY7FWho
rwhmP5yCWTK6DL1OGVA89xR4fhDXYCGHyoH4/7hziUcbe6zCNBqsi5fGGf6eSwOrfaHnSRQxVvgH
kBaUwNkc3c8UJya11kyVMRiJo+pAE2R4datE7TamQRbR6Peoz32E9Dxkt5MBhqZmAP4YS+CrkgJ4
jptjabZuu0HRzcfilYG+4eRcgm9NhDxtDd4RT3zFhm9WGtSM94xwk9QioN6uKxk1fM5lwxdnn+kI
4H4KM7TNNZ2IVZXXMwMNITOX9sJtBYvNUUifeyxFVnE1mE0hf17LX+81+GmHPsd8KTWpm2KgwVRk
KBPLNvjdMSKeJf7ufodXnSppqRkJxw2yIk4yyRh6hszI7F/lA2ssZpeXppRh/88xCuDKF8Lny3p/
EQZLDmsfAcfNBirx06jsUJupUn+qvRw91Zq8JchDYJSUqgtzRT2zo0dhh7x3VU0ApCHmJd/nDjv1
cigUCOWGn8wRYq5QT/377CoCZ6D1fQiCAUEXFuxuWQV5uCJfXlXrwXsqv5pXcWspEsiXo51pIrsi
g7OT2t4bt7/dj0Q2EzzQkcRGaZvBaUHQfrhqDkSjqcXw2OoMxF92OD1pjuEIYWz/dlgqN3zZBS6f
i6z6ZngWMz/vxgRn8NfJoFL7arH6fKWRDnuG/ilIdabXyVBwueVyrshkB3cts36DEOUjQ1pGY/mP
6IL3kPhu9B4oTh+t9K6rasCLYda4/Gmz8ODSa2wlQ5YOtZlJHHrYp7fIn/7dfiWWqqSgpdVNbZv7
VWu3xt3PWfOpLusPW5m0SahMxSG0E4RJUWfkc4U3Zn4FxSLPIBlE7AU+m27ZdKI8rs236nCC0X/R
lQ67eGffwKDIOuD+j0kTC4BgppRyvihxcAGhf/yZOxpgt6+VGs94p4iVgQBZOLGhPC4S8lgU8EY5
ElUY8sHkbdWoOMQ9tKExtQOeDF1Q2q5uDYXw/BjFqg0zV0M6NI6C23pWrefUwAaQnI91yAmERBVX
MQfoO/AJ7Q4+9boQMUisHy2l8JCQys64Us+PdZigwIjbVPt4t4Xe1i5GOok/iZLTNnVLk1kh0TdZ
W5mhlT+5ytBTGPNjqugctCqjCoxt8RfIww0jLWT3N+JSwtR3wVcedzM8ZWfd0yPAnWzmoY7+ecps
5p9fh9A2ybcB2s2aW9ZSXeHyrKVmTV3HtJsoa9/pT/RjCh81azrb63vmiZA6M311BNrweJl/0Sjt
oerCBjDy8qvIJtx+7+KX2H0NNUoLXnk5QyWLndYudZTsiBESwZvI1kDnoijzbqBN3Aa/XdRQ+Ckg
spfUkf1BfK5DbqpLPxegNpHcU2QGofHPxcpu2holZ6vOnox59WWYtuEBl3txN1ZgjDc61Y+6Ypcz
Ohh/XaKXP2AjtYkRWdcr1Wbdp3NEWEvcc++XeqL73q6ny1VGodjkmUh2FQom54dPuVnNCIcSsAS7
VQY4fkUt4XLjKr64BOFEovAutCNCJuKLPvfilS8mDDn1M6It5qeiGPf46842wRX+R6H0Alh/IPG+
wgcnXtDuJ0xyOCfWfF7GX8M+HqfbKwuD3IL6IKM+AgyDV1OA6uGMBBfXtoyVg2w2/YcXc0f5xZUG
y+SHG8fgUvtfHZqnY5UyhntloPQX5/IBuNbBhoAu0YI8S+M9ijMcyd291Y662p2xemweLITnCr3Y
l9FFCieEoYiWa/27QW0RMgyLpHApDcu/Ik9SGjU7h8/dI3menlgHtd25FqfzG5EW9e6zqgyQAL9i
AB/PK+w74E3AqQ7yWFNdnGoLdhSPZj13ljUFttFdZ4ZaLzakf28dBVq/LgNCw9PWbZBQPjGGfJHA
T/tT1XJTtmuSMsX7gfB/jWOl5xOlhfMhYQf9ueNKOJ8CNIJuqPibPP6piYaXRVggWJ3hAdWV+i90
htTfZvB6yCvkaIpJOT5QoukXNYWnQuFQo0MMRp8EfKpbxsFD8pKNRyrUeTH70odYlP7Sq3ocHYxj
8frVL1oqAmsP57dX5mZ2EcuaoJl9+VaWLQpR9OiEKWn4X5X1y+vJ8ei1th4aPGCR8nqFALrAUWN4
ZVX43QLQi6b+Zb4p7sKveKR6pyXo6qdqTKLJBVpbQ8irrixTm9unTWSM8KZ3gNf/aU7PswwbYLAs
suEZHyTCAubRkztcdgcVUaizEbrd7lZaDuBcS+tCmPBPP8FCAZQy4a7l6bxV1GfQpdc2CYE7WHcz
G5Mws5T/ZIcvij1fyZ/2uy+fgFCSiT24it4JuJOg0B7c14BJZNq3UBbQgWuJXmLyMNWkxXeoSiJx
/591zKUGfN/zdfYzpnh/e/fPTVN5GhD1yaGYVmpwmztLevnuO5mbSw1rkRy8BzNbGF1N5eOPgwKX
u4EH6NZHE2nse5UkC7FGBXC/VWhfPMm4n89kOLxO7qn5AajMUCa2YkiRWcp9peuKeV+NePIQEvuj
aU1j6XRESUo4tidNe+ihvhsQNOsN6rzCaPPyg4eBthyHYc3hp0LVKQzaGsYHxEiueRhl18bfv1iC
WSZsCPJi0Zzyv1Pin/CqYdPR2k9VO0M9mqUuiSYjnBz/7N8mJXvbk7ekU5nHIqaKooiRqgJxg8on
V/krqM5577sP1LELgupvk4lkimw5fg2r9bmxy2vTHUhyad/jKSNmYTusRT+oknsxkJ5dWlBFEk5q
gn+dQiFXe7VjveK+4owc1W+RiMwmlly8BvPiQdKCkwDS3FPKNNDN+35mycb7ii0Uu5m4MEkcsc5b
Arym9UfrjFJDPIQqo08DibBMimMqSRMA9Gbc0PFGqSAWg9fipxpycaFTP8W0t5ipbZHfSHZM0zvc
vGQxrK8qLFe4m769I//TPkebw1b54Pc4CXw903pyiCIoUYPQMGvLhrPYFDwe6OvuoLGY2OABwACq
Iz2IQqz0MIqHutE9vPwaJsjDnGUTwJp4zdPM1IywxqOLTTugMWXvvmIr42HrMpNfdko70OuDxKA4
pjqUeuB8ue+xpeoM/fiFw0G5TatskmjHLlQBz4fCTnlewUNC3To7kJJWwvcQ1aRnlRgTAtqhSjWk
VCEA6y5KoXbwCPPMbOCf3egwdf2KU6tcXg//5T+4M6tH7a281UDsGtiLNvWe39d9srgOZIork+4n
awoUXT2HrSbsKsbPhPM2u9gstv3oVyEYyYkNf3hAQX3dpOLWk/8369JLUt0vFDYQ3B/0KakKcevG
haPBaWhhf9B0tQ4eoMgz/V/ggB/ub96/JCEuCqzC07W1PzeKMXa/Ja7/BQb1rQF6mOz66Z+xuwDc
C8OYL0butcUX9ZMSdYHJ3tNljD5Ap913idzAhhdpFfQoFpOqkE/x8uxKYsxt1oMvZj8/5q82SjYg
8C5txgZJ9BRy7Or90hzKGyYj/nnI6xNTplJqheUWfNWf+kn0+KmgkpycBYKYFhZBJVdSRnCLeASP
U5NiQwb0viwNV93AcArPmFGdwkTJ0XwXLPQvuaD6TIUugchp5mfYwgsm3pAXv2Zp4mg0Vf7WHmaQ
inf39zY8arm3wD3IIJYhZR6qYHtT7aoRek8zV21O80XJkqapD9hdAVw+550Y9HDbYN9e6TU8lRUF
2t7Ey3y2zavtZvum+xjC2Gq30xfOtb1Nz9GyCF0VXZBw19cYDCgg/JIPkBb5lKZkYOOX+aBb3mnu
oihhf1RnwEWCDQXied6xpsdQkZu+vRnTkJKVL3LhxdYKgyMgof6/c00CfJAR6oAZ+qZGyPg8TrXt
806OZGgSe4BeJIaZkNskV68bN3mBmkaSXlwhWnwSXP4XfZsNH3dNiYPUEZ/etf3EPxu/eKxW/yWD
plVAKVtOMNSjIrmCF781zXnJ9XvX3ciysavQgBE2BbRQRNcM44aJxnrLXPPeuQwLYnD+cz5qs0/q
jRRNOaBtonklJW00mX3kaFgyhF8lhiGZ6UWFd+ssoOeqrzO4z79Sbr19qwOAJ0csdOTvxYI8QBA9
YRkV/exW4O8tph5/TC3/Cm1bViAxsxaakB3RKKJnghgtdUQGvW9epRiUshiDqMiFEw0fHCUAJbbz
7DHr2ORdSAM6w8MgzAFuvDqa5KAQ6U+64HLL7kr34b4efmSBwwFC5FTkzPmdVY24Tb+VqhI9l4wP
WOWulOaqzAIKe4TF7yWxgpFhxQI9n1x7eMBNHYPBEWl0uOCXuR7Yn8x3kMleZPlaeJp46QN9hEu7
ZMioiEuWy9XLFV7HxE5EBgwUzN0lE8j+nnEb02riDArMi/oV7TbUy9n3sXTBrLGZkD2TjJNm4ujv
VsC/JLfRQsB+vT+kOhbSRQFVnqEPFkC1LPRl9qSy0x4/qnh7kd7tQiu8ldxKo0zI608pTRsuD2Ar
sdGi+HA1zRYe64sDDHxuiBWErip6RRJinrw4W0vMT8kw1ax93idnO8Q/48rAAU3pqDPq5r5Pjh4M
nBDIP0agCzknPxMm47INenRzVWwKsv9OWXdgvLK5kQbktPveTbxHh/yBsdqF2wiGQNo2LjEImBKj
ic+q7i05dAOSu/jUOnYxKofV0TPf6SppI8jSs+9yCGvuMzxSIhArWy0XBidDfzXq4OLgFMw9M6Cy
mcH0ZL2OZkhghkEGTVoRwYfgL8+dwPMHn1jl4oC0MV9NFktYA3FGEqRXgwrokcy3SVPXQmB69ed/
u3GkeMOoNSRBSmdggnhdT+W/XVLRz4FlMtezFPWnZ8tTHI8iMWrV15BuWk12u63fx5gKa57lBCuT
ed/W4ZbXd88ARB6kCcQl55asqjk9ZhBHFBluWj7y/98EiNt2dFNmj2Epg01h47bytlY1GNUKoAjG
AJQj/iPiLL2njSLj0UpuRxA+5Mz09Rl7RnUkhl1pRLBnHvPFuLNhivqQdQrk6q0S3vwPMMuvBsdF
fXm8yheTVVvnFSXyVRNUAq38YV4ZazJP8441P62InO/bHv7rTMhnw2FOSrprgdKTRTbQ0t0O+xso
IZH73Ib4jm+5YrTcuD83VnbEqD/kLrkNlRPmtANG6rCV5gzPU28ryte54RDYTxX9V/XLOD1kkSWU
JyWHaVZ8c/0UIWrqcpQGoBDq3IGcfdQhmzpvBj1B82OyQGEXbG479q44GWB57e6D2nwD861R8WpQ
dq/xAZQx9PMGCbMZe4z4VlTUEU1THwJhvSZTMlab9NMXfiVAJBYuF6ed//JGWSlsfWhx39r8j98B
cxAOUUHaiQY6S6DkeX9tJz81loiMWoO1fQAkbG5jMkEy4J30jylpKI/hkbRcQfMWbMLV6EOzORIf
K8x4PA3ibgzA3z5oOTC/6lWS9y7Znwmf033xJtX4tZivZQeWRPGmuSUL5kCwsY7bMfAncR6xWPcp
Kz+1iLMPHUc3Qm3BExDpmH5kOh/+zwSxgiBLy/CWVnKo4O9gXMDcMUn+ovzWS9//IW3UO9mjcqQJ
A1zZ+lTV85fHgEyhCKVa6So+7N3zBWcw/YWGo61eQHkA4TgL3IOXXHmi+iwstEiS7OA1W+xM0QHp
vQnx9iPHdTg/nYXhWI91Vm97wHm18GOmqKwBbL64PC8mFFlSgRNCPUajo1e0h5+wG+aPzM4dHaSY
/Ro/TIIcFnmynLCF4GtXBZPcUxWzQ6/MW6nU32yLf98KkHecWlWodci6tSyH/LE6wgy0bU3JLP+S
QzDNlUI1pypJjHkCEqBSKjXBXrnL+gVSDrsgbCQUFmzQo0B5B9NVpna6t9tHEnIBnrWHCEfw9rsK
n/4dMsO/pQy1JhtwwozhNutXAHBp9MxCwPx5aFieA2uUD4+bwg0kW9teRqo3uAY0vE88cz7RYvU9
Q7xqnxzC+xTdzh+UfhNeq/fYexa7/BvX7VIp9o0mPMIlJeb3iAON3D6nQA+KEgi8XfKpiSCrUjSu
/4XpO/DN/ZAdGKbR7lQ7suD3/+UO9r5BxdpnT/OWkNOdjLmWXhPo4bctN8xIW6D6XWJppUG6ogGk
klSfCt82jSNcOUuy6y1aO/jWfrIH4/6jP7dWP2hkjf62hdLW9aZKf5+O18L33vZ6FgqJ92cxMKOl
tvm3JQ/VlSz9bo0REs6u38f5TKGkTSa2s5qBXPGhRPPC6NIid/KSfCncQSzDcbsR0L3j4u6TzMDI
t0Zhn3yDdPDOWTAmW2t2fq0FEigGWTWm9k32U3WM6BX44eLyqaI70TlEBxBM6usubDVAe3kak1uo
XM1cXlw8Z42+41Y2+qwg1NgvyDeznvA68MeJDy3mqXgVEAaNcxH7BKbIA0pPiXwFf5LXXeIwE4qj
NbOKvuprbWZZGaH8Jg4Ud2hcZPGzedBPY+36W9wEir6Aaczl19U9OT2aGM62ZIYpBKOeXl/Ba0YN
JV2cMGHV+k6xlMnS3Obg+jNizuGIe4uS9su/BaVVmCAb+sLn0ThGPyRb77HCNVzWmAelmOM9S/yO
u6hvjg+y4noGacdun7pIIXlB7RG18abHg261OP57gElV3HpGcdW7c5kxd0PkUcMi77ud5chSv9wd
3p2uF7KM34YIZ4KM4K5WGSZCmxN+SHuNdZjUDjdibcAshICLS2oUkp1UDojK9duL3RmpVPVCJWV4
B+7KSndszdavdtAwu+7TAZbCvLcI6TDUZmaug1k/u8qqO7AM2YyE1BhTtN5gSOaBhhnI3vkoFOKW
4hppGoiivwIrBlbTS6IEiJfw0y4tZTsmht7qrYr/TLe6Kl+6ta7im7GHKv8pvvecZ64ZxI26hG3m
XsfiuR8//RAWXXNOzEAXsaI16KNgt4VyCXlUzZm+6zJCYlUnL1KnkJBMIp0bYvFzKnYCFwhJ9UDQ
6Xt5OAjht/jLlVylltHVDv/oeohfwqVwlfT0vOVsBhFmsuGPt+aOOSKFQ0+ZkFhYhBcOR60wLGYY
B8C0qu+oSMMbAml+6pZjtB7tbGbxn3dy2iQ6QpI40H1Y0BYI5IOFA8vaFhZffOUrNymSQS/quNay
sRpPhmjbhVPOb4L2oJP+i9B7CeWD9xcjXFqDn8a3G0bK1vH1/C7vSWl5gkWXeudIg3A++N36HiYS
674+pL6R7WYhB5qAIMkHjb5LW+oOmxRS8rRB19P6TkyEv5shlJX6EBE/VJY8KR6dEuNRFnYnpMRh
nT6JKfk+r3alGc8C6JCoCyrfiOEH0Wtxy6bUyPE8ll0pQMgONRG2GMBNqJUw4CnuSzLvsN9xSx98
TJNcOiryHh57SpW4E0yO8HiADvAsExr1k0xuYG2iihqkQErJZ9/hqrRWnpFeK/EWBtijgYgRLu35
DPGXzQAM/hOhi+wum3koeRv90hLtjGyRAe+Fbzn9Y05S2jlZuQKIbqxqf/xNGYFWxwodO7dqMFYm
uF1rwYECPZmx6hV5vkNwWg2IowlDmwRRYIIe/2yhJkCzhboKOC5gH6NWhQTMMB3qfAEXlhQHhBlI
JSa6tZzOXswkTa5j6rDst8mATzQE3K8OVg1H7aCNXNEUGYF46izw0Bvg41HjjS/IFxi2gKAJeKdG
AwSjaZAZ31MoaX6LH95QOjQxqFPDH4Iel2wPmyi9UCV6XA5R+vJcnML3hLtkIxljiqL2QwCwu58o
DPaesb5YmZQEL/WednPxXXeuZ3s+LsO5/l3cbIttBUq3jr/nCvhfVUbZ5qkf1kYzdRBiQWRoOJGP
54JJ8SeB2vqKY5Enn7O5s4M3IkKSWJPtpC+J8slir/WJHiWZRdnsyQUJYwqMF4dSm82kK+yzB+PR
LY2kbLobp2k2YKklz17mZx2ngkh0j34vxNmoab7m8I4BBjP2AFBrIaIgOYVdpd4a73yw78vbo6Sh
4NzFhyTYeQeAoSeRmz8FxLaYDx9s82uGIxN3ZvPUBpqyK5INDQf+/jxH7gwRsehhS0EFOSdOrNW7
Q81PSZ39nZGWWJ6GZzGaZK88WZrXQH66Ysrtawtm0cjoEnvXUngZ4jyOFlmJB8D3JlpnL7CMogBQ
2jBDG/WdSBwHhkQfbEEJCigVD53gvMb0jODUlk/QmBm7jc++Bko6chO92cW2RH2xDPILOX8pLr03
GSkF4ugbUxLsbGEk2QwbFMYQeV44FjAXUj3bLDgkZqxXqHcTR6C4ooa/m9pEWI8Pk5+RTj+/ikCw
1Y7JO6SVOP1dmCXhGlxHfbwZ/4HEoCfMGFLVbZx1RzuNpYcXHChqIPD2ZkOceybTbnx9QMubRyiO
34GVZSU13OqfEmjDuS4a8Us+6D2XWxY5HiQeWYhb3nE+X2eYy9lwrx/BTDNJUejz6VKK1wiAkpGy
SUU1aQH0wivFDDUVSuhv5EI1qg6qveGNLLUDBseWtrI5FyxjZ6wRtpGB4Qt5W5vjg6uQxBB940ei
e65WbVATO0lNffqG/AeomYiLIGVTIS88D77OG/nVY5kdz5yPyAHs3xFeF2W51rzdGuilDtXNPJ9N
xXhmBfnOW7gJjXvyXTcn3W5E5NKgXsqgXcp3RiXKbs/KR8q0gH5x0j5hEPzb+0Zt12TRaG08zf+8
9UdtuJCI6CG7MRFEVlgqNS/DHRQbBl7u9P+HtGKU3k6uMnIpNaNFZD70UKTmJfWaBAVZkBgy94Od
TnRBXIoHKx4hZekyAF8NnTMic7jDajRE61vsBeSy/pQ/+V/9bSDNn6ld5BJx1fd1W31rOluI1hFd
AhP3YohFCbL6bag+o7td75vvKevweMS402WCziHK2tp0B6glTummeFlSZfqT/ajk40hFdsD50NVE
019Xu6RaSJA/k71XrATIF8QNXN/EHPuMJ/sFOUMTwPiBY5R3h036au6wYMZhA8Bwo3nuCcW0eg8+
Uls2SzCG0lX76fitiSBaU1yhZ90oCSjhunaBpqwm6HsU9YbaxicI+V+zKfOGnkJrcrGRrYVc9I9l
qHeCdKb9VomxINnMjAg65m+mIleaAtfEN/SvleeTZX37r1qB1DMHJtG6/xRPbX23x0pNw0tht9QF
SAj+2PeQ26e/6PkEuoPjzg6/euxQ/PqF8We+Fhl9xJqZrsA/jXEIt5V+JOtccre1pBJH4jyuKwIX
l1CimLirz/gl1QCLLWTpM1GC23vIaXQV33r2Nz6Es3QaTpR79kIiuLdhuL3t5JbY/h+Z1qhEbhFz
hWjTrEaiUP6MKcJNEkCzMIP89V90uN4a/VtmsiLNbdUVfYlMvQiTimwptxBSBvv8uNbAw5gaiLpe
7ClWbaKPfxKiUi+CimnnMug1buw30xywgA/DCtQSoV52dPFCudCsIshesbozr8f8IqWqNRT8LJQK
Ak9dHWDCnec0rzHOiQZZtvL2pa6hXfcaVS0tVWVYtKpR89KJMNwscCdCRrwaM9HRWZ3Zqxsy287f
VrAL4/4BiA89DnGuH/XNCnxvTMNEWjZWMcXiaatGXWu7r9hq6gH86ynJAPj+x8qvwdCfmsXRTgg+
1VZog+MmI6xumFVV47o6MjR9eBRKZI5hHg8YR81aUvCtd67ztmp72ek2eIkTp0PprCz49rfqRHo1
5ILaOmycD7Dz93VUyU5DArmoCkPpXoS0x5iaOhMma5RimmFlhuQhR0WQLIPeiSQ41scimWBx4eo/
w/AtWETwqp+ZoFwZAR/82OI43QWSmGCBq2qTrSD/GhsvPlho1uJZuI7gvb0FkF6SodU8KAAf/XXf
h2doatomMztxOwmqXn2SiHZR4WjPb0tS8FdAoMeM6mcQyFLmI1w1mK4+Qf18T6c0wTFnwsFMBml/
puGHF/RTKAEY8XpEwchMfcSCKjbGbqCBQb7YM4rfNbZr7EUB/z40KajGf0phCTT8D5H2ZgCwdiO3
ho2Vt+nNCLOgBCQO8TbvKxFWKZOvi84VfXAMPfxrj3rr6M0JCIQiBL7uW9SvozShQIMoAOry1zjt
bscICsHynDnESSgQEEIdWTBroMCwgqw4w9HnmN0JL9U3EvUkuxHt74ZIzUtZtOnMMUz7bsUjuMUW
Qc+bfnpk/c/kFsJJO1Bn0Y+8ItPj/Yg213iRkv26Puv7tBKV46pvzSWhCXy1VOB//3fgVHUyOB2e
ZvLCUkdgRkz0DSKLZ8ajvwDhoLaU+c7h+PB1ULFxyoN9TKUwl4WnWgC2C9rAHkaqgewzNCHajk5o
iwhNPqdRJGMj54NPKfFtuaSX257yJwNeZJiAQL6QhR/aBpOMNyfb2j5h6u/K4v9a+Nv4TVHyWcxI
U6bvvbhR2IzwqltorIn/06qYGHQGzn/9vmP9SreD281yGnL7MQNvG9x3U/Biq83JCL9ZDTVeIBDB
Scx81E2sRdVRrFwBRe/tKli6PoEmM9OuQ6Hza52zJZoTVM9Kr7SB420TPjU5XTaAbY7yWvfKwYLM
+aQIU7iMvDK5Cjn80rnkvlt58UuEf5uuKg4JgSpg7tW7V0SaYPp9kqm1wPl+IookjAeNRTkIoUFQ
G3ffFkQmRZKzepu6KbEDow254fwxgusfrkAsm5ZmXUWXK48ieuOqeQ0iTS1yYmL+ZKfSSO8UxEZa
zBEjV6tMy55dLVwU83+1pcbuEKg4QmFZODE7/aGN7L+es5RrLAYCldBgHJkKI2j1FOmf8G44mibp
EymVNwsdZ1jJ4rwLh0rE+8CYBmuEAQiX0TeH2wFv+f2YWmoX18+v4eCcI92P/9gpT6Niwdx0Jywx
uVXb8Wa8X7D1xMKfgntH/0BQ/HwJhMgX6k1jQSrmcvf8TO+NfLqpONvCRiGlQu6yZNDgVmT0o3s2
EX/kgD1qIBzU1ddnbcLn4KJqQRBXVwKZRKZeZzr5NKojjmqB9NWKkorgTVRDRqojl2wMWKAI3b8d
v1ANDV60ZIdcUhYr2DsfGnhrGwvoYs5MEph++v8rNJ5xdEf0+Y09B9/xzVSGZerkmgtq6dE0wIu5
r+hoyvHyK2iw9D0tNChXCJYmPceYasDqY7MLDuCZUgZDWlb3ki9Lzj6/7U3Mk04Ae1zsZ8lkDokF
AJSL9sEGd3Eh+/jdAAlKcU1ji5udxnoCYgtrVWL6cHL7Fs2wsVv1KTYn0l3CaKhEKBEtiTFSyBHt
kKcb1FStYi6DdQrujytRtBk4JL3Rp6RpYmrWbRlOT7oNewvpqHORW0mtAqa4/fznuoig9rKN3rqN
g5XbZ94iXaTtA6U7Dg+0kxHWfFy9pxABg1vs0PQVZh+AgPAo8RrDV2M/H050uDxvN3MixmNCHFoL
OXIyuu9XP4SGZ0xDWyGfnUZq7ExrQXyj/xlLsU98h0iSaOz6P1xKZkheRxF1in6CFi4emoqFCDIV
uTGuEsGXkgi7RPYk5Radl0U7lv4myLC9DOSwgwxA3H2vGm4RkqyDnKh7Ib6SJFrc0pSb1bxoxB1v
JdSRv+rngJSkNT9uUF0QjXsbTQhG1Ac691DIwHW9Mt4qWVCaTmwzWY0tXKVNfYLhCorVjOvBTS7g
sNyR+EPYMQ+X2PAbS6TM3KX95Pcdp096njD6XSfeGItzHY7aATJNnyMRDBxyBp7lpJXuG2rx1aH4
MPtnbQVwuW+OgdxMSroO7J46Ps9vNe8RJrGerYjkerjzXZA+MnNZXx+dJOd609wnbROcXB6LWAkM
nFMkmT2Xye4dl4qMUlFQNWWnrr06R19hu3H9HkNyXyg+Fmqqo3Hp+8M2H+3Oal3QJSTOMHhnbty/
KPPqiMOG+AVZk1VEEYmDSdu2TI/xtmrXfCze2ViEKCta4bmw1dyOcearKOisLp8RlBnzATN/6Bfs
Um6LMhqiCd5xQCbRxfrzL/rig2dNPVwJM9L5OvsY1V0VVmR1uhnkpZXuR/VFSS2jRQqzqeGmmNK2
y73PIPK/SIbHjOETr0HzQ0B2mnPTAyRAL0PuylOSb5tGDZks3otVeYF80d3v4lsEWz9H0r4dnZVE
Wd/A+e6lY/+koSB9cCFqKv+uSj7dQwYXF8M1OvufD+EJbrvym+dbDbv0iQ+wGfqLuGhSI4V9j7xV
gMGxlbnIjP3910+bwY4/DTfpe4SxH/ELsarpqPHkw4L1diCsNXZLwYEXQDEsdVbj60/uCUIDJQuY
m77/eiWGYLN3cI0gKQbvuT/gi4qs0t7FtwXragwOjpw55GzJ8/ETwV3AZ2UNCd/1uVSyYL9lbrXo
vyz5vI0QHTSfP7HZdBWKAMnR1LGcl9L5bhlPsmXjEGpKzKaG5emtyjXmgs8drYin3EtEO7cXCSpg
LnBqfi5g/GZOwWPw4ztcHdamour7yh3UjZhJmYE+QBO9DPE+LgZfHp/yypOZUzCutUdXxof1+Ose
F5f46EqrzjRvvtBVZnE8QypskNezZgHVgHKfvNwSzq7GMxOtKQYp1vAuBeLF/4JBr1UoCZK79Dhr
vnqbnbaOXL9aojUpEpwLTp64CqfOCUX/5A2S5giDVc5n8cT7UDsJiroH8z+XOEehCC6HAG2QpZnB
KEQEAQG/k/Kgb+Et12JBHvGazd1y9QDac9qpfy/3wIZXaD5wz1+NSp+V2E3sj00Gog7rZzLEnw4V
K3tTXcYoHARkc0yy0tWYsME027kUNb/22twvGSbX0LCtH8PsY/iDxhOdpfsa/XzEYzgFOVonMfuF
qx2+/tRRH8dOfv52Fy4RZNgohfY/g12kcIiGhIsEEl6qO6bie3QfKmV3ZMgnDVW0RL6RukkwBroU
Ca84Joo9LwCWbv8As24bDE85/EQCSY9B2Aol60y5jM9Vz9scorMp+jA74DwP7PzkF/Jftix/Ea2a
zEkuMFB8jUD3QY1+CN7aGKXgqulbNfhfIT1l/rzII9Z7ftfYRsipWsfm+oIfTXys3iI46K52ln8q
X52+DiPSFXQ8oy50jf1rbW4N+pichpwnN+eMbU4kzayD7N9g8cRpZHV/JaK/EL1Nkrys1uylnTom
CnIYds7VXC/As0ZguRjdrRPFxuijWkXBSIv6wkIhHM3d6C7lsOZlITklWdMBAOih+KAp6P36YNBk
zmKFT9Z7Hru8wQONpK0dIDsx3Z+QpqcMEuBj2B783LjGTIwKO1D0BMMRoOrM+Bu46sOLnyqqnDAk
pvXzPvnGIz/iIreOzLrOrybYC1/TMJkFYmL9QALvOg9Hd453+Ct+fRjOkOVHdDFPXbbN7FDWA4Ui
4XZEP83EKY8j+6ndUJqFL1tkmKqmyo8svD/wsQiD9Skd01UXwU/Dcc33RnME5LXmnpbXK+MGPvHA
LrSrEfAtFgs9mBTofdUc5pixjDrjjXzbNg+xXTo6db98ZCSpPESxWyHtCKl2Io6HJzZ0fn7sJOe2
X3xxJFKNDPeL/opJ92pGOIrWV2D54rFAd6AZAyIP9F4i9Kk2dME971Yh/MEmxX06TIizigYntlOL
Wqajz7MuSyb4Dv3nEId9xyx4lkquX9W3lq7kbpCDJZmC4MKQOio1qwFJW0qbUWCMWSKgC0O1ndmT
5w7thlK1m/Ph+EIfLpycwpaQEvKBID2MXens4vq+djcHDWAMiEbuMorek2SpbLPo8g/I9Uf15Rp3
bhWo/SxosyBJzZdddzylCe0mUVG5iTCuo9y2DRJuHYQeFAe9ZNk/O3c4SDQgDRtmaPNNQAApaGOh
CIqTX42w0OqKu1SEILOmKKyfxeRMly8G5Dhb8yTHN2uK/CVh5oGFdmdpnK+fNJ34hchDsL71oz8h
zqjAbYSRqgJih5K873iXyZcr66KAoZ+pwayjsp+9+Hv1dXu4+BAUxt2uQRh3rI7Hbw9//ItK5EB5
XhINHHKXj+lsNGHGaQolWqYVtGPw06Q38hQL60UB29PjrOLjcGy8CwVkz012HfywclYef1dgmuKH
rfoavmIujZNtEL24ZsmRRJ4NEEVaNvt5tOjj1ZruPzgegV4o3NJX6a8RtnrOzilWH0CijHke3522
+nel4JkiZkO/e8XCUkwOXJmLbcOtLSs/cqk/Mx+7RQLlJFmJ9P0Zn3dQY2v9lwFcolAebkCwEVXq
HYlc2DGU3YeSqZrdz4WNBySyTkZNeMOHO8ozCZ3XJXGVlxGTDEBIVAH1z1ebVGO0goXAesiMX4jH
tdIMfg+T81FtlDXY22bZZAeMA17IJ7yP21kIIMnuNpGH0Io+j8RSUUxeYleKwr/OrKx8V4Me8T0n
oypzLnp9P+R7QZCKP9sSJyBYSlSHAsRRr0rP/tfCHxug+lGtfbW0ZNcvJfQZ+bJwKzG4FrPtbx0b
SFk1KMSfbviMQ6gj8mRAGQ0DOazoyaU5fjct7I1+WQUrvjnhe1zeE2J40ORqNPiTYNVvsEBk79XX
vWTCj+UyTQP53Uet0EKtlZiymqMoUvNJ7Pn6yz1sMDuGObhmXle97alVajpXaDtSfxcA23YaSP2d
kiV1lnxdfco9jVHzqWDadMZBy1D9jmm4arTZj0pENTtcPeFb/R4bZ+VJFYtCzKdpJnaBNndK/EsN
7lCOrqMTU0XrQlRdji5U7ffCfOOg+Rj2tcRqjNqKVPsmZP8aR6BXaO2lLxJD5EZxWRXx6dYxmOH9
B+2M/Q8t3o06p1zu388GHw1nIwTN4PRXVLAwJjg0fLiVjXuCD/Cs2O4ZJqR1dUAv8dig0wJG0pIj
tB0rMx4pD+OHaOwBSFrvpHh3YSh7d+dGDM+IDd67N/3F7T7jtOsj6WKpAcINtAvxYnFFknVQv646
qxoMrTR39MBUycPvJ4Z0Qi5yZSbUenbUwVJy9ah7cf1fHzCSVy/6v6uh6QPu8aQDhCxDEHrle0FM
4JzPon0SKriSCCQQMpf260sZXLeEL+mwpoVe5yCt6hs9nhH4mFmaBS7TnesxAxDK/Yb0KGzc2enI
qrhy65ZuTmz/9IyJElOZe2z6TS0Pq1xdJ1CRJvKkCSjR62oLHADVJDv+jNiSPOKhlAkPo7997Pxr
qa0TqpaILrxxQxWKmoSd+5MCpQRMujMfDakIaArX52te9syZ7WpKCoRHxeSWcxljE9JZ5rBzE+X9
N+8zP9WXtmdd3nk/L0dmPtbhVlnQn0759nM9RBRnnQEbwdyTrkYVrtgCB10yMRHLaoJUgk37SNW7
c8H2vhAj4H5bJCZw3IEyoxKS0+2VWmoa5YHbD3X39yza8K2zRFBr5fEsCGv1ScK077H/a10bG+Ik
qqU5PSPpjNYgbc3q1Nsrwcl/Y9TUid3ownixShc3Nxz8tAGJYqAgJstiDBuJDDB9qeV5pYHTjf2i
ucI4PY0uq2km/OWOLMJ193pvG5BpJYZyzag2DoYswjMaN3/qWExHNUjJrsSjYVe1l5cDBFz/grhz
eg/h0VJjsksXaGbRR8iHiAWxGUIzv+KxCRGqaQaIvNc0WmTydrtowSyWtMyLfyH/J+zK5bG7mLkh
e4P1wBA2pswZE73tkW6yYdfkMZOjLmxPaW5kS6VJD8hzxFfmJVOjIGPDgN2W2xTf1HiVt46trhq3
K90Jxh+qrV6xRKHOGaaNdHt39MmS9lO4M4bJzpNIb+VPkAz7qoL2EtEW4LDvLBd+oX1lVyHTr3oE
fyaEisrMj1h9VJaX64uxj8U4/T/9vCOvc6GuhjTTxge11uxWImWhnLYjWrKzjek8HN8J027uZ8zD
qaXtKv/xZjBusGrnwxlV+313Yvydx79D13prrBklT+yu6iZWxaqjdao3ZuXkKGFWbS7YCmg9NZBh
Br5hBSK20b+WMPs6/B/wTLp4jvv/YwUqG6mtPsVNulgVW6G8mpUDk3k3Knj/nPKFMjU6WjlXFIG2
70wW6piB2kISTcgp9Cqkh6oGyoCFwdvJO5YfEGDFu4DnTCE6SkB2qqi5IBEH2sZ/SBqlGwMDRtNt
xmBuoILil815x4TFUNE8VCoPaz527uyijuFa0g8VH7d5jnoSFA7cRfbkSOdulqch50fZLYKMaODE
eq97VcV+xBlPlYX0kUBAgJ7/usCVknpFwx/criU7HgTqgSntQtlzEgGI5O4WjhSxoRodHrG30JdF
7kZS7AMDxfbCTD362TuzyKfHHQjFsZGDoZ1iJVI7/bAM4POaJDBB0tmoZ8Y12AiAlAs/GnohsHIL
vIzuDVxhodftTgHjM5rGEV11mOnRQGJM3k97+4pFo+nrgHsQY6sJWeKXi4hHQ4lpOt+aC19ZxSaU
cnzRjNy5hOzJXFLL9dt2yooq7Z+/8G1ReteKIkPJG38tpYkdeiVi1ugIWPvNmk6rxVmVgXhW9Z4n
w8jPaEHK7/ojRueKAim1CiIA8beusvJxXuqGd2Ujxq7C/NqraoLpWI60iL6l2oCCDs6Kkl5HzGnN
v8cd9gX07AaDsDn8D2jz3ixiOIO6xvpJGI/l2JboKHpLsESfzLn9o2tUcnnjYCHAm5EAV6w1/1fH
jfBoa3GCcsAkm+LWX/g9QccQoq7TvsdNIsPKPD93NU3+vXhserjue1jQcsgBD4nfrdHh6bjWDFpV
Bg8gKEZTeUyVcgU2XmCcPeM9a3IvKb8SNGm9RSpyYA/PPr0s9S+8od0J3/fj5K7KVderE+DCMH59
TiP9zmqYmLSz3iO8CIXcPMqp9ZVx1QhhbVV8To/e0Z3/6K35i7/gsLSB6Rdf2WJADE4o7fk+TLEh
SKtOu7nZAaCMlWn+rJ2I60O9gfkqDGl7M2LfRgJRcHjNt8bPw+TuwhsFxycyreabdcR6knxVzs5W
Np/qDa7wCyy/KcmpHTziBozVBsMwmzvhaAiaIRIbhD9qGThseXmpERH84nyCdPcQMBW2w6ZRXvTM
O9gXJSouHiOo82XQeCEMMpyarLBw000RwzDtm7qerS/UDfEUv2CNyERGIVKKi8SaG1dbZCLE4Iu/
gtMJ29JbG/3FJ3ddu8HRSscvLXjwMpwuVzchpExlMDwT2qW4HXjemHwGmrkwGbPc1Xjo7UDjw1cs
1vBZ3pSJCbwvuZfe4NwY9ONkVgaSblhJSoh+UfX9BPlPLTKNfS0ltsy/KriQrUK/xJG0w2MW3K+q
XD2pMcif4tYhtniFEL/U9skv8L8rX6xES3ev88cgAPWKClkVCYzH5i1oc9eMXiZtyEdQQxTxZ32P
KLwL6h0IFclq80Mw8QLHFp2LAceGSUhzQRP8s0AmYCyVodtaZp+NjEMKpSe3wvu6VNgLe2twzX7d
hhgF2iZ6vfi1a5fOuPe8u1/2GJWccm/uHQWj8tCNdhUdixCh0q6VxkpRyRTeWIQAJtF/i6sZ8hoE
7rE1v1omense7kzkzdng9yM0IDhWMe+X6xGyiuYqkZr5larOAWfYni/KLftr9EfXjVzstVWCfIe1
Lf7JinA5PsfpEcaHa4scWrzPUXAd7oG7wsKxe/cZiSFTWcIC/dzJTrBiQCFRqOxbkyW8Y3wyxXAQ
rNO4YpIe4lLrLH0LBq9Rez469zsKMfmrpsRfr0oDzYpvVCU/nGlYJAGHhxh8RKwSSAW2EKnJK3xV
OU3fP60CAjgHXApsFGeWrHSV24OAj2vStKvoWptChrL5VzMClzdgluXYKK92aM83GoovtfLJRAFw
EcRWccoZt8/vZSHXtWW/m2fj5UNZozSuBZS7tnAmasZEL4y9h+FmBqjezpn4sgAaBEAlwdBo4dq8
IkTUdMvuoWmt5yGhnTFmBthauOC3zHOqwjM9txrPfTYesi++Ozn5KwHT0Vxvx/knI4rV2fnoBXJc
EnsifjJ4T18I8oknydRgoqO48W0jDkdvXbQwmn6RGDIEc0XfBOXv06/0dnE0Iyf6hbFJ/lnE1uga
NphNtaA5iyQZa8EmABv7faZIF8vNtZf2LDyWrjsT+inUwPn0/60Piv8RoVJTbninM0CXoGJNXZ8y
+rnGS9UFNw268Ozgqz3hcH9+1oDjr9UJdt8xKP7kRoUQLo55A/lfBP7oCDHXiXfZfEPi446Pq6gy
LyohkdQePCnYJPvzBcBzHagmiMm7q9krcqwOCd6bVQZGlvOLtVNyLrOodxEIAylDQ1oyUK1A3nD6
LQdwmnzlHuYdbBKbC2t/quMztn9eUx6NFi5HK7u6esMVptN33ZwSrtBEGtO9P1csPC5vRiZglt3p
C1EFkUNRcim11Eg05mBuIR7l4nsc3JNigR5cozhIYZJKjo5r7u1C0tDEW1DG3q+Bgr9G0lEW2plF
zES49TL+bf/gpUhw9YSX8jKU7wZPvNYY/eXGE4gizSiwb47bp5x7M8CRE4bseStRNWQFw7kRJZ7w
RUvsZMB9F7BnBwLzskH/Ocm5vcuZspjsmP7p81IrvUxp2cyONljKSKMSoq2xrnvYa4dpz1WWOBz1
zsij9axvZZgAuWk8Q6FahTSAYFp6LzaKo8SYaR8cd7uWwU1DEuk09YwuyJa+xyM7+UHPVgxaDpx/
iBquS1IFBKg+ys0KlIF75p8bT0v76DlwyCDGN9RtTGIon6lDSWvS1iu7VZltnkprikbrXWJqVfIF
Y8KQSUTjjzC9ZY6gvQz9exO4YQHuMmHJSipJNLgbqmI7Z0TqR/7fIUV9mo3zkO9GneetM/DgDZ9J
Q4vdCkBQBwc3+g9DWts+sVxBzevla/46UCJRzfdwbWGuAyxNgmSDP5ZfV9fIgNepeZ1ZLRyyOeHt
hG0saxcbmMkASyiN/Ndgor4s9AtdNSDaqutt9r9Sg6iC/FC0f0/lIyoCO3kWLAKIyNt+2lShjNzz
dEEHl3cV7mU15OgnsQ9JS+4U7cbzPBqv0PcRXAst3p0UeSe3HxhFSWZqUHqiB/0PNpl4jEq8CMZM
T5umdYocwSTKrGujag31HH76X3naR9cytCB2ZrA++f0izRnhg0mWUYMSsHNU8tCmn2S2zgacY8R+
Y85Gr+6yY7MjUPgm9WD/wY7p+20KLVjAmts3RQYIn8fMSuXj9AHPTpDbi8NLQ3D3k4jMbzI3Iorx
VXGvTIgeOUOkzGet6yQ4TJGGFVdPBLVBgnuVpxSjk55LAKmKahNF1Kal9MHKsoRYTzZd/bKFilaP
Nz94GDuvdQYfhihHAGQ8AejbfpuoYM/B86TIxPaMOzb6g8rE0NUWKYxjuvc3N9kEJ0QwhXuBonut
6NLYtTCL5dF9om13yD6WirHxGz6T3Ad3XemsFiS80c8rjBBbbwCFwyQa1ey8omZbVFsA3/+cuUkC
3WYCXcG7aCnxqwfHMNLSV8eplCgNrJefGKQuutOpo0+arjEJbgiQ/9iFvXiWTXrxAtKZXlPzAkIc
21IXlIz6M2xPgJRLkXgi4rMOO9Upw6TrbYDZAVraDAcIfmUhCc+50scun3tUY89dhBC7TNLDbo8C
ukehuF8yhkeWK1pj4EXNLzSFCBOc9j1jlzwSpV9ALYtZh9ZHYfWzRSineJwXFnivHUqA29wuSfGt
33IuWCsgieomtom4uf4mwmZeWieEuNLdvFRWUaCHS+IbghcpKG7tZJ4w4NCSfYU3VpevmYtPbERQ
A/DPW51+HwYbSwkokHD/kTHhGnkglCceYpZFv/TzhK3JHxe8Ch23SEprKoFwQFih7bZ8o7iLPX6q
qzbJ23mfBEUgKGCai7g9BnHdwHTF0ZZEP3mwKCjfwphB3pLtlgbqAtO0J7qpM+PsIHpHy/eU45xJ
DXNb5josLg5B8VO+MnplByp27wewn4KiHt/h0CoKfpLXG077ntNWfPHqopxGTWNZYco1ZHoeehf/
1WL5gr1h8uikO931+9Z+aakrJrsJwS7xKOWt6lAmR9BxGm2D0gaqPCy0BWRp3Tlb+Y53loe++qkn
VPf12z2hvK1IyjmgSarH98yFwyJoVumZ4SzftDbNDuS+7CCm8T/mAzK4PaP+7Vxge+L+o/Z4DBXo
NAbVpui4trdRz8WBl2gBDEogHl+WCbs0mHz92k5sz8von5k7XObGYRaJnqGxpKHDYjX9WYNUpyOo
t1WVC3va492C6bB4g34uk+CB0GnhKNPBMiVU4Zx7sbfODug1P5Nuj0u1fMGzwEVjYg7afbpV4viz
OYxC8SOAkyWcK6DWJLikpXtKlLXA4/omL5SktgkZnEFuSRzfWRmkYfjwnoO+obJ8Nz2LHGsWpyT7
BuuMIgoEgYMWr7EFtykWEaVGJE/8SuLkeR8ck3slrtZygv0y8vIenvce2RCqognY+M2bhBOfPUvR
Qj9gtSQZv8fbiP9sYJrOZumaMNGan+S7DspLxmeAVR0gXvZu/AZnfVz7UBvN5a9m5G/0DBI4EonI
p0Zimn9IIGXw5ztWBDfBBDGTsDVk5QPHpaXxplUjkK5KEJ7fnSRzfL/oK5JSC3MMntaL9wuwqV9e
jnLi9kGL5NvzhqzIqaUpj2P+jhs1eAQJu5CRhI5oA78FgOvcz1b4F4yuaCVk9DEQCU93VVIoMqGS
JAkfnsVk9jeApZR5Rpc/+YqpLnyUM2ZacvM0/8J7VqPzTOv54Bf+IGVqmqiN0Nw4TeYpUdPfihuK
fR4h/hZ5Ya2WxwBVK396HCppF0G5+pZTKT4arImlZtpVYtkCseAct085Pl9K7Ol3kBX8YofMaLXe
+WShn+DLR09eeECtgh5xSLolkqe0iQo7miA/lsWfcasHYCmv7TGvXQqP5ntm528TEiiH6qKVzNHM
Mc0CLQzcVNizqFutitY4t8ZRmTSCfRykN4c51Sg2w7ng4HLdT3qV5C9bu/ohOSvp+Vz6ib3uPH7s
c0D5CcXRAnNzgwlhwU0NnRFrASc4jbFGO+YB1m1TERTwYNlh1tbKanAius9mA4h3gtivCFpzvEjY
zCUULGSfRpmL/8pcT76KLx5LC5DuqZUnxPdlkbJvQCXXowFvXsikSKYkGk06GuinjvtqZQU9v2rb
nLnyrl/0rARNj49w/rbbB39piRaS3dxCFiltnkWuVIuaC6yGANKI2vs0p9RF4seis2kksxCZlP7d
EKPrcxAst2zuIuw2pxTpTHtJG4udKJBmaxSp8yVERnT+Y/6DzUrA9oyTVBRiYlJfqqH89fWCDidp
q5W4n3FkTooyFWewiQ5sxWw6OQlHfOzmvRdVjDfCinwA/FBPbon0KgHCMigv7nF34j9iZdjKDOwp
VHvVWZkZbZ7z0GmOak/sTP/USfW/3n37QQryF1NlX2xEFaFh/j3/RAT2Xy9tSaDBF8Pbw/Eysz9z
0ycryd/i85Zxhv7RIAa8+/ps4FHIkL3mGhJCBSJfFS2sT0VCGrY1a8zKyUrbVao8XvnUcMMyr09E
CpHRp+sSRzMx2b23al/2y1vOBwW9tG2fguTm1OOSlKyq6c7JnYefI9cyyevMSe0IDgteWXYaw6E0
Pqz6oFk/xYWGxknBnR6TCgTJ6DFLJdujXx1xm5/ryGOt0XUJz7SQoOmCPvQ7ldHX2bryyNyl/PqM
tvl9uEGNsLYd9hzZ3fX8vPkVgKKbMcDfmVO1lPW698IG2U3X74QaFUebjAaX54RyfBkvI4VrRgyH
/lZR1B5pCfDT5188iwGJJczFVbgSigpH2Zrnk0tRl4D+Z3zr33KEqQsbJhUrQcJdwjO/s2RDA7fh
qjMRm7voMJ8NbNcTXbud7txdpMZrFwdM32ExCpiNqv23WUZ/lVWOy7z02vjQYucBsNoo97AWc+2J
Kwcp4JztBL3Ndqre0eFLnkMV5nlMQCWsCfySe9sr1gKzRDZv8KmXEFlCalUps+mutZoN0b7Njy84
68C4DhG2oLQNk712X0LUdEMStg0ZYAug0EBamYZMqrAbfse2usw2fT7aHSsHa3mX9KmtFlmNE+cg
gsKns6pLboWkoK73O+3/7R/Z9xVMkf4el8Zs0o5KPy0uT4yn3qTRUuwcXuYBnxohrpYLAEn6C3Na
n9eYsRW6J824Zsm9Xh/lVcKOzkI1uj0EEaDQdLhf1xV+6vAe1isT61vQ++9VzipKzKXfUkCcR2Se
wpOFU4Cf6UrlVtbitWhfXVbdanDmWTYhGtWPHIXcUJfIPlfNX4Mkjyx9V1LS3xKUVByAlMDORdel
Hg6OlMQJzpYHxDHgw+4/6o50vOH4WZS6VhSTVoFCDxoO7xncz3q/fQePa7kthIFMD+RtfzvKn3EV
jj6jV6WNUhHfE1waxXM2s9qT8jU4iCoJ5o7XIGfqAxrWI1R+XUKY0yyFr+DvGmEtTmcgwZdcSgRN
2C5G3C6PKUYFPtdj3fEH5RGdLrBsX1O/G4jIc+qbQeZPnNeCJvbC1yphm3TkO8p2bUJsmfPjkiCr
X0iuOzV3v8dmQRoX/PZJ6IjLl7qcNmTuCyXoftq+dC62tZRg0SQnO/50BeMjdkoHTEbZEm6/XeHB
C3cOhehAQGTF1YaSMecjMnCzE1T/hXOHOE0Wjj0i+JasKpgpfR+VXU0Cqzu43NK1861GJck9B5R3
zbkMWhD5KIiHwD0Rgof0WizOD0r7bB90CsWKeHemQ6tJyeRwGVRR2Gvctd1LMAoG66IjlY9b54YD
v7PT7AccBSGKQCHG+87grSANsWjqRTzzPREVLSR/4LiC6ChJMceTp6XLC708EZad6g73pGhq+6gt
t1w25yY4ab/gcOq3zj8KfwllycYcejWq91uxYI9M9vl+dhMH1u124LvwkpXlG+z3Vc+vWqw3zgWH
7Mh/YOlpmpwopD5GFCoNrq/0uWRwgJ2W+QQbSW/OMP61wdsr184khdyiSs3JQaLLfErJ/N/UDWgX
u5kWhK5onTaPNtOSxwD5u9G3PGbX9Ix4VHBgaOzel8fERC87kKcGj+X5xjH9Z81tIBcX4uORQ2gG
8YPErAhS13gQlNIOQeMl0fhTB9mcSDJBiox8BtT3EAueKNVNKDmGc+6A997jKP1o7D9J6fxPMaxp
r8EcHvCma2lDWOoRpjBU3w3V0dqezFMiW1a0CMoqFsDZ5CVQkCcYDzkQ+oT4TdXz4UGqCM7lKKEv
cW1K7yeTH56tGYnJrPI/VfyJrcmQtTwf+JxYbHBc2gkaO18XJBVnsMQhtrfPu/v3mEXM1cUTBzuE
2K9xCLeXElvmqywOAdWdN4KrttPBV8DX8822xkEIzJ/7GrfO0MgI67xyVlkKXj2FNaIaawr/MnIA
sNhCTURe0MZ/kiv2ZjhbhCz6n69zj10B0vSj/hXq0fDZvvIgvzprmniELrEjgQE6LHx1g2OeClaM
BESQbYZutW2ObOd0e7pP5i3zzjoR/s0djQHd2rkt0BEcHdA4q+3T/k2/YJ47gpbeo036/wMC+Kfl
98kY+0kvDAE5wZmCpdd8oeNS8072E+f8aAZ2FxdLpINQvZdrePRdnnPU9l5DK2zYW/dyzpV3frz2
8R1O1UN5i0sMVoWVvTezW9B7AcG6Yk4k8l+fhSbM/pOV97dzVjDeBThY6Jyotn897uR5gVRlZcU1
1oD+04OZng76+WZViyrtx0pRUpsn/y9wAtGnVJdC9+4jYM92ckW5gRCJsIfS/Pk+hPjG9oztorkq
qtRiAZPmzqT9sRWyEz/Vi7A+grnReXr70Yy88vC1h4jFoZNias81FL0Pzmv1kIx2POack7CDjzCc
vfsDE2WG0ZuS4dGSnwLPXUT0eix9RccGG3qus4Jszr1ZTf5aDykbcVpbk2HYZ+Qslp5JHcB/Rxcp
nf24yLqjKwakQ6g023xb1JileodUN0YOAaBC58Nq7aPISZxfT2bO6foVXhDTZ+mRUjf0njk0eLx8
GbruoEqXyjaASFdApqRxw6wmNcQ2zPwM6olaWOaJ08zNCp/LuSzOQ4oNSxrKxXiTvkSxVjNl65Ku
7nmPt6yzbvr5DZ+ZmFnzTGexyypfnIJIUZwmyllHhvUvzfzAJeSMpVVTZ4nTRac5m4h4xSe6L+o/
VDJOkTfVppY1pmtztZluPtufQjZ2AgpQ6bHIXd4OruTQjQ1PTUHfYuPIefHZD+TmL9Gs0JMDjJpI
2EZnfz9GCup3lqXaWir3yaV1S06yMSYeFmR95cvJBzLRu5gIIWBy33Jxfey018Izqu1+Hzx4GEjp
ro1pI2FkJcbSsSbHQoSQFYfVZWxWyuYdYjVOb+f8a85uChd2ZUOfPR51XIUtZ6y9bBZiLzQqdMga
7xhXE/TGXPg3ceor4TRE57M1mWJAm2p3iE5UKQrSrgL8hHOO6BsmP7Hz+aSp6Qo2ZS56BTUdqOCw
AmIDAhE7tsaLzz2nn2YmE+1kAParIgYIAe+TT44ZQXIkm0eUnAW5g12krvBGSFINPVIHew5zzPK1
Dk2zjrPvDmlwx6YNggonf8DyJuH4loRndGiuz3bTYgPcUVSYYa4NxIrObCvUdWD5ku9cW90ZwYVz
xaDuml0YYWIowfTwakNDvQEHqD1rBJc1B927XGzT0T8hM0JQ0mH4RHfgmATSr89uIqXf6jlOXhvw
+xYaJZqO5rP+oDd0vx25UZ1OVkjGZMJJf+CKOSF8GHLl20yBQHNQ3T+ZiQDAc1uUvS+tkpKRbIOw
8BGpo5oGlY8OK6PWdy9YnZAMPciX0EuN15tI40kOvLPiC3iFy3uWDF7Euwl1sYVlT9WX3jfgCLpf
l9UgL78lAn9sauQpH+hnzjqqax40Ie0cuB7tDvQDBCnJAGwiq6vV7+jwWS/NWM5Rf0rmCn0Fhztw
ik2Uv6w2ZtnZxG1Qr/nTv7RCZy8Cx9nGoYO8xZnNXAVeJx0f7TRi+6YHwWGw4+nrEFQ9hmPXJ9k8
iQJuMS/lLFqj82RmFIV0Ao3C1w6tjoFZindCna53N5Z2yuCnnoi172ofETnbDgHl5HvruY636sOl
HCb1tmaEvwFLidR5WX0h/75Gt+8+WH+ZnqNxvYbh0zYdVlEYO/CekMIEcTjG57KtRNf7SmeRFs4w
b9GfLg5EdU3R6LDYGcnTiUKDFAWAamT2t5Vq7gEdmetGDOrNawOaCJ+6HcIiIZF01xAmFtLDVCVl
7n+shU4bAkFw+qKJjkVT1LwN/uwCcTGCydqmHs8F9f2goeDQlVPPA4LS6QPt7WiFSiLTSMgIL0Tk
zIXWnLKd5PLSd26XqXR/Gx9SXdBW8h6omU5hGzobWYnMwYssZ0HUKP/mG9JteKq5W2oriCNtECq1
qCfqz66pNV7sTXeQw+pIT0T6Y3RFl4MxU2IbyySzEJyP5kyZJpN+UnQI0DbZZHCO57VVLIHVmgRD
jmgScTKy12ne2v71ohHfmM6Sfu2BZGdDP7ZNgnH3JuGimx7cCuU+m1ezJ54Ej3sgtcSCqQN1amzT
SHGi3FL3lcdN6kdNiisyT32O+wnH0LJOme910I/RjL90RMYzDVGcuyDgRklVgw2DCwokKxApNOe+
/LyRUDrYHaE/kLl/eLPBI67Mbm9KAA32WeRqNL3eAN+TtPXMmBccgaiKMpjQYfxYfVT3bwyfFpgR
OKkvb73jusuZKJ/iPyXrM2mSvXfIvAt2wn2XUdZUotIGzCKKzOmOlDUq5hkxttQ18YjgJlC8Lx21
1kRWLFltgLmQIbEyN1k+4rk/V5TCcIrxjkKc+pgkWJQezcVB25gcyubJ1+EvuHWkeyxWZ6OwNxJc
yMPBqbq/vM8vqn7e1dmM4nuHTrv5f3kwcoE+/OCNwEg0/5Do1A3PGAcXezaRh3tPmIXeEHp4g9gW
G4lcCx624VYR5CwcbdBHf08ghhKhYI3f/+Z5Jjxw8P7uYIs7770NswNg6awO5aUUyU6dxTJ1PweX
6ewaZ0CVwTDbZ5Dk73vXqzIA5loLGsXJ76uutrSJKN85VNZUe/FVIAUtR4ZuY4rqrBYlT1vndjS2
I3mRzkc4jY8qg+M1onPkzSJ7VheKEP1JtYAGFt8/KS2OcH6vr0dX1S0fcvyONv8w8kGwmBQcBGYl
2bANK7HX3JW1YyhBG23Sgy2o39Mnq5pLLg35AXo+8Z/HUmG7HqYqBRxkL+v0k/mhOboCuz3tEL3A
lQWjZTjZ+XptifVCpnM19dJbiCN8+t7ex+FRC9ashO0zV/KSexVix4IWIYCKFFsl9W1v8Lp+qL2f
UNUvgeKkaA00b6MMZzBTfpsrzgvVB0pqWB3uA22k4S3/xhcoSzZoDhodmjgck8bKwzdNknMnmu4S
3Vlev9mfyRU2KGhxV75wtVJ5Op0kZ2tYpq+KDoZbdpjl2lenWaNdOfsI375XGV+cUkoJJ3KFokiB
DcxbhauWAY1E+gOTbg4cYaf2KNB+bfNHzitW9Q+Z3baWX7iK3rGRKg4rnGeljsNt6n2M5ozzeqQE
2kaYHzAh6cNmH8UWkxUXGLT0TNL/h9D8cFge814vrzAcGMLmHsMdlMBRtbntE90Xkv204gWvwTX/
935zsgJ6CBuZiK84C2EOHKXDqMPI3Ld01+m+iWk0UCE7M/Ch/GVFCe1THr86khOQdFX3MVV6sMox
3tr8JaE6+8zQlo6ggl/t4yp/tr+lubQDU0/EGxFs4koG8bmkeM0gkLBReab0qx+8yJThK9PRbMkZ
0GKigyQF/PflLqhP7s0aLLjZjhuYnBAQPQnOoW7/xGAplgFX27LumhWQThOwtVWsY7JlFy8IT+2H
+PnxpLJA5EY8eBSzscVBodlBsl1KE18t7D8ifVrxZLJJioC6O4mJWfwL4u0ZKx5ZzR+CLxjjd0/Y
eFtpdIOmI42dtZKtu+kIRSKoz/OF0t/ddpLDk+AQGlA9aPc/o164J60c2CDbdKo57FQW3WdCvZ2K
canEx2fMAJ+FUEodt61j6OZhObH9Bg6BsGztb4UgWjmpFLJ7ZQbmIytu5rfLH3GexddhQlsGYJom
JAcwZicGKMvJglo7pXSaUoZ7TRbtuhYcDreeWDvEpmEF9aB/o5Njcba+v8SzOhfrPnCK9Y188NNU
4uH4HaDNr5AVyGVrQS8pvP1oiWRKxi1Httb1x0uIvxi4Eku5tIjWssFZdzTrcQqBELPQGPAC8wKF
1H/istFWsSaSwJ/gtSm+NvD6qb8xQkg9HMDTBfeGkE31VABUA0PEWUCbmxszGieso8Z8W6yNOir2
9EFU3LDHakUqIPrDfPELbQn10DtrO/uDEw1NnHUc+3hDRiT3WPWRI23PQDfsttbP9vm/xL1KaZ5y
RjNmr9ZqBhAf2Qvrn9+aqWqbVOnd2Xzc1nCK8QRBdQTvW6CONZL/2XAa93N7tuDno2iRGEd80m5m
GEf7rC/jF9royJENVHuJhu7S4VgDldFIR3um/wxIxJnJVJuy4ZfqDZIyMi1co4guv5QWLQpz7xrF
uxtw2eQVRHjFiIvckmE1JtyOYvbQqH3kBhNr1YhnzK/9U8Yjmy6s8PQuT/o0Xf9txBs0B+oHNOCG
UHHYHZDWgQy8g8tuSntVAz2dF9hgeB28Oj/0tS/Vc3IAn5EG91wNo/d6J2w9kpP3HLJzba5YwuM+
JNjTQd/gaQLLeR3oMT+YHnyRwmOv4ejxcWTBd3NLRL4RBXROEaIvgRwhZkWEO1phno9Vr4wKTzuv
lI9JLhuHYHohbs3BcSGBrTmsLr2vMSLbrcH27gD4+OY76QU6peQLwPtOqKYNWr314oCEbCveUs95
h34dc60kXbjlTOivcODy341trnh2Q4by/mUWv2kPBWVeLXDxpyp06CAA3y9HtEed5I4pAlbBB418
ZRnNkffdxKb43RFrX5J4FRL2KiqiouW+Z1l12Xo+zndxkXGJoQQCjNjewepdfjH78+vUaElC1lxU
edCYJyYhpzXZI6xcyuBsIRdxoKyL0VDcKOHZHext+F9rNWsVvYoXTM7IHq9OxpTdG5yXhqGa9ZOD
kifHPv0g/eTZkhQXvlLOlcLsowkYrcMgAoKpZSUluTDfLx5E0dSjP26VV8P3wunFEP3MNeemHgQY
9OQ8BOkax1cKD/jPX87IVHlaYIe2ng8fax4zx+8iYZ66jKTjrKAE2meHyRVIvR1H5puhSyoQfVJb
rkve2GU3fg58n7IU7Z046JFYBAP9lMVrIqUQQjQB3UGheRCUVQB/9tz3Fmxy0vbtgH3kML53yyU4
vYU0c7l+tFxCMb2MDleWXMHVDc4C4zVxzOoXglLLcQeuGh8LMqw1LhgD/P+YkFdfqH0CL2ZW784c
hk8R4hvozO3mbQ+qd1PeMTzs9gZhG/t082OiL0MudPRf+ffqCqnp2pE8iQsIQSp9YpV+Uvrb8z/+
GupXpzPf20U6WuuSuWhSnJL+s9lVsoRQSLGlfYd5buZLnzAbClAvM2G7irChNlkprbqedpTKi6Rw
JKMduovxZU9BEkme6xpzLwCspcNMMVzIxcEoeKSDF+3EPllHiKgKPjUJPGYr0X1usCXbN5PEdN4r
2Fdp/DrW/uVPRqTFUkfk8RyYrGyVeGjNxh6hNaWfpj8vcmYOt3CRoZiw25rWGT4RPmrJswdRXF1Q
5UHb17biT69zOvNnP0FOI2qp3L5JzvzGXxDiPqEtjq2qM9CDeQ3neDpYz3JsJx4tfbXqoMGqDCU0
2PuLUfw237ZDqEG7rbg5ctK5F+evtN+tBIXDzQV5OIymS7MKmoQYiCQDPC6k0oj9d8QeArrrHyxZ
pHPN1wSmHDBUN1KEfFwSf4fv9CFPooddGNImC7c+0+UBs4qEpTFeGFA63ad7q62XDJKlKX5cwfJm
eEFsI7C2YJLiIahXr4bYlgzgZ74g/Sa923Rx8Wo2OMU368zFovYj3ngnRn3U8DX1/sVQ3Sb5QsP+
vuTsdJCMN/9i2G4cP5uhxxzkKVNRUPCi2CMc1TAqnmsgE0zqCS3zrvrByFmhnAUMJK2XepkIH1JS
YQgmCSrJeX0MEnXYawkKuFp1WPmIiET5ZEIodDCvlGi1M9zd4nT89/LxJuZ5KQlV2EyOxP6FagVx
S/zj508VC11rXX0NERgcnkno3cSnERSPwb6giNxZ3sRiT4IuZ039xIDMSdHrVvXNqqPBxoEiHi4p
Ef2lO2fHWUQ2blzpTV0/++SyDHihNah5CYB8kbzHdkej3Zr1sNwo+cPDOGkqj9TIrEUwgoTbVgOW
JqYLGaJgpf/uBBKJwSK+H+UJK1cTaVRsfeDxRb/nFeYA8AtNdMh/5YeyPlQNkYeHVb9UXNT40It5
XvFoDLKLJPFI4l3dVoYmEuWVQQLLNrretx6e2zaFhJNnnaTyXeZ0Zoqb19Dq+zac3QG8t/HWQxv9
anhb2OSS3AV71YFUf81DvxoZuScKR7ywpw50rkN8YXLht/2YgDXkmrT4tuXCevtFCnZIgZOLSoIO
8FVf471jfYb6ffeC5ZBpIx7IyIIep2xJgipWAa/i6yQj1egTmYvo72h5jST1Kd3qBEJFwF6XTQAT
dyEuHQBC1n3Hn9BQqjB/AwTr0jK6i0w0cnZTy7eXI1WGXkoMQuZuMxcvqhKRCfovwJAG5Iumm6oT
NmFyq8YrYTB3kCBcyPak1gGFRphAIqz5tJ6j+aRRsGh4EKptb20jSzExciJs8VY0a9XIvB5i7mSO
cVnkUcLKKKUWh0BQW9Km56zwUoH8/55WDs2IBsaLbLY+WDommYiWXt/a50chfxw5wDOXmyJEKL8u
tZrrHpcBq+pJT5VWCP9KmaYiLoCwcExYnE055/OphJ9xC7wsBn8zYcKXTOnBmf8tJYoc76MN+r0q
LOprNpvIHkByRIPY2izForNwAJ2I1mUdnFdbVtbI+wGQFrgPPOAr1Ir6hCXzO4x0iokQKoGXI4r8
a7Lc+5gVxlytayei+NK123mGmWNL24yi2HaGJRhlsqrSzDC8cnNfz3ndLnsgR/0zajTgz3WBk9nZ
utetxgq+6rzHiuECTvWJrYmo90WgLFcyOOLnmL+ycvlFTQox7szbbHzfXNeps3JdeErN0jP0LlJ3
IBQbScfN8pga/XBJCSyWGMe7UHgLR7ppb3Dl/k5Z9UAbwUbjavunvU+8bvazTbSH1iHsjasdLeEv
ruACVDr5xd0d1siK8MKGagkgSkEjgZCVFy//josDZo6MptcHLK6+udXjBpD8g0NJDORsoW7vR4WV
lEYTWWUxFOp4rc8yZ8oJALnqPdJoiT1dY6ogQnUK/4UYcQ7ECmWa/Yg8gUpQHfh02lUzcVSlrmbC
zwdKMUkargBPJ0z/wx35OXDxXQafCnZAfvhygrYXIerNpYsZyU9pZe9waPO7XXLMvicotK2ss5TO
UUUkWlU+d6hi0gQO5ViYMfw2fq86Nd4OJc2IT9+dKuimxV5JkBJrEWtKr2OunR+PNrEL+fO55ER1
/iVYRfkYgIquNMH/LAkOx6MGKEqWymXQCFva2mRNRMyXZD+BlglJr9acykqUr+gus5g/PYpaZLm+
OMV/Ly63+0MWuh9xvC9AiJwdHUOmk8QR5kf19ZKyXblDJMR6j0cYAgGCoxRO8Ps3vKt5eT6+QPP1
tU/5OvHCAxWLjYMSkA34kpE5r/rY6kya+QzQEHuiD+0AFv0tiA3khbCGJxWEK8mvaChg1XIHbeRk
NNhe3nV7LRS75PQTsZjnTaLrJQc1SHUQZcxE4J3MX0nPOx6Ypt9Mcj6uf95yoteAmAdOWkUjI2iW
8O1cFwwD+MmkISIucGUnk8Lc3tonG7JXnGvhJtgczkoNVdAwAfG8U2i3s9yrt/WTSvJGViNfOuF5
rYchK4dLCDb9FOjtdiL1F64xLZu83I4ZktRQWrSdAx3IAQe5oZ87PdfyES/I7hc456V9325NCIac
tolIbsNsR5Z5VC3sgKYCBQa3kzokf5EiBiuobIOeTzMTbJec6nVyXJ2+c0MHKYF1To22xwwzxoYN
RYBuvTHNPiOp0k5WN2HkxiRrW9cTNg7/ozUpOAc+bosdvOZqXW4TTPCs4wiEs3QLFajxWKAu9d+V
iiWwGGMYh6UjHH5HEKasjEkdVA5JQn/otd4er5swd17iyjOMy8Aoj5sYvtD0YZYnxQdiRIsrZsMt
KgunDWzE/m4F4gsAG/P3heMVBHeWuvr6vPh7x4oftKLZQpECMdXc3AMScqm4YguutSqVeuvHyN4M
gKo+WfU5OEBL1VhPu1T5QmGjWxaM1MY4qJGWYrVLkLyoX0sYLes1Q7d6ingc3HT8UFoRfTb4A7nJ
YP7SBhNoIbQOtp64Ivo5bOFaFD3rKB3llhLpTamIKTjosqNeim6F9XMR7YsKT8S3aXZnkKy0BZ5j
x+a426W1bBp0CEd6jt9JZDW3ikJlclDfNOE06tIMh8Hp5KkrdGt3/Yph84OLdx1zkV1gOBir4jaS
IwS+DTwhQ/LzyBHlo7Dl1OfRzPkJDVKbM2SNa8zmlnRqdqeueSeI9WnZ4PKkyR8u1EgJlihYFmJP
vp0CH6vvN8qRoDhHnlz0i13DuZ6GLtqxEaU0uZSHnpvmN3nWdXTylvPa3/ougu1JShns9xV+r9AD
vf+3u9ND39TrXNt0WnipUm6w5Ij0d68VI1cNGvOw/SWVbCb5xS7vt2h51i8SGM0w6XbvCTNtrmvh
OB3LwJzEGtGaio113VWgKrt0fd+fVe3F9MaLU8883cdw5MRtulSDA//Fq+gcVc95tWrRnZvNjBHR
3eTPDw7BdOlQwJrWjzT4fcr4Yhe8KpQW5UjRwmRGyXenmN92O+Sxxn+5Z8Pu4a0MEgYsabbGVV9/
BiUKj8qPIXQ7jwNIv3Q5tcsuJghT2tOaoMT6RS99ViXKR7pTjZ1rDNkHgPtf6ue2yEipWxM4AW9K
HS5F4EpG2GYTLgeDvv1j/mPacFWgbN8dgLtXaX+wtWLzCVKJS87h7Hqv3DjkydY+h4te4R9m0ykX
5R80TQYJ0tmq4ZsWeoPyUDAZZRftT8Y7djKm3Jl7fKrdz9bTBDZmUNXotGaVxzpR5ssQj4YF6+Sw
DbcqSpvKI786sLK1e4OPl9a2wYfHKSQPA0McKPZ9d9f3LRLiFBEkMWIryVzL7HP9orPCBG5YSSth
DEbb7epLnULiOSJdHmnTCY7C8Px/UZUGnt0fne9lDHfVWLZcxvAhcxslLJYXUiLIO4VZ8vrVRxaP
l46xi1ptsDAc366grUMUj2nlFokW5oyNjNQ62LmSUBkcpkOJaOCghyb7ZUH5rprgFlEVZGLx8NlI
R1YpUEsebYcrMjhteyhLNSs1hSQKzKgKQtgZ57OSzL7Up+ESM7hB5Q14lWzXjvtY0mqqYauo7ixZ
X+v4d15cKY/xxJ3kPqkvhdU6XUV/JnFBW+5LqP9NoByEZmRulCMazkTDGQHZMZ2vnP8mB19hp7r4
BYM51TjYCoqH7OL49acTgIA3Zfvpp1CkS2NQSBauL2uSgkz4JUAd+iNrkPMvgMZS0d7K8pCtNFnX
UD7ENtmQTeK3Z4bwePMiCIpFu1Xp18HDTnwpg+hTXMPSs2qDjeGeP9z8VNPgEosF4GHaZVrbHi9f
iij357gO5fLBcIqP9iOEQjJFpG28oFMfqMfco6VVibpmHW98/mG180InSg1Ri5BXhJd9hC0/dJVm
i7Qqz2FtuMS3bVpwn2Mjxah244mZJaAhs/X9uYM19+iqIM0BgpqdA+zREM/Jnrzp4aykyxbeHVa4
+PG5294HYgM8fGqwd/uhsEoKdCCCtDkSZqTZM+JjvoWrj2zdsAvepu/XC6f023LfxeUcZwK8Tta7
br8Hc36up2dgREc/oatZ+fm7uKsNXZekLOA64vkF5/EC6Jk8VqQxKPDqdrTaWJOez+71CoOxg85P
x0pcB1DNdcS9ChRMsQ/UUNUff0HzNHIF+Hw00GX3xtS2VuUMVsf0vovfaL2fSe81mPZzl/olGmXH
fv96yMRxYu2Cr56Yggejkod5X2wAk7umFnVUUeeUYC5L/ZK5tx+BvO17n7WChEf9oyzLnZAjEEWC
jeYjuKO3QjjOVkbvYv1dPjhVgheLW8n81EQWlqDYrn79Y3B77On1IrLWnbRmdnn6+MJtWDFrfkyp
3+yk9JfLieAbeSoFbVUmSBcU4gVkhyaizW2EvRNwwTLpDclBJOY7OOnXeO+fMGZHMbuxqpsXoN33
g2Xi9YU8bJWAUgl8wp5rFcJjImjS52AZAMN/7WmwtUI5oG+mfwuBOqfbqXauvvOuey9Zfo8Bxuvr
sKgvMyz3hDmEePwU2EtZ/2amdMhJeEJekcHimgvZyvXghJtQXu6Z9JeVfsLN8G6YjHBQ6GsAssAK
3+WrD999kCgEQnaYZAOP+72rBetV1I1HYP/9OJIdgqdxjyjPOOuk8MXWIQu25lvqLcTdGxJaKLfL
9X3OzEHNtBLeZC/3mnWeCVb5Qv3Nd7qBRS6DXNErhgEtxAWcS8UA8gZ2H2n9CaIr1gO27HyTooo3
dwCTwGFSY4D8Mcq1B+hTvNckpAEg91FI1m0+C/5AgJ1CA+rcqGSU67j9OeknJrDn1npjU/4XlK7S
zhdmaXQhpHz/XV4gbcVzqu4DBNBr52ATmKija8kWEd4iPsz7OoJQxzeQ5lwpV5GtYAwbmcfrRiRq
O2K0RMEBYt6+kAs442jUkMgwJXQubfLjrzeliGw/znALUpbsGYbrPy23YckswTyw4bZFEYK2adTV
YZ0XMkOLtMrxmdWwRgLnAMk2myIzOGRL3jMS7eWo2x4q0LKQ7D8wWrq05PE5e3HXxcPBEY0HXSfr
dgBZ9lyOYbRz7SoYywzBVpqRMbElelNf47suYqh0r+B8pXuVx2DXSDvYiCqXh/dhCYu2AhR8PlQo
hYciFXr2mETV3TcbojQBsyOC7TNZ/FE2LwqcHHAK+x0FX1PBefM6KVTWaJ/OSb8lokp01Tc38e2X
FWQ2PIy9T3G1jFa91xqcjuWosArNi/BTRVYjpWa5T2TC5XC/+5bi0MxViD+OI1jbeb5aXlcLoplB
BS8hrNOVx6Sl2/MCE/dCiqoMIvGgKifPYg16QWnBVtJ5+hAApTJiOM1FwfOwsxSbo8YTBeU8Gyv3
KIYvkwUVqwCJimxpH2+E5N6IP5M1lf95LlYRSoMPU7wdUEVt82NwQ1eTTiQ5X55z/BCtyHOYTiZa
3eb46AUXRTN+8MIgthfvvEB1SKlgUAF4x9Rg3kZLAKKAmFfm6UUmM+HAE5LXkCKgTj+lGcqoyK6c
+qtW240lX5Y21mRzilVo1GDJrC8/aWKcYVIQ7x+unwYpEITFG2coVrDRcWmbXg1GMnOLf+NLBw1N
elWuVEIuA7WoeQ25ymEPT/azHcGSD7M90oFGYNOodDIB/1K55iOwrv6TjlPJWRlbRq69Md3Ad5yV
9WZVeMZpU7RWjI7o/ZLRJMF42u4rO9fuqdZ1jDnH/pt7+chJz0l5CyLW/BLHmCBom5d1GGn2Mbno
aazTeaqjFvJh6yH4ezzi2h0QdAWaLD8HRYy/ZJtmRPs2JKnymtb9NKK1aQTPvs6yDVkq3RsLrChh
KNJtcl7ybWjjj1NphyQ+nntlJc8yI+1pScY0BANFHNgKyoPg4uFzysFTglpuIAZJK6wtjfPqXsdK
Edll8zvWhNNRCs55N2BrKgOCbnWcAfEkQDZ9qap8Ju3Ns7PUnJKbzE1lUdwq5KPkc/zxp5gvL4T6
r1inKEmI9tb+zp2HAVJ6ht7ye6ZW+OqCCO8a6ZV+4Nt/6BXh3noRW5dazljgJFZrkFH0pwelQxGU
gGOmW8fYiDPCry9Ff2dtd8YO43AOfV3HtMOFWSbuUpJ4KBedfm98OFijXQ2Xi6Jp9x72zXh1xInh
noNq5YFDVTa2XBQOjWqDfnYFkUO0tFkzdYy0WRV+O1LlLUAuCMkveneuaCOwicfxsA7KfgH6YioF
jn1p282R9HMTuBPsVM9CRnPUkbNTmNqCflGRSenB3gNVLR/NrJz4lv/AiVBY3xmjkygbT1fjQ7C4
KTMRKWapBthXY1dZpcSqOyrNEinue3GwsXyWioDJPmiLd09xhtnHISqX1+SBxM4k1ff/BB/pDNmO
Ln4KIY8Ik1tsaWWChwuNHC29YxV4V7hBGUGCPGoQ/d0/PhmyORqQdwM4RXcWDyx2yjkLo1ADyTaO
KQQ9N2FP71aoqvXeETRiG8RSxufvjkz7w7cjn6x5c/50uU3o36jbbQsSpSEX4NlGJ8fcclKoOA38
UeGHZxKg1ttJcOdwLH2w+QoZ0oKJFvQMsvnt8dyjS9ro5QQaL94oSHzz76zOq8Hatr9ZRP84XGEx
vDnULi/4Cf9X3uhUmu95GH7u+yDJG5yHAyxtDXmhc9Sck9VhS5I9h1pOVoeWogd1nM93vtImkYpZ
FCz6mb1KK4msK5BgR/4rjaXqExiKy8cTWkO+SlgdeZ8slHSgbG0hYndtvuiB/L2pUdhwOrJpnvlp
784q8ciV3j6T+6GYqYIxRLiIUgwQ5GyvM6TRnU81CGBMC+Sf0N1PO50HmJRIIPZkzUoOmUR3nnyn
u5OvAcg8EN6iooAbUaHRNlRlHEXCfls4CaBm/FC/CJstrKO2BzXe+XFUKyBTjyD6nLIDZOrTBp97
akBIx2cwv+q7Giot5RWoZbVBRX5GKv1sKPjcAjDIn6zG8DgDf4DiMNQZ5hdLI+ZUP/T3uHyeLAg0
ww9S1fc7gDekMf515czZGBFsRzF3o7Ckn3P/DmoAVbd237PqfUGFxzvwwrmKfJvNlE1rAdr2KoD2
sfAolIEHD7D/p4p1YhisfMxZ+Zn6nxp0KFVSvSikSRuUcLMbSVJoUUNzcDHIJGbAyCXRvo7vRXgH
DyIUvVyJAWfN5+AR6xIee5zB3GOB6eIVqyO4Ty9TI75bpVggLHNV8Tiw4MasUnhl4NghMOYfsHLc
QnG1ycL+I3msrdsQihXaUTU+Sl0hGpGUsXWkw+c8TIYb2wd+8cIy1zb1edFrFWXQb1ssfQqXfuu/
O+Ooi5eT/hNMJjTmAXE+71onfJEpitL3ddu216BVC/uZTampIMHi4I8Nrmurg1XYhKimjX2mAgs5
LQ0IO0aLZYx52NhdHk6FXsOlwxCOrwZGMQsU54jWy5RxVqBH39kapovXfOnMG1tqT41IIoX5Jy3W
/qJGhsWcf3+FD7Xze4i4UdyLDW2BaNBHLN7hl0thUbaVe5leoRXQlFi2VFOAVkHl9Uzm3x3sDgIz
1Jnm+9TNN/lbrZLhxITijU66I4lOgtW7yG0Zvx8DsnDsUa20Df+NZfNqPXJaN8HKl1w8Z2UM4PpL
uVBduCMyGLqYwp7teHXlw0nxQc2Rd94L//sIKrZPA/c3ikWqCX1PKyS7HmLtdTKuGlQWk6HrwspM
pr8Dhk2YU3eY3da/xHcpbfukIRHKPjHPMI4wer/NDpoZqAw6u7ND6qROIsaYqOYwcyhjoYSH2rys
2KEQz0HTpK2OhM+vcJXHIq0Lmpnc5+yVlls++va3M46ja1r9LckjY4RJMy/MKQUksIZCOXTOlkLX
pe+DXU88CESHACVg8ljBJpBMnxdTkkK7KJJ+7AXszmZDx883U2UuL683PCg3IFYdkKHW52KVj925
upMx/af/VdZU8LGKPLCgqBQJWrx57+Bo8sR5FAyaX2KGuvU9u+2U07UeV9EhyJggnn4y+AyhTLRN
m5ADcHJkJeBmzWvu5N4/trH1H2vb0mbeVf9MOK+C9brFyR2bpHyPl6FoiDI9fggCYAFaxE61PwKe
e0zGHQuYCI//pUs+HSw7EAmDGnGkqd7/01b/QvZRx/KYZTuJ+65SsB9v1j5p5YDdEshfF87fcLA9
4xmVeGEPvhJRTlCGsh2wKXNoLUEyLhbj3MlzlepfrElWiWJ73cwWzWki1RMqxD2BwauxTc4LXIT4
TGHE5DOA6wD7+jLD0BLCxj1Qsr2xeZTVi5p1nWn+UjdEk5fuwvC84KR0F+4IXAsn9wDazvIh5alX
AanqyG1go52Qa9XAPSyFAo5l9rrIEaVUuix6dpgjA5LQ/vmoQVTIjhwAXG2QygYQXpBPg7GJ4aUr
exQbMVlPBPCsIZ32eRu+0IMJ0vD1X4MAc18ixqRXgXBCHMQH/0a5hbw3ZTAHYDNe+XlOz8sYdlkm
hxqBUmyKgTRs07CvBJPuXGt8KqplpJxcmX5j97+/KR4SbkmcchBSota5yFHoaEZSRXsyvcjxq02p
niA0tqKxo1tdtCe6PFl1YyF6f7ku2Nmufnez//M7xUNOLO0YWwqtlBW2EmAziF5gJiXVLimteIeG
VXTn1C1LYWjoY+Brv9/W8vQZNhoePBmNV5QCvDzmZ7xzpDjiTXzZb9B5URAR3vgsPObY++IlPklR
4agF6SooxKFJWcPC65OBXoKH92hyIyppl4UseocbZfJlGDDic5v7cE9FWcqPZ++YigwDqpxx0l0M
TgnTNbyUogZbaFSFAFRNMbIMMTcee+apKY7bYnTbK36MLGmtqkdonvdbALXvWmotJ99HEorf2Ymc
Ldmpx9eVLu+IFtTqmy1RWuFa9i3V4+vmvBljR79qYroA81MpMyV966wcXvGfNfi0KyO2SYOwJZWo
gVXq8xmyx0K2SYCD30pZr9FFvH6Y4mW9WNiKd4fkwZTLdFq0PCHU3qkdm5T/JICkmjsmmSKDfyEE
wC4VY5ABx9zgsjM7QT7fC0ooLUBHrsCaWY/3MpUMX16rxgE32JqqRICDTTssM8Bc5wZ5HNVWG4vJ
4G0lqHMX08b2nzI1Rvh5OJLM27efrZoZwE/5CvugoFEimDWmtgSVwt40CMgJuU2a2f0m8yWigRDZ
tP8Fqayg4FM5BtGcsIN1hPUf7pOwJfAoCMaJz0AAhYSj1JFhesTA6X9x5CqJ6Xa0UZpfQIRzKsMO
GhFcO2xDI3sR9cseFx5IliJXTAG9zb3oui5e2218p+dWix/zHvV6oMGMZBElnJyrYuFpiQJeWfUl
rGB98e9dfcb8aj9oWBB2nPS5+djBepHHQ7orFx0xZ3q5zKktJUQ2+ReiNnQwcF+QSUXFyANtGGoM
oKZSfz2WDpne7w86/E9xKWSVsQQeGO9N9mLJsMEPPgRkbiRndEk0uqJN9SJY9Q+bSmrlZ/wexDdE
HNd4fM3EAeHls0bpHGsK0Kxd5yiqmeumuPj3a8UWUWjIoCt5GWZWRjr6MmhZOuLXOyXCvTWhxnS+
goqYaaQlj/VYFGeARVGLiHH2hQZNO5jc4Xr6DUTwM5eZaCutjeae9d2c0XLnGKn98jhcgUvPHfvX
oFLrHtTP39S3q8mOTT5tGI6voc3dCkEmBAYPHdAnoiRhTNUOL5QY5ps0PQseDeql2Tyf4p/8hz9D
SDXfolfBYdDr12l581+WL7aTxepG+Ee0Ep2ZZ4H6sl9HYM125oXEqfYmnJE9AJtupydiJaYqh0GU
5czyXKfqwLIjUDEcSw6RyZBj10Kdj44pL0PkUHYSc5P9Sh8OAUC1I5jTa1OJMUJ3b0+wiyVmRvMm
Ez2WSFnNLWU0IvkbhmxhLQBSivB5mXSidUBlYtSK7hhCZmChlM9UehBAT7dtlOGy8i+nPxtfaGSr
pDxZleZsekCiPNqRxQhHvKMwZljOBXQfXj7YwnR9p8Y3ZtXxKNYk9yX4qdGf4yawEFAB4v14hv4a
62HsDIIN4Eqeu9YnS7PGW6T0ORwdkCLoFG3Hw1sY4lRRwI83WEZTqA1+0vRH/EgbjtqJlv3ZuPrd
ZHuaCiU/q2iJmTMyMheNEzScMauR63ntLMHLhNdd0ojEVzCpg+dSCBiwJKuawPh0YDHAb6mMDw9S
wKiraTBeZrWdvCLEH6GLN1UIRWCGJ2hDX68D5TE5UopxuH2sAmSDeDF516879cpRB+pEFaTVkZV7
YgLtt/vlDoZdHhH7EEN8+hLc9W9waUHokp8H707c8WjLF01gsmLBs5ngitIATFZcP1XsihgQUwkU
ocvjDqtYBhlbLWTHgTbrh6amdoFl+CCtRi5Dru8qglD4VisBAgTKKAGmTk6XP/I8jDDXlnZFU5nI
GWqkzygWMicFn5Xfu4IAZ4i0OileOuCzidqVtAetctISrVHBGzJb57fsLt2n7WomXuUGQHEhz5Dp
Cqw2hTjZXMp46oL9ul2LUCW4l55Aebquz9PGrRLqJdgsFKaeGxGuNZxK2dx7/1nY+VXpcnKN1bGD
nuo/x/XbJbzB13dZlj0FUJnuMew6eq2nhRgTSD4pcR729AynbyvCvvhTF959GxwLbo+yeqGcuQF6
IHkRe3TJlcF0tZeIj9TSL4tuPwnKdJ2khc/RCXfKUNcoFNQpHUg/TGBopQ+xU2S03lYDLLsucRV3
alh+dLY7H0cM1VV97sNzF2ia0Jn0IhqsCrs0jANbGNrr/N/+vzTvBiNQR29DUcYZ7iMqutoydJ+e
BDQZrMefUr7bDgPNJYRcksf08wjn1OBOjNuZ8u8AmrabDUqpXj0w2fYUp9X2FVp+8pRfLFv+yVZV
AE+7PdVne+ysQZIf+tsuezbuNxwpiotlemF97PwVzCq7MudyQgIOi9JeoT5NR+zppzOqXy5LjQEc
BrAljOT55YqvvxM3xTjvTyNvCiN2XOyzoG3SABIzsopo6HU1lFtKd4ykmAGge1NEQj4P10amCam4
9vYcVWx7w0cipcNtF8ii/L0CCghrk7N9+asC3pdCgAtkVzBFo2IPeHNNGMzVYyBUgf3J3imfbvbN
qzq6zvOdvAipatTkiGGppUPvUvidGP9BSPiYagkF8tAZAPsinPoOkFATFzwtT/4U019ZH7NkbrkM
HZ0CWswgvjCkLboRI9W0a7wDg93FVQxK+KdgZyqHagmkMjYKaOD0y/DLA43UORUR4W5gRh/txyLP
MPo0o4r0B6gqjz/L2PxduJfwvDTKxIi6UAvGUSA1eRcCVauhLRYp3mYRmj2BRW4sgAVSw4hjb5yk
dORMXCUivbk/EP+ZRl1kau+hBW9DlIjt+DMbUjZUepKeKlpeT5IF9URkeEdtmUun3pyaWSfqK6Fc
6P7h8AzIYtX4V2Jjhka5sUWNmCvIt3GRSxkViv8mj1YtVgZP7MS7/9CUh+/Vg53jtS1xkjud1+Wr
E1NXpxXrEkCRpqShb/rmbjqLU6ruPVvvZBpidnYPRXOOkOKBM96RawaokElTe6RrScXeM3q10phw
kPvbz2kn6VDEAPO9X56SZWe9zSuD094vYXRClPI21mAHzt/8Cs4WoErbdiWWmFAVMpSLwTXAeE++
CbUOGm7JdwoYcNVlxq1FrRdRYBCrxWdUc/b8LRNt7QtKG0AbkvkidhKGMJ0Av4g8I6ta9F2hy3BA
SpRHoAPEulyNt5RzBkheF6SoZj1gXnZVIRntwrkH4ARWSatBvNgAjAO+NbN6nXOWXsm/jofJXBuD
gCULc8M+5Bsm8W8NdJUj+b1ouLCRERgnlu9KrzXQzumpRCURTrjn0kZInvIv5ElMWQR9XxpfUJ19
y8+9sHd16X9HtCjqUOFCPfTimbKkSDTiNNLK1O/q/gPXkoyQax5zvlbtKu0q7hkb0r+QdTo50d3D
qhd3KmaLDTo2vhDMKSeinENXFUOMlzby9D50hfquEiccyMNcpZcGDO/AAEaQ8zcVu7DLRI72sgKd
0D5acSdIo0ctNCnwtAsHdkfICJh/C4i91lOml8QbT1ZM3h8usDnhqLz6xdVqoE+A2pPNNOMLVNJH
NQK0lbzUmWfJqVsRyLGMVmOYBN6MSzbVAFNiPujgJyrveAHZWncPaM9fO4+d3Qt3KB/u+B7vhXMM
1RynaGrQjS6C1sKOEEm3SurE+W5NOv2Sq+qLM3IQvQktHw3qOXOEmnkbMd8z7dhPuP0W82uGPARL
fMYtkVGFtXuGL8IqSHSHf91DyWGybVmTXYpGyn9bRM0iw4TENcxRfRv3cah9DKzYtVwqd4haLqLW
+7WglShhARq5efmmAk7rgxFtYgTzjORXO5SWnfLhzcVO8iS+5EhmuWLtbc0w1ZIHffR++tSN+L8G
Mk2tGvuH7QXKCsMW/vJECC83krO9gS3Drp1xhd4lpstXDJjrL/Sa49Cl/m+EwslLIzQmSi40LCPd
tBjRtEtr6ykFUB0apbWg735MiTGt3s2O/lojGRvtb/nhoG3XJJmtxHP8S7t3Dcx3774+nGXvUYJW
Kzhwe9T9CI+ot+Ei3uqFaFMgODLpGm7ppMGkntCGlOSw2T/0xkB5TgsjVKq6gTSUTKS64+EiR+jO
SVkrxXvy+Yy3p1RbT2b63R8LZIBmgxewDSVBdZ9Zb/QJrbFG+ketf4g7GVCUWDTLEcYy4uH9bt7T
VaECnaGBWSK+2/rTFc+tlNdMb288WLeL6Uou8QWwLw4FOwqvVDjGTlNiZxq9qREGjUQj6dp1CBz4
CpYJ1YivS7zcY/meQSNT8W4EgXInvjri2qI04l2Dqbzfed91MaCV4vJ/prZbJdKsD5/uZgluL/Ko
4YGeIbX5kcFZOhpZ2e/8qYPkOAPAUVEYwx+seA0HpeDs9+4x67iqLtqvQnp4U0n/iSUzEwRf2vS5
luvR2wptVnXnmzqsSnOYM6nC2E/S72gcXftYveeSurJg0kTez17jKqMeynSyyqO9znx+iUmhHESV
kfgTDILvui3sJkR1DCQ+5g79lWefZ5/aH/yTAIxKtih6gbPvVBoDOMZ5cryELFwsiQqYg9wxmqWf
3FI8ZI+gkVVIDjKG58eZyOtRWoiUMV5znN+FLMJfOnnY3yUNb2Q+jDkwdsnUy1wsZ28orlLwgjtO
gmK1yKq00b/s77o9vzacqidAlNU40CQ0abD3ZZt0qVD68pWhX8/0kS9RFfzacATpuhdOgMTgG452
FhSyG1z3NdJzZE9lZjkMJH/5ih6iJhKXZu/TYCnMEkcfj+89TAFU9cpnTYZJIXUyYXvC8/Luip7z
m/4iK2/cC6+icTQArvFcRj41H13VDobbbi9UnG4zoCkDm+TNgIih3xR5fQtrNtlkBx7Q+pRXjo1Z
FnyYnbGLziB/UyUwlZ9XvTjhTuaorVPfGx0o732MdF7Um7fi/M4wiIXc8OrnRTL/OLy95cf3EIRR
VwpO8Jgcwca2k6zRcnyS3oPDR2bPcJoZ1yKx8obohn/NUc5hqMiHEuKPBMPMCxHxZytq3Ne0haTb
D3Wg7fKAhPcoHedZOBt1TkMnJp0woX0yeovRjZHf+ZuEC3gfjQ3xgxRLhws2IJrdyOOZhbalhHpz
qWHPnmLYA0yW0nXzbXnXWyZVQmkbv1AFKilCe6ozHc0yAGIcGKGCJMzOCS5qv7xU4MAExj7EZQIy
jWJz8KAwQVZ2KTrmFEOFQ5LUAQv2E9Xa7t6Io2FTZ2Mcm7LF12QIwh6CNSd2k3w1rt8s9W/S/bSd
AYTksNp3GptCLTxRFfApCN9EtaWAdX1r3i95yChXweiZFJl9hI+oM6dMQNE9CJMZHKe8PJ6qzk1Q
HQZt0iTIHYeRFVUpE/o3fy5wEEow8NKkvs80OV4H80H6JuExKwhBO1KKCyKko0o3MOxcH638UWh0
I+nKfPromjY6A188beXcDodXq+ZYS1KQnH7leqlLrTaUmY8C9jr2V4N7sJ05ihId0oZVI9peUEEK
HtlneYYUM+C+fkIDQgwn4roEWaatYeSp6vCGewtJZ7QcLWaZ3M7vJXmcdOaXBg41AlX7WCFD5eCi
qIbupssORw7oPONBBxBuDIcApAUdTxR6QUyFgwkXK6xCLL2lcbVDdS5+zJTlV22giKXLunSbXzfw
ycLt2b4vdS1nxK4/w2PnfMybPSW6FEsZqPO8zKKVKX8I9fH5LYVnBFO/fDIA3o9t9FyBlC+BoCXn
xBPKBTbwv3tZ/JecXcw2BLrcWxaeczrKo4EXO9hiJ4tW8POvj5Pl6tUfuwf4TGNx7djJ5uxNNT+T
QQLCbugalSOtzZwlaixykCU9eOJ2zK+KpyqGJLHtUvKwdTL8AfnIFha/kyOB8X3td9PsE9kmT10v
syDc8Us/qV/ReXq42y47fuc43r6Sx78VMlPXPLrW/9J2qA7GS290tbLfC8uDRxzsM1VAoif6m6M3
j1ImbFhwLuZMgWSkptRpF7Jz6XJS35BoMxCwc3oteWCXSk8IP8ZxvC6IswG0gXZSV5I0W5x1nvQq
MEE6hV9EK22GaimU7QAp+3Np6tHE9EhdLf2KEKd0su5MhulNiVHH/FrEWGgnCNgSHwZJ+6du4SXU
cXjyXdrCYEZn/QJJ5z1tKjQEJjjKs37wSKIA/7Z2CdwEvnW5Y2zHvG/V9Q2OSyW2uCWieN7dQj9D
SuE4zEzREUHyw6qA3lao5/HOqbiTykf0yMwpGAtgbX2OD9WoGO1/t2uKszlbuskOjj3R/4cENC7v
MzBIsDjv9SKip1wVIO3UBLOvFz4HiNoNLC1Es3H7OPbA8HyvpQdkFnfgD3TdzcwvOVevapGbYoyu
JlWHrzSif6vv5XslQkzmz1YWStJXPlRNnh9xCt8whaXGBu7duBoPs8LwsH/vWE9lG+qZKWdzeu/o
8/ZCcKP/gBcN3YwpjyTvmYMQ1a9gjdDuBin4uKOphvFLk/VDjdhKqXOjXYyvIFioqeA9XWG4XJi2
mg+QougY+z72Yim1PfCQmQ4EdQP8fPCXjB583enwhrYww0FGBrmhma3PnVL2SFzy1glaIQVMGzjh
iTZFMPZJEPP1pF4N6p65IMehl0w8Vwmix9xDul5cbNHIjPhp1HGTHn/BUZcgn7D9jsOuIEr8s3ky
hs8+tiXnkFplWEBW87gBhyf6swYIDXHMFxWMtHzGiMiyIIV9kbQD5pDWs1C6DoV09LzFA3MsqHge
PHA++ws5F8uHOFXqBsSouwJ7jNHtcrFf4OfnZgunEgGE9yn+HyHHeSOQlyc8jgyJKoDAiwq99Qxj
Al2HHmispO1chEaON9apBM6y3iEEs+A2cnKC1UfPptb0BG13uSNgq2mm6eheKCH+TKDmKhIPgglR
YRymNu6n6dV3gOeuSeGrZNycbKWMTJbo/vRCBEIru7C7Fq+Gzav5eeqUn/B5m5SWq57RCgmAnFXO
lg2JccpAt0HnPrjFmygVeFI/w/Jm7adrWJx/mKW9SvyFnSkVWAgcuOETqfNwyDcV572ksZeuP/Fb
uSSNFdAH8Rvt5nZtpGmgM7hJD6k2tefrs1SFCXDFJZKs96/U4ObL2EkIt/Ysv+XuYbN2Wfg8sk3R
+cOZcfXHIy4LV+/OO/Za8q39/lFGZcM+ybIJjiMXXvtQQWcWtsEewox71+oK311kAnT8tMFUU9/m
yNsNsvKyYiYSF3cN5CrYE5ayziq6i+MroXPc58SarHSoq3Yr3cTlRCFyJRCStqg8opEqbKEi1Op8
xCEmzWgSWrFZHZq/qaOae+0iLH6NTly2Z13MStdPNfvpydA0Pv8BRTxC6W2LXuf+in7+Koes23A/
Dg9P2NSZ/nz7odywXQmRB5SYkRgh7JWxYXgl+EopTqKnRqkxv/06vk1Rfra0mUDA1r/7jB0KnW4U
J77zDiXYSxR52MwNZxXbMy+NCg8+j5wKFOqbouKWqjPr/pJ1zM26eaVwUc20xPEjXrMvl9h+2tFz
/apL5g4ERwpQO0RQMLMu8/IlEsItVunSLdeuF9D5APxQ4WUfzAcreYUYMKtDfKWcjQa7PPHqNQDH
l1rJBt8DYAo7n6VGOyJSGMNAl2tzsKZtGrKIx5EuHbRlq/JJH8MvuLb1eWFkQBBWJYS4pmXSOvVh
CLc7C8htKuXgSbkirugNNKNSsNdaHQVfqPNgwlCekj0sv5y2ieHE/ms4RMCT2Nr8bcAz1vDVtyhl
sWUNOWWxamUhqXBQtEJFVbVUXA318v92ghBwNPOaPrpWJAwJP8DFV+McFTEtSUNAW9pmDk76Xa1n
FNxyt+KADpxW5v6XjwUAovhEn6NM8PDGeBbWyAChLESpUfMmrDsCtV1xYk7JECGcL2npbN2NyElI
EjqTAV/est9rgI43AiOfyPl9iBXMxYQ7bslRtjQLzhe7UGF1Mg0PEV5XvDNxkIlNjtR5fXy4qI91
1V5P8XXJExCRz7qETIP+SU80euP9LZcJU9flM3Psd/3AF8w6Bg5+FfGey0DAO5is4D4IQ2Xly7Ky
qDHFMg5eXQg21o3A11eUXJNBmI4sCA0yQN9kL0ynBLfQFOUSeHU8Gm4H6hy0Q6guy54+zdH5U379
SC6/CBrMa/5FCEmchzW84yHf+7UIAcAWNeFDOl5gRdt6tpDzW8PfLsyG4UIzKtVY2DNpFlNz4wc8
w3cgRHHR8Zh0ijmzoIGfvQQ0vJ8WDqmMitsvGHZIk6UeR/mU80YglerMQ6ltTwNkzwSkyA00E++P
hkRTU/vGInD2al9wNvbVhG3lr8Qi0Y8Dn+nWwLnQX3SfFce5rIopjYNloQDU20RNnFBDzjQUcBQ3
0O3A/CNtF71juX487FR9B5IMel05h3x9TfDhhWym0CmyYND6IZUbMAJyISoigr57YWorazoJPI/a
Nm3OKr+SRFUNfJ1mUIJevK157eIlt4nA+akB+ud0Uoymm24Aer/nA6EsvprQvqKrM7aWDQ/+MzzO
6YFIxAc9WFivSOLFZkZBoYlrv70KZxNaXCakAiFub1mJRlz2bvGdfyZuUU/ptiQ5MuuAVEbU5+tw
X5h+R8gxWrYY2HBiJg7jlBNLe5+t2i7ZY2fh2l4mtv5xswWNFbkRTfgoNg0KdeAgaO7GbwwCVCEp
Rcxsw9RqiijvI1jDGinWJQMLJMwlQg8uZM7SQys106ubmhnUxv0sl0l/aHld0grNx1lJPn8KGuld
pgjmFeVMuuXm+a1BYx5PdjmJOFb6SrUOvjl/GYwY9Fm7NrlU4pWz4qQbiSb6Rh1OEGfYwB8vIBxm
rLzWqI2YVhRhg+zoHmlhoSRsuWfUFy0ifAYHcUXLUL13yyhuZfmqWqgTGuXJ2+RmYm5Uq6toFbQ9
kWIIquv5K/DwKp7nwJMzDu7GgA7NrOXMN1tfRYK4IADLyDRakr+3hh8WI4owhhLToiveUSNbCCJm
Tf6Tx/aGhiHwNREbrNtrhNF6hmUKPGGKcq8iCFp0lXaaalG0iuyqT+KIXYlT3kV23ZYnc+Y3okEQ
9D48+Yk7Ze63B4CxZ+vt8+tnqCzPeMzQlbxhzTMHsZldDPpshFL2TIYFMGhsRldE+6qV0CgPWjSt
RZ2Urdnqa/DR8RyYQiDm7/Clg1Ym7rNOB8JbzWpEG4AM1vTTySehAmlWO+YMpck03GZvt/BaLAun
aJF8JeerIWZ7Tf+cAKrnfBag3QUNVsQQJD8rWJxUWlU47ytwm84bmwsa5mPgCLqYWC+f1JPNanKA
AVgkViLARwxqSIbi+9klHUM9KlYypp01mUf6Y1ZtLeVpac8JDhzq2mokZft3bjn2Cq1SHaafymG5
C0A7j/RRpWESirCd61xl561MT6IRyeBZ0rkQQcKCJS2upUmzhhr2fD+sNLDP1RMcr5aXGVygs2zW
ZpGbsSkyMIcB9Iknzczejw8YZIhudrYAQZaWqxe4rfyZ7M5WZj7VOqhjqpoXO4hN6yC3u5rowC4t
ya9FfS/5xvjVvKepg0rNAV+mB/ryCrwWG3YilhIgQSl/nAbl82BcVekt25lkDZxylBQBM0MMYxn5
1sJyXXsusmFBDxixtxR8SDi1JHybjeQcUi6sL5CW5z491z8SQRjGuz1JxsNfU5SqrKfvkxYKkI0e
PdriQL9AwhSWkw/PO3b3Pm8pfZe4jnNcyT3kuD8k7Tt30yIaSBacYdLIO33WeVum0i06mgKC8vzP
GHv9cI0eQoftQHfFU9uU2KowhVizYp0Ym5NXFPY1LcT8R6XKMTc8RsLZfL9/LEwtsdKLJd5fi9Hm
qIsmsjEwJDCpGH+MGpfkptYZ+ZP7G0e8C1a7JipyBS9FPIUi2bDZR4oSJxaSeccKUIzc3nAxUmyw
TgQ7/KpqqTzEZ0bcdXcDJ6hMmrGbG7Rl7Ent/oN4c4Rt4+ImOjCDzFGYYuAziAfJoV2fS1OZICBo
DOUp+zTI3UiJQLWuCmiP2dndGC6JYhK66qVBD+ef1/CwvHzdxJbJMHyNUzYiaD7kr3Od8zmlQW+R
FV/kYVRp7u2DOZ68HytoE4uRZHcNIsZ7mPUJtTe/KoOOSPTuKjL2hXd0dqGPy6qsD/DPzJOEt8lE
fv4tLOjcDhk9FdsTW2vlVBp9Uv0a65ETuXIbyNgkdTVAxvRDMH3Kahd05D0f3gAL9aUbsTE8TwdA
/l+lt6oJp9LLbCUxXg27jbBvXclonwdzzF4DrRCvmOr0OWwZTWFkpZot+xVziMIfg5EKc/qa43KC
nF53Alv+YMont3r7lFOwaxhumksHGKq35xXsJ7eiae8ghVxNVBs7pHlIcjwZ9LjTkzTUhwl9iI02
dIncqf3R6+HVZWjfs9aaqFuimwRddh0YKZ+XFWXMrfEYexcAySwTTQlPAs7eQc3hZV/elC3S7DIt
sbJLFn+UWm1dV7t+jItb0igHJWl3+tmkQs1K/usbYdwhSnBPRBQvAV0Bcg5UvpYR5nBkqE+Xs/UW
T2n9vR/b50JG2D9Ql3SQ+F41s4ZTvKA+dlhxaa4Ni/ufU/v7yhCLk7gCbDtxiExqns0pPeHQJ2yy
88mRxo68y7Rr2arbBvT1G46tLRv2VIcMXbC/8Jge446h4RM2KvBoaRJBFajvVfC+Rrgo9Nw3SIzd
hS7bc29pchU1RVY/ae1Ozpoqii4ZP+dDw2DkiqbRx1/6Qz8YBzB5cHvN84PPfGjdT/2qiY0/PjpC
XH+S2dmXh7v+0Q7ka5sQzhPkk/MzlHt+O6o6C799duEKqvMkU7kba5PAy+Ykhs+/3LZ4ufDUslfw
kF91SnOcqHWtj4UPkGTkTd0QIZM3zalJgw151kCJwcTvGMSnTxpkUPqhqPsiB8nNSQKw8pqo7sUA
REXLvxZDNxGOodRwYU00JuwHeMeoZgvHwXTiiqY83h6uBLQBRqcidMsggOjr4KeOkqXYhELpvXt3
wnTR/aCgDkQ0Kqfv2Ah1G9jvGP9TVWUO1bJ4+a7txT7w4I9cDZSu2faa1ioNtLwPR/3Q8wL6hkZp
Y1uHC+k+l8lVLH3XuVCd5B1b47dCNq/TFmhZmoVZp8+SP1dFKPkAKqyaRN0k7h4ZgvFm+P917/iQ
Jz1Efqp4c0DTsoJvN6igovalyOcCleGHdNKCdOGcjqgToMN+7Qn1pNXWMfJPXuk7zRRBJWRv53bU
yVSmRo3WNkQsCMUNFnbI8599tqGFWdzwHP2dr9HWXZnL/UR9ZdjuwnjEdOxUl5oXhym8s3EICsR+
PaYvekQPFKb6fSMz3bQQEB3wkiFyDaeWbHbc5KC0mh5Df2OX+OFxjOSsfJrNGM44YLFLrsLp/Ohz
rule1KnOaHvbBVxqN14kYojJ0+/id89M0ReofEEuEs2VUikKShzUQIJZfLrXdBj6t6hSvJ44B8Zn
PkyVdc5ce4/H1+pBrfUX0RXdrh9HdNYUkVXghY7qORmM1MpWog6zxkU86NIxjtMJB5pw/nnFGM9E
oJ94aree3+PDeXck1WSR6pMH49nwegCAhm+1ZkU3E61M7ENYYBECNxkpa6DWJzqlUpYpibDLGs32
Aguua4whhTtBcHPRUGbzY7x03Q0vLbEAxW3gRWqAPqrAlH8mHTScX0dd3YenjG2nVUMVY7bFQLPR
5qSmpTU2wtdPOkw4MLPY35pcYG0Fg8h2w9wJv6vcRmg515J/f5ilf3kzUr23f87zpQUv49FvKCS4
8VZxwYuK1hlwStT0aISYM9xi/frvKW6Ai4HTG+uFgiROIeOQ5viRVGp21L//wk2u5y5eBXPG47EX
NPG1WJYmaQNpcOdSnxgy3qCiqq67STFnj850DtwL0JPHsSaHlc9CbngZ+ZX7X8nD0jZs9zYfjqe4
lG8gtuYyZeXoK67sznc9qyPWNu7jDggVJc9WeRvoyz8AnRTS4aXYc8Vzs+SgKjs/gOHp40PouNc/
fpX1tO1rt/6U3X+LGXzpUWf6H5tQcywAcZEDvv9kpGyNIiDSi2Ql0tt7aFWzTbA8PRz2VP6JfNnS
6H2MfmCq0Wv5OXYHD2J9Y1hiksxlvbMvAlJKuQ0blWYvoHbfZBGXo5fxlZKw5l/wplnXXaRa9hF0
H0IzEpk7UKXg9HQbsjpXPF1w3nBN9hePAUavWQ5qOyIAVM42HC5n9Tx9wo4MbdhnCbfokFm1yZyt
AtfbFc1Lef2Cr14pXafVTBk8nRXaHtBUhizmjSdRIMymlaqXsSQbL8MgdUFEX/NwXCT1gWQZ8xh7
fC8W+qcheTxjJvCbwK2sDMrwthDcws88TdnWWvns3DxSr4MonPbB4CyMrqBQL384vYhSkvrUTIfj
s4aB49tSjUKQyiYfeawq5SvuR8GKg1ekY8Nt/X8qAi1x7f2KpCcp52r+SzaJDsR2LFf4xqDIhtUG
XwQhoMuBPF6AE2cnKvzuPl6mOlC/COQOggx2SQ/mGwgk+OwjnEh/0at7ij+hZ0HJ6gRdnLn8BLtb
IHcFhZilT+5LNwhdZgaIQKgIPMbUNXlnsEwP/BuOtLLcHmxRzsLHpVx8moPJ+MVHjBtiTGL4lRUY
6O1XAvRSjMcY0FvQ/9fupM5waLblQ4LlmbfOK0QcyxVh/04LHM/ClF9jR0lMPMaZNf1bYjGb8Q6C
Al0j2v+/rJzinFlS2wUSGXCoIIDlX0HJ6T39xhhzN3dxiJG1qDEo9z9cqGoaeh8QAUKKoBNwhxqI
yQPeNbT6ViTUseAUPBj8CATFmwG2jY0KG1AmhgPTSnFBUHxrFUZm5HRozzESZ50OQRfsQSlJv1z0
VJYpxfaI24Et6r0VO0y5p+D+nBhBupEl2znfXH1TytHbWOrdayQtfyHVwwPCXXX5sFQ5HuDhLS1c
UCI1hKVNEwxdHqmacgA/GCQBHXH8/BRJD5xVh/7ClarQmArDiPt+RqMD/54xAn46q/H2xOvQ2qGy
nAn1C25CEtp4kWMw10EKEV7hUoGE3N68mImTyhwnlTiYCa3ETlIEOGsXVVDKN2jHSemlFA/1zPA+
ef7v/u4KRtttoumZB3e2CdtwBApvaasGl4Ir78IbrvM4nqB3vRSAQlDx0kUxMwfuiOj+91Ff9gTU
wSxaym7+aoX2/L1uFnLq9ppAM4wubMTgbzZwmQhk2hkHosLC/lA0FW2VJ9tTyWRXyDvwcCWKn7Uo
hUl3SIMsvNDgHTDl6kZqZQBm7b0Yl/IXowdudpa5dlgt0fSgRqwHSJZRZWXdQQyxvzMMy8x9zE3B
Dn0DNA6Xek9HVXRhOVWXstmkBrDvCZY+tEfJhB6wagM+9JS9wItwI4Au4GMuxu+cTvnyicLwFqqg
OXGeTQKLenDPrvhrzkJa8oxwUQ+LIagvI1RaWxsCvP2Fz2jpAs2hdEgDxLxohdbK/HHAMF4p+FAP
IPEDTDqeoMSDl/E8q5PY1FmKdMKJIKUcaEClIfZfPq1DlMwexkK2pX9JTLEbfih3lxxpxhzzUTd/
rAsFhfpHjX+NyZkfNptG9yrBZfPJIKSUtiggQ1RexqvnywT+hqKgz75Ed1s6VzreGzw+urqdVB5D
blRhl3LrPn7SkkoxaQ1hL0HdrRgIetOG6UAEQTQ8UJE2AEBDZSLYQbWpMoby3AJXMr07o8f/fhom
FnOyoTn0WBsXRK7EHGyCapzLJGiA1NqXwxvDurVvjd1AsYa0doXz5q2GTIc+NJ7r+t7J7SGw0Hms
JbZ6aOi8X3cTWZzJMrc6dSwupJZWvHtMrBPKuuUImbAwguibWs52RKoOxKbA3vEjreakD4cFTURC
+HtefYWT6VFl0alxyx63/yoJswPvFY22sXf/0GW+3djfYjveh19h2uQ5LvyMgC6KmEs+8PsDMKYz
sc66lZ1z/DNWSFrWODmhG3iyZgOhdJ073vidRB2BPGYKtjUWqafb0VmmK5xBQv9+AtXY+1m3WSFS
saLu7uhqDV/d2IUjMvrXOf7KqQ3saacFYB+Q26n4aMIPhueNmMwv+D5OP9UYygUaUuLXnft/TyE/
hWDogkVhEZLxOhSyqkhFUgn+weTdZOkxwdskH1ezHnOCPMMv41y1jfCGtfxUn4IhMuqzna5EwmWb
PcwiiT0mUYaVbgkdiLQCNOQE4lAM4m2TQTtJBoeVy75Jew0ax8h9adt2WVKSlK+KFYadaqFPGISt
1xB0NZK3fTyKl1VdnOLS46r95OPpGeA/hjN/0nGdKObMwys5acEmiUPDO58H6a56eu7QLNslLL68
Vy+OIedF9LzlXbu71Ak5C/KmozzFzb42dULzErrtNvGEpZJHWW4Rw8MHUprGpvA+wG9sPJdhO3U5
pbX47H24ewSxF2JAABKsXZcjhD4363xvdncFykSISFICD30/JuI16Xft0bbRNX73LLlvTH+9LMlb
XMW5DXT7T/aVP37pyx+jti+4HnZIEx1C687/lGtefzDATAi1q3y6fiQ4lAGncQyJm3fB+/CaEjKE
4Ys0K6IMuY3HA8e6OCis8Ebxq/wOZnK6Xuvu5iSFuTFYc9aGEyYehwn6GNlSio2AQoR+smxFry6v
+Wjq6gvdC7YCpMS7MwdxoEtDT4ycV9kdXG5jRWVoKaJPRgUBQc7MespmX8hKzDRO1uyqVy433omL
V12SDhIU/3BN7a8xdp6O05JZvmNDGl5vtNvlEx+RPxWSbEZ1WKx8flKhK3dSTAFRKsaAWhNNbcjd
nQyKzJ4HIHiQKYAh5PUx+lRu9eEyohz63fnlFzI4DkciYqRCuKJKEYZf9z71XYRPtzE+dtQF+oKV
zOH1lHfgmS+4e2bc1HkBkqzzwYy5Fjgv24C0dA+CrrYjCKjt1fHACGqltaHoXpYbpHb2S6e3dIB8
GEWC6w7YKuEA30rZxtWzU8jqKEyVbGMirZyrW12QYjfrBC421clwAmEZRodsQ/xsRb4kunECVpSw
kkzsWk40azM9d2Kjd0M+p5BjYEy0suRq/Sc5HTO57cCoFKAgoI7CX53EktzUJ4Z6vz09DOCAWrPh
3RtEiB9qlm7uDreVCozSWCHs3DdYt18aKzdwF6pitCfOwpmxrPGdXjhdc/u8lrFn3Y/jydS/TWMh
/Q4HB0rSaarEdzvgz7h2kT/Fg2uv7/8g/hBe952APAAPsTIrU4ZyJWzkwB52SpR88wQ9BkycQ+Ti
3EzJP8tFnouBLvkkNKr3YGLmUyPfQB1C/YZCTV9xgfyRZsx31Jr0EHySCsJVGMeHMqDeAoCv7Ihx
ZF8Z3mXtAjbqSc0ZXC5Xd8UQa+pF2YoYLDRgIJnySUb0NaNDPkblZsCu5ExBuYdoKqfX06YOA4hG
AKQ6yuNObsIrXzoaOSuiSu3HCzykMIG3objoNLE1d9GNvoxJGAcWeFudi5vB8sc155wybo5XMLY7
GvfbuHyYhiV7ykrDA0biiziq4kCc0l9Y08XTVtbar2BfArNkLt8MYo+MY7XF259pCTaPOrGDAaWr
WfGCaGreSQKKLvBTHxaBk61+uZjcIZuRfTbDzhaDXznVkqbRPL7uvofL13uhOQ9UzMxU1TmlzM9F
bEliq3oxwaoF0zlDcl0uj6CMjB7nTy/FUi9khP9cQJp3vWRb1D2MR44VCvQ16aWOEK2L3URQxb/b
BsrS45j6P9i+jG5vOmrD9r0XHXMo9fmYbeGMxbgT8mS0hl2A4jdAme9g/3l9rMNu6u5dOEIP8Q+K
6D74tJxQwaYZccQ/9WEYqrhJFu849P/fAYU08ygaN70pyE52tp74GwxaXXvO7R4hOqXHTTN+LI9i
4X8RfnZIyTM1ZpkbxVQXxJwec+1n4pRyfhNnczqNZ6O3Or+FxO2iHk2JZnhwfSzLDuGgxcRvgDIm
UHQ3Oe6KxUqrClDjVZLSYiBpm0yOg85T/JbVpXBhEKEdHu/+eKNLE7hZN20l76QBQBebZiu6XCp2
WmxXSctJZ452oiGnxMcj35EMaYQo/4+1D47OCRpRXL1j2Lm+K8amS8hmcTpnt7sn+rdODg01+I4A
BDNzG5y4mlndtep5/E0OCpQaGV0VEVB7KhZhYrGcxdKk7L2y1pVuspWHziVB1a3AYAnDdFaOGV6H
BlvDxNN6r3JUbpXQbpq46OAQOH73sAXT9Bdq75feprgvGFtf9RWAdwmxmIMW3D9CFIgyb2RHwukb
rakAIsRkQWBPGDuj/nH6RzrSQKpeJemtv2qAR4m7nwF9/gxwAJuAWaIiqzmgUwk4pezAfihFPY27
WUbcV2TX1It/HP/rFJQIzK36pHCdGbw0pVvsjY2PKJlin59vawBbx9Ud44u3olhVdKh4x/t77Bhd
lzdp7cPqEcLfYhYZ2m67IA6cTm2im/KsVKLFek7ECwA/VzgXMdSukIS+/HOxrhhBJzPtdvk2X8ng
/H+3CVqCIdn00gzdQsATqNytuL0LZlTwJc0u8R6YwidOpASJAQsiQ6JhP5obaGmhhYowo0eTb1LB
5aXPQfgu/JtD3gA70Iy2H8b15xs2LBlaXJsmKL2o/65bpMPHCLDg2Xi201iZqJ59orTTrMKbjbNE
U3fiYcHc39NapjKysEmUsAXnu4wXsqViYrJRPw9wrTGNjrUCSMo7VuM2GV3S4STeww9RayDFcxjr
Iia0clmfp7Bf9l1Ak8NcQwmIh1QGBNkPWz76CEscZWcjuyINHZa/TkK7xlr8Bf3r98ubDARuLiwt
MHRJmWvw/OwU0V1ai4Xe9qGGX8klubYPLdFiyXgmClMqUEM0BCBt9z331gCrLSG9lxffNvT7Zvwc
63G4AbsIGiXd7ly1YyTcxCVf7heFzZWiOoR1WYfY5Xz11CZrTR6V5K14UuFmmWGUGIhWEJSxg+W8
nVop5H+g0OHUkvJA+7bSQTNVvzmcnx0uVmmCzfAMT6WDVY0FWSnoNYlkWquu+2TaRECP1NjzOyL1
N1x5g4Ar2w0CAMfZCc4ifYrClxNXzW5ZGy2DtYwDkV4jslOOrFmfi2/Upn73wUIaOGjcPhwEBmsx
MIijS20xGNZhYAYEPIKLyB/yFK04I+WdS6q2Oa6Gn5N1VI4BrEOVRB7cmIKTwh4pprrDpuxEEBVm
ClVUK3com+HjsASbEYAYkR3HEf41RaG2XocapTwn6c6ooxp6KVKwXiIpgk7ihaVi94NNNxWjhUEQ
fS3KAKBUt/Zc6mgdAXV9CHQcsaect/ldHqiWVpukwOYZFmYjOTOpyPzcpnZcjql9Z/qSU2bg9wya
vhFtSbXwBIPPDqV2x/NpMsKvXBPHZHGlLDxdDvRjRMTua0KTr6uhBAsZ7a1DNIkbqt14xOg3x6Ay
ccrS3MOSHMU1t6p3VeGgT5LHQfVtDMz0L27KxFNkIgOdY8CRgevU2+1569ncrhN2b6Nfj5u97wMK
4W5v7l5aUmrrjatujuE/KNUU0bOeWIEK7sYO9hGEcCpBsXNRNDD4iPecHKbVok/p8Xrjl3i24hsF
9/oY4GdTUvVAN0Qz+jMAZoQfhqWZzG8GP0YWz8NARH0BmTFJBzXAAFy4Z7vFrXWKCzB/hJaXQXho
icVLJSV2CFTzjk/JxjLjTcBrnKxx1mlLXANGV9+VK7ozlth6ZPhj24Lhw28XTfJu3e0hx0M+Hljq
X1gfG/aLLBQRMsIAQa9iwm9/RRNV1ksjClhRHNU5DfGZfNTJZiqqSqm17GcWglqg1Kz3fSuJ0h/P
IeyOTMsAVVrFrz0HdG0VzjjzFFRB+0RVReLpXscDiCEGfqxjOpzv4emLJLmqE/AAKJ0eCLy9E6Up
bgms2KESK/y4LAyC+KbZYfwvljvUxcTQFTBGrpf6PyiCXWZm8sJvun1sxQCCcXOFQepDxI3YuBc9
ufskaGC2UPasGcgoSIMxgCbfMhRfHelu2L4hw0pDUFDWSyieg58/eEqdgfegc19hW7koAUMoQHoa
G6INst4luPzdVO95lbkIDmwzWOm0k3z/meoggTobOuPrR5IaagQiNdkDwqS7NG7K/8UqstcQcumt
a1EoWZRLzwI5t9PY2HI9wuinpLIdrIp9QdtHREiZz7QSAb3KBd+czV+/VpDLxlVCO7ImhiaGAx1v
Sf/SjQrk2TyAxL/L0yhZdJSFvl31M5LtbBonLpMfIXOmNyLR+AQegdcFd4JkXmmwIQLaNhcLBGJg
ffiVgfj/VHWM1r3oQcQDEPnXQCoWxxBEpRmPw811KTUrNnk4vKkm9rjRp4C4o3nX+cOVfLm8W5/Q
D0q06ybCuzbVa+kcDbGyeWMDnkUkTHAj4G1BavN+1uFXBglifGW/JDiM8NQjIw35K/OU5vGcBrml
oiSa2naeSXJb2fL4KOpgj5yk1e70MD8e8UJTs4u9mi0H/IGkR1fQl6AYIJxjYW4NRD3AIYVdDLgs
44xEIU8RD2V8h5FmMy3JpAvlq4tW2m3GeISzT+ho7irOxTY4AuJfe3d+Q1zOxHgcdLJMoQ+Minkv
EQMUkwnXyYZBLWW2y17tm0x1VDbvtDkKC73n6cCpRz3lfcLtDnF48LQmSsfmqGvS9AyZs1dmMAjr
/GtQ/VeYy+EpfaCs3ppeZVCst+RM48F5ij7zuNdQiLUUCBSuIodw8dVkTUKKUyomCjUC53vveyCz
y9dgEzCiIzBefShyLNQf24VfD1timQ2Jwvy1ckWJX6zY9S+Np0pxdTF9d+wjFFEccqH8caIQdLFn
Qo2g+DLT+Fpab28zTY49n28aoobNZi7prV7RnDIcY4VMBNBC9h04USsj+M/DZtYF/670isMs3whL
0/OadPfnlf5224V/WkwAaOgdwWCADV1tVhNaCLLRd8t9KMLhOOTje9n5eCovLjAYHLPfpIpn+uI3
kBLrfihFTLIeYkEyiPQzFer611dtKeSicnSlH7Nk5+Fk7grRad5foHX9Te36HJJNsDQLv5zLnVrF
0ImWa80/cwAtkWlP3wLDkY1s+A6Lw3LPJMQNmIJMsiLPFZ7qcqq7N2TCRBOehPeOCtnK7rG4fl1G
hnm0PBHnS9838piIO+kXiyPlW8HMll7YMV+/VF+Oyu8ZjNxUPg5uv9nsv/yP9Ru/C5Gy7O7MEO7Z
VLWlXWpMuIVRzjgXbkivXz6Sut8fvzZjUpwVPdxAcZh65yfaIo0fnGYATHQK4Ktnx1SVaiSW4jUF
kIyU3ephu8qqE1VB5Sf9oB+BtE6nrYfOGOiAW66lUuCqssmaxtZHPv0WNRVzH1VWkZv7dfON9ate
tQZ+mWr8P4Q6i+NJem0jm85TUnHIXlmAkV1y8TsHraXmLZmig0fI3e6fNk+ikMHgHmxS/bbwYKeN
JKqaFQfg0xHgFNzItRFMzJByXB8rFbW3dgjGSAtHZAV0RT5UJDPNznFPJW/BxDVOK5nyIFhh4+Nl
FV7Vdi2SJUuMF1qbk0D54fAubrbtXTRQrVJw1MX1Sm+O7Rt0kk8efpRyj3YaCALzWP4N+Idxdm5v
d+mQhQPh1odMqA+ukxe00HMrtXsStkupyIQl1F9OYpPAE93iYCbz1krXO5b4swbkNT2J60ol9M6b
s+UvydKzYrOVMH1zsrj9Jl5rpEexyI8Yl9mEHQMf3Oby2saB691CLktsCa1Lh8AtSvkzSw11CTFA
XXZL+DPUOohCuhh/h7Fu9YK+bQXtDMaIceWNROIAbhxOK7B5HosT6wNFmpObhMKabjBCQNL+vw5S
3pn9DRlkQFX3fZGfS2jQiaKCl0DhWgMMFsydh6oQjLv7WEShkMoeJU2rad47/R9AOU4zrrebJr3o
Q2bmbgrMbQ4mNn1D/LuFd0SkwW4kDoGAgPloeO4NvtDafIc1+ZiKOc9J5DDmDjO8rp1fs4OHlT2h
cMOGMZEIHbWaM5x0yv1KzEmR+OYH1jsKS9Av0XxWr7TkDTii270bCpUs5NH7nr+GuEZ8ryb0iVf3
IcSHwn6wchUPSCB71J2ym2x4iXdilY4JAbiGa60OQsaLN26xJoJ8rP8VB2R/36kQjwWccII3FU9Y
oFSaWpoHVUWeBye5TMUHJIO1Kl+4zjL4VY2mhidVLERUTz2ghIJLaY5j+PwN2Vsg9TTbo9MwnL9B
ym8Az2qG8NnBW5IDHj+jsZbN3WkF45LvzcZ5Nt1lAxWn27+mQGMkkOpXz/vdcdOplYASHnW5UBLE
qiKn9y9xsMnaXmj1jrzAF9HlJwAU26L8qLltt+AYO/ojPjlOkzcNZuZ+HN5nTB90Vvdu3p+lNdOG
hDvG4r9mnIxSfnKx1eM0S3rxGCEUHI25RdZfy0m1gFujiZ+DSIgcdDo/BJ6f3g7u73DYsMWWOXY9
jMLPK2nXRh/oP+0gPsDd/gDZQdhDRxtX8BhynolxaRaVK4VibUGHOPBIIt5n7HGjKONEHk1920wd
4yhLJ6J5zzHtvj8ESPhwee6oW6QxSOTx1o+US3iAVv62mab8sDwTF5DSzCqmv+rcB0SAbcKg23Py
nKnW0XAY4z1Bn8r4PZz911Et8eRMleOfg9+fcBi+fM4lgJ3/A0BVr7R4t3p+hxCMLCNwM6hqEwOX
iJOPGX5eU2nm3BIrrueMfH9Z/kUwvPr8zB4T270J6g7Kn6eU6uWSdF05J54QhCCSeYNKONn5wn/P
9y0Jw1xYKAxaGmTNrBDp5OMEO2snl41woumiRSNEuDlSXY8Q8iMynHx1BIMxwXgFtSZnoC6dUmh7
RPGKaHQZn1EhnZ2sv+iLC6PYF0AZh9RKCwds/c2s+LgAKPPXMPemGocrVSyIyg1GKt+uv0G4cn8j
zXMZxSZ6BBXl1dbwVdR48LOs3w7tlrwzTjsmvp1QoKYsqxz8tZpA7jCwZU7Xn6VjrUFX68BUlc1z
E2rDNaV0jjz1SJIRECgD0RNhPiGV+s2e8kYSZ2Fd/wmN8FsBY27N6RmdNwTzLCkC+wiPCJ3BbRH0
xMTH3kOa/zbwnPkQUVyW8/LFu08rBqar6oIOAMwqM9WZYeK/CS/gWFcPsgkaiE+Kbm9cVrNCtlJR
CLEiM258X7ZUg1Q/xVBrMWHuMrFp5/OCdTzRg8XnPxSOZzQxUMPRX5oD00b8TLip9rM9SICVA2xi
1ObeoXfMJKOoNKJXnhstsaBNGXct3jWYmu3o0GoFKWH5+8Pggki75sc7wJdgjNq++3xJwuBDLSZa
fvOYRgGERQ+X1uhWzJqp9mhUcn8uvy+ZE0tf8TLlEU+k/65uP3gTJv039FfCZ9xkmO6JI5YRqzHE
iILTlgPtVeQ4b47otGZ3iMoOiczTkztKsrLbJmES+NfZdJRRDv6LUnRyCgXThjPA1PKWtYb2YHw+
ZP25As9uua5q7CyYl9UQIAkDBLDW/SiEowLf5IuiqPsOnlIfTvYd5FCYOUHM7Yb4GB2r2dCghaGJ
fBkBcYfU9CjFhLFf6znVfl4h3O6zXMehYIFhID5QBSjcU52JlmlTKCcU3vkzcBkUIDXBj65NPfHM
TfLPmODw5/KX9Up4T4XegI2GbMdEiVSNjHrmZx7ZjSMvJwmbhbrRSBUnG3/p5f1dwUXeGlfIFzUc
s5YV3ws1qnx8Pm3wB4pc9stdxhm9d3hXSTeg5eZeSKjLnT0kAQurMze/WcsaRwejAh7H3elvqyiB
R5JoLeDfFfaIdl13nLDhvtAzneor81g20WgDRKJDdfkL7idgf9Uf/Jb5TraLOLHeVEgYw6zCv8FQ
OvGTJo852/DomW0rPVzAf5tkBTJX5p2i4UUvfKnjYnAqsQaVDKtia841PWEn1D46Omb+aNN8SXIA
PrXOZFxwayvse4DqFP61kyP/Ot+V18+aS4RRl2dz5q/N/DYkfaNhk2k0wzxSAKUiktB8PF+4sHKu
++pJDPk/qEzg/yg1kQ+Hqa4EyDQdpL3sDu+Ztg+iDQi5hO/BquZ9n/m+uGUYI1RwV4CbSZlwvxKP
Qw6LYSEAIU3cr0AN9raUzHoKRnpVHWXJ18JwDbrodlR3mCGYc5GNC9LIkxLdsVMPkrHgm1X4TN8d
QFLlt/CJq5NDa4kETLii7SM6NRCM5ItBvHxBP27ZWwcZEv0GgQbLttFRvuVKDfx6lZk34BwWqyrj
vPPukTki/dw7LwyWpW93bppczGa3fLUAXjKBjoX8S7nLc2NHVpmJNdxmm4G8DhYCSyx1V2P/OOgs
TKGsjAOyCz9Q7Wnu/p+N7FKUrHm1SHp+BNMUsN6n5rrUEm2D60eGeFHXfupzItQgdjFSpTbi3P3P
/jhZodODRXmH8Xja27RkrGfnckGCzvkFuDdUk+OG2IISRnNMGG3EfNBOob+68SaR4Fhi2NR/jOXr
79HJgN8NyVEPh6IRBwlK7f4NOmcTe9KAa6K5hH9BRgJzCiuw2bvKrxEvpLINklgaW5R9h7xZG22F
GpXG25CzKiqA0WCERR0OVH8XOLiZ2a9/oog0jDMc6c9YczBWujsczuWe3WnYJCHW26GmMUzwLMts
HhZgumcHs9TzvlSbNM0dO7bHcZBCET7ZcyBOXIx/Q3grIy5esLmGdDTasFxRYpvZh6TlH2W8rQbl
XaocMdnFen/iOEn6Ef31/f3OKWGDnd4pWes3RVn+xYUGEOeaUt1joOfkn7BFd5i5IgTkyEtDIdUV
sJBWiznBd47TCiRoTHi3pVUUA3O0n4YpxKESlotTXt6+jyQyBUnAO+Sqy+Xlz0ChMVdaMKweCSgC
4SG1VhiQxds6bBR7QT/AMaaHoLoOFhldxvCUQc8GWEmg+9bpbpLNDfL6JD3OAVtwBMM3K80Av5ff
QpR3IbdqgEhOW57gIFS2waRCxDaNq+8Q7qtItoEeZQxh3cWoJob98duU0dU5nFVLIUcu9d5C9LoW
D0LBgvjJxKgkmmpM57kZGrLdK17zgZhBGWzNvOJpc33Ozl8dAQFhlgueRXu2WJLpZEBB/r3C4xOd
yr9fA0wRxpoMriGHLdZLzR1zBdNNj1J0qyalfm6m1G3uDwFLme9kLRW3mYQM4/oNHSdjyGd2VlsI
Hw9EqTcxSyYI7WjLAAykBbVLGJ7k+4Kz2sUXlwFAaumJUZxAR4/lebhNRyHVbGw0QnUjOZ/K7AL2
G5K657RsPaf5uYKuY1A0WAhyICCGMpKkNV1baOPbu7Yj3JKoTr9OHQjXoEGqEskI9Vmw3vNz0lee
edjr08FiiHjXNcyuJ6veuCDjS8UMunP+T6uhLb6YKErrDZx94sDfkOZzgYDmS3ophkke4Ms9BXl2
6LkeSiVT3C292uBuAUlLKxTc/BH67SpEiBgffk3ax3ikee0PXyJ6BppFieX9K5py/3ZXB6G9LJ0e
p8jygOYQzt+ZkYKRUspNVejnxw7M3SeSaMi5zTFjB2gjXZ9rw7fUt2JW4eEB9UJG/NvraZZ1Xpm9
GBWpm9B+LKQogNMHf3rmziE2oIaIeQUYQq+NJrr4gIBsAgjSRTt1xKaDbyVe7+GZKeYSUrqt6NcG
GQj6M75f0tNLQTl2zRbpyJMgoDaNOWHdG2gzjc0LKRavxQ25S/CnBMW4rBsASMrmttBnx9xyGsF4
CDaxM0NAJsnjL2TNIfvXHeAfMI8LK7zv6d/eh6y+FG0LwHnczslS+Y3Kxkuu0hH5fQXGhcCeMKbb
CogUvfqCpQudQ6jEut2mugw9xqbz2HwC2J9aUPRd6miuLjYrLD/A1gbG65P3XoEwVtPqtZJi/Q4i
Z23QWiiVhSZ5xfu31oqcfd3mTJWa3rT5eKUPyydmxrmGvQi740ZE7Gsc7om9NXiR8XO4AO9kr8K8
1W3vB6pAdocoEZF59UJiF+M8NZhDhvNIRBRxP9mJhQVmxrJaymgSnL4V+OFENCWegLxXP/31LyB3
sC70HY3kdYoZkcr+AjBEjtI85FdE32e9aH6+5sAlKavndALZNdSpGZVczpGzxxo75/PMLJEV7i0Q
NVGyukY6XFRdQML6yHtXOXfc3pqop1cQ7HJuVIxAO9U3gzt2oa+TH7cDE26TpzXSHV8W4TQ1elFa
j2xTIKqZ7sJ1v6bwY5WNCvoKn9TSpq1LPuAuP+4nK8eG3+aVeCLqv/cb78hmTT3VegOpg/bxFwIv
PjufBsNok9ZSapR8x4YRb82AlJlMrKq5DYAf9Uy7Hz3QCOevgtB182rr1Sa1OSvaIB7dv602Fp7O
BCuvOJ1soP7vnH1VWKnuMFBvoEDA7ZRSthwHsFMic2gFvCgVMRu9azNG4D6wsYTdjibqJCl3kncV
oUvmvGcnC+B6vieQpKft3RmwOT4uyKcxdHhttiyUF1xW6mEsthdBD1Q608GpiBlxCXmbZ/wW76xF
F3vLBJW90rIPq56r+fbNTWiVkxEMYuyNlyypx/n5MVsMnBjWWmScZb51Vc5KksNSlEAaekdz/YLJ
ey0iDra60HUMdBLTipsmbJ3xix96FMZdJqO7X7T5TFuNwAhkVwNBqmspJxgNp4+KoVSO7vP4sstl
BRA65z0yb3ll4o2FE484Z6m6va3QWhVI0ULjdXeKgtKOx7JQR2PEHBAgbXzGi8kgxXRkPSlqggEJ
m/diU6B7X5JbDLB48ku/nTN0SRtUQzol4Et+qdbJUL+gUh2tMvNbPYZWiQlp5S1SS5AV9ReRjbnk
WUbyfDXNUjMlR0qo7ah333SryAKV2qUn4XPgBgDYfjFObGdkVDTgWtbxO5b3RRHs02zqoi7t9T1d
XJmNUXCsN+QIuK1kyKJWcXNJWFPS9g5y/sywdsbtQDEGBhtpoB8Be5emJA9ikiKE1qxgnkDXfx7c
nPOro+fLAPZXpfPgvo8/PTCPTl8QjUTQPWjqH29/p1/PooTrB+zdwd77CR3L8vt75ndSoYmDTZN2
h0XUn3HfMpKIkf0K3QKK78MLg7Rs8u5nOFLabp2GvaQVTIcnN/f3rLdxD/8g8u883qfnj8SFZycO
7nEpMW//cY/Ru9feWV68pjj6oaoIyRqqsBCLYB7BbqjAPtrftV6ZfMbybP1d8kvIKEC8kd5c/LFP
UXkB8E1Lq2r1+eCulsSfv02f8ZBwu6EeTM2Vn8nE5Nq8tcaWQRSA8o3B7dcfTeI/xAG5bF8VW31H
aG8rIHRcKPpM5Sow9zt6Z8TEsnUhF6YTZKhBMTKQIqAZm0F6YxzJJaG6BI2XnWRv113NJEXMWNDN
rKp12/88/w+Xcbi8sZygXwst1mPYGz5LF6RCtYkBHoW2SZgOyoTwoW0U5khEmZvRBtEvMUPtlzDZ
1BXVuWiYxV68M7B0p8hwz0x15Y+YVSYTpCJLtAADChcDDpqRUIiNz4Sb3qxTvRUHXiMr7WY9jaQm
7Nz2VfHD5YsQX0cXyzlxmyocvmUqy8So9psTj/QtHSYm1U8hQhsLyByO95klSchOXLoj+sOd7awC
bZGEY1sEXh1RmEiWI67+0g9wtmeS9qGC7F7tDpJ30uO6iws8mdXSzQ4sarR1YuLIgiKUhmgm6rhs
ALzOsNoNWqduZWEg7x/UU7gYFnNTebv6VLfqUYysmKDchi6Dqa6miggt4WXeEh+7GbZx5M7V2lLB
SI6poQmbNOfgGf/jH89VmJEXta1sKynoQvVARcgVq9eOi4SOYhp5IPO44lOBlsWc3gyrgload7tw
KOzzSfdWxHNGa/UzSQTgrJ1jLQFUowFriG3t2zsPa2uSLHVhbvYonzXcDDYfS2r+3m+BAalTCgYp
xoUpJYbPL7WX6VL4dED2In4QLGtMS/iKM2C1jZZvTn53Ck63wnUYlqlHFfPTvRavdzZtBDMqz6Bi
cGokH5V+ThQPVcnoG+xcnlYMWZ9GbZU5kWFhO40w3TqXhuqHUvryngxwN4p0KNnDsxvTsr8Al9KS
91yJvQYp06J4aAng/Eokjs5W7DMRfVmVZrNCUEWV9HxEQfrAWkTcFARuCrmVxPsRUOs+kxbaNHSy
af6E4tfl0NXWNYQaeUBu5J80EddCXmdSqNJY9L5OZzkwhEs3yXdICVTPNJqK7mICm1H/QH8hltdJ
eaJVJyvLmGw2GP7ZEopT3aBUfXIM8KWex/nqPY0A761mJTCk1K35QPEnVX4BF4Vs401/gdWp3ifW
8ZkfLqi5ezHa6XKTQmBhGVmjHJPyvy7ejyamadjzSo4LOmpFVgFeDZdFIXPX+Amtiw6wEbr4yGvP
nfJL0E5Nj516vdVMSbYZ9/0bmsXvW+DCG512CW5XxZ6NwB84RHeSIgCPMAsxvMx/ryikh9y+fQcm
UouUw1E4KALmoeaTuEJqQ2iIDSSn2CHYWJO0wO4tJPyTlxgkD+7Ij86IcSiibKrHuS8NIWfCEPkz
JwAHy1QCHQm6uYTD7di3RU2UoB6VNSvbzXaWakdiZNH3ZyKYd0mcsLn1Kt19e2i337YKwNmrefoa
lAyy15l1UcSLuW0JZpDMiJJcLXo0kh7Vx5XMJGrS/1sfKT2stKWxbPl3udcTXu0veWVU95aHn2iI
X3e1HIrEt688u3ddh2SjVXR2m2FGSLsU4JIbdM5jwt0KQuXZiXCV3wbH/rp1B3HTtP+1wzYJnoqo
/SVAs5WeiUZ6yiK1JalelOBWojgKi6hIzivAPv6bHl72JiKAagONuV8DPsHipwubZf4nn+eW6ORZ
vSz00odRfe0tf7BHI1Qe4QvYSAw/vjLKhGFInuf8LRI0zwsvAoGMLUw3kqhbCJQ2raqA3jVbypoy
S6LHuP7QeHzYGUpVdiKz/irqbZ1W8RseAhuycXqxA/1Ir6l3UqfuY0EtkguiQRDkLWudptqOGfLa
jfPJxvDYkabMqmt8pAPwM4QaX28U2LQ/ivHNeqKCxUJpzTUIGBaN8hN3eAy3r4wUXHTQgMS7ex8K
zX4EmVU79nx0lERySU0T6QuNaeC+dasLo0fCRZ9Y71ZqObCAHtpGLnV1I1c5cW+YamoN656u+qgK
9EIejQ5vAh1aj1BTHT9WYKXbAXukpuiapu3xvE6OinJ5Bm/+UfxqXEIlACja6yeVHvvA7mZW77wz
bOXpbjsyL8GfpIBmqSXWfaed/u9g3Atzz12lDG4Z75l3MBBiTpGOKYlhYud6uTUwFM5mZM0aZ71U
7vZsOPfG+J3t87rBY8QB8NFYB7XKnfur5qhnqSCS7UleBP40Pq6UC2uwyFOnTnq4y8PCQivYiI2p
PZhtYnUXzhuwa5eYFuRUZACw6LWhWEvF5MoUnWQA3EychO3WoKGUoI2mCIVFAs9LfySIP1WdnB8L
taybyvzsvap+udP0xzYr3pV108RobXzO2XVyPZefmC3dNKQsEuPbyfuE4JKo1GrDs/GBLzXb5ouA
HdZNcNaU18rZK644AkidTj2bueD85JZ9FGTtGJn7zoIH8qb+vUExQyVXxWH6c3w7Xw0zthMjBTeC
F5yJsqQ1lNZS4x0vMjhSrOqaQC/R51h9/LmIWqzAKm3cXGqRM2pj2i4Hx2Jwv5JvVpm+fG36VTTZ
engVOCHGCQtR+ZjMCj0AklUc6qz7oLOwrD0Yc8A5HYR8XYlGfI68tO+T+CX0cVeY1UElWiaQINQP
1k3vhM/J75e9nDhqlmEcmb7/kbS1V2ztIkNtWvRHUwEYwpblqg07qVg8iuzBjhOGldwkah98wq3B
Diu3SDZ4i0lMS617tdl0nFubEubOIIKUtDe7X3ta6iAnknXiHK2SnOozh79yksqbhAqARJeugPPN
iqhx5JoBqezCKtrAm5N6LY1Hz1rjLcHWFhNbFCGoOCLQMAH8Y1Jvv/OvyhhBCeeN6sE2MYGVSZct
TKq7jUE2O3Ueuy4xk8VybB08DQGA0tqsICF8ffUjcJZSAtvP4an3ctcnr5zzaW92FO9JWxgnB6OL
IYCpmgmiLtJLGSE4RINFSNQYw8OymQZ6dtQSbypSeZe8rYNkZi0IbWVi8qZSxckDYTWHr5sAEFEm
Pw8Tbd2KZZ7xAfq2N2zox8tPGTO6QWZ0iMHK6hnkeL8jyuQ2mt9EODbf6p2+qWJWQNpK3FLR9gwS
otrHkVyxPxFQ0xftaoMx3w8gcXUL+hvbAMT1zXb73EfMRmgb3jB5RzBRJ7rwwiXgYaJbGtMWOOPP
xJKbSUwsHiAz/QRmFCyWbqgrW1w5erMdYvheoXlRW8qNqfmTb/PzdHpIq+FGuC3gTpOx5B+mUlLB
z/pTF6LyBLADYrlnSSYqlIdKqlLWCnR94RK/1T9vfwBBfoWfbz92y0XaFyFwAsS78uvj83gJsAIc
RR5AEtXNc0ApmCb7p+ZxTNAQZ5euLjlL5Ya0vOdYEjXxHpTU8X8+n+fuqy5VoznLn3Q5f+Fm71IW
9U65gmydb8MRgNJyNWRf0XUOMeBY4y5d2t6RwUH76o0HjqixzqJey2cMpVWeOlu0P9m7nOsghAJ5
48QJOYH6wJcHz7SHpStVgC9+vHsu5FF8vFQzfPOqtgBzm0yx6BvhWhquk11ZBzF3ITN/9PpJOU1I
b97lQEhREK66gRNtTBRH57EPqXjHysYl1s1Qn8hZHzS0f1A5cZ+o+ZKss2vqevwIcjnkQ97AtC7L
YDcExx8ioDHGZXO8+awaknpxjTgR/BkbuJtdbJB+vAwHHTaVyin/ezEMxa03OVBiYcaYtLjMa4ln
KR8XBZl1TBD2ClQjIALBuvu5v73dtrLjXqBGsPh1rqVK2IkQB3Vh7GQTdVBqvXpy9w/RllXgjDLW
bhExxJ+vcbJ5HadWaYrpCV6Uar8LGK6083caEqMb5Srxe0GqCgXo/MGluKNNqebzWEmGONGEeSQb
dtm/Q0SKlFD/F46txCRuDnwAlGGGaV7W2Wk7+8AtmqZ8DsleuE/YoYoSih73HsIe2KgZGXyl8quH
fK7SnKghnR6YFns8OgS31dHS0DhNWJZNNGoRRcgvlPJbmUvyR8X96n2fuKPn1J8jFPdkD/GuUbgD
hw1IrNaruP1hpsDZkN8FarzPFWdDbMrBsTl5a2FjO2poiwPzL7VvXWQhqhZxNeRVsEWaN0xwKemV
DsZbW2efseqx+hDSccAN8KGQRUonvDWZmFOinzaQrHtXXGgHs6YwvLPVJoMj5cKAC2qxsz4vfkSG
DyfjORSQ6TNQr2WbxhTQ9NLlKe7IXEPrXSUZNtQACu9VlRW4x6UMtUK6y56C0CK64fnPMdWk9QdS
/6GtMwmtKuK12KZhbsucujRV0on5GObY8XjbzbTKoiDv7guRX5ZEASZk1VMJslX0iLnH1e/5z9PF
6Ge9as4zmSek1HjIjrxe/vuFjZvbX3QJsqMMwZWDEg9IZObP1O4igdS56d/bLSpIuszTIFmfxH5X
AVK38mDqXty+tRUgIvh7+qJmDZn357fDjhJqJerAGOK2lgcMAagWg8R02CGvtPOF11RB59DUt7vM
yuH8qS9+Dx2zL70CGZh6pRl20EEsaEd3DUbcx/kLBrHkXqkcDelm64xs7UUqadXGkD30gy8miId6
3s1Y0jd8BUVUCToYfVCdXkXBHkIXGXwZSYXQOPN0tF/J6mGv26zbkIK8CPPq23g+XSUu++6eWSDn
TghLXbyZ5nKpjCgX8MVtEu3AVGE1Mw+2apd/sFG5WMt5Zk8fWbERA5hqFuE7PbspNBlDOt8CZXa+
fvKmgAI392Tnvs/5voBLt9ntcm8h/HCICVpb34EyX4yRO4iMnF/skX4QhRbcGuJbVdGivT04ib5p
TqLs5UacjO9E0T6xjDoj6whNay+QZXWl6b32Rqr2FUcexDbmj9wlcu2TPoHuhBksbTadaAqjBOFk
DHBWH+I5bDkP+U58V4lD8v3yoLrFPZ3fAgxejvjUHG447GEwApA0PZ6dEQ0eWFjeKD1EoIK8WfK1
yuAhui3En5Dt19mPuQnQwPY01QHk45RroueXdWOXnbyQM6ufo/MkruL170O3MbTuASq6ZRgcDIYU
SeJcT2dzVAoKMvapewZCKxNlro8qS/k8AMbd4pFbHMWwucp8QeFn6LlWCGoaJcevWH/z7MVPg40M
EYwfUBlRGMFRbuTifz1Fgerk2Mcn+OxxPGTfiQzDQhMi/KWI6LPUGnSv4/246Nhc/AePixOU/dI8
NJLI4b5I0ofA4k2obRkMHWGPr62UPE5NKbEIMoe/tY6j97WTmxhh3GIxiQcWr0QZK6xoJnpat289
7vy+QlJQGtmkW2UWbF2uNAq9P+qpLYC3EGOzeRV9LVjAr3fJXlbxr2lPMg5bzAoD8kbIxcrM4/de
WPTTb8J9zW7/7KkaQ9Ygh0juiwe3QCigPcx1G/8dqr/JbgcbIlijPBL/i+7q7AURRkVHb5CuHlNp
Ntfr/jlo9SSmiSmxKWirR287Z4w+TvPrhK2OPoN69Ncn2sR5FanB8y1eU6AyD7fPiunZGVO1Qzrl
DVB9t80+dqSd93q5X5i1iFcfTDM0yimdHVsJpylrfKora567/A4d+EIvtf+EDYLRraNEDkiBZsGT
NFPoMy029zTi2shEyHKsIQ2CXgTvE71SV49RyUmloiq8SfaxL2Pib8vC3IM2ImYdcoPwA2JfPaPe
B7wqHggCDaWXJsPi4JYEOLpMn9MGgi/YxgeMez7wJfxVCfbhtUyNWdHZ6cn7eQj+yk2A7HJoBu8E
wSjjrKXaVDBOJ7C7dNvz5L5v34S0kTlHuQ4NLdeFXsOOGFUMML4i7v3Y+cqI4NccMkF+1oiJXQit
NEYCvhRDOQQHCZNycZ92NcnFV0Ul6hkxBKRBu1spF1242N/b3MU42/BoXJsOPLZTzq3aO3iUz6T8
XMT6CH4KAWX35fac3Y8ff819XwcJjgVdBW1bupFWgA2oDJcb+BJvyDzwux0tryoAcIzNliwNfvkG
iFhXitSAFpwrqLjDgKqSFNjmrkfwSly7UxO3no9e5esIIOqCCYpKVIPacDmlbp8bx6I2irXTDABR
5GEYkfJGzg9sHhtG98UigJEa9/4KBCe4kd2RW2A8nIP7FMtbKp865odidA1RmC7iEfzJI4L3kKHc
STIHIYA9hUL2UvaEaFy2W+pL6yKx/P6efUd/KrhLnh1I3yL1yydCfANkfmq3Hz93wUMEFi07g20D
4WKkipqj3bHpTonZRPEdAC1qnsVNOSF/EwQen3JV70WjMynoNMpkPdXteYqdhJeKoB+rBrcjHGAY
b+tXr27qNZEYVm4tqfVTYSNVzja+8kqgB0CDfcJF720k1zwngJ2xYbrsR/HmHNmchthuYgrbB8r3
fJ+w1tp99T20UKz5T4Rm44pEzx/IYpeYnyzcBySW0JT/xLtUieewc7Klz0PbNW6mzyLi6DNeL5v5
pvY8ztXBZXVCNhNnmAHvkBu2XAv5AySehzSTtiW18xBb4DuU/7+Lv3nsOfTa3gmHToTZMi+gQmeF
6jnsyUHLdwRcOd3oP3K1VHCMLPfGublA1dLZmZtrGyJeg0jZ8vq+obewdQUkyUxVailbr5LAPwUz
oUZjG7QiGcy695sLqZV8x7ed4/cGIoYXjETP9YYR82v57n/SZkXd6aTfGTXCxWf+dyHkgRV4FlrA
xBSOBP9pqbrkHl8ObmRQ9xq/hJcyz9r/5Wd0CxCjMd8RsTXuN1q5jVNiGgRZTMfcEhY3dBwdiDBY
VFHN1JzKiIhqFVOHGc+Iaf8bL4vrnc2C2v9/Ib5KhOEBDh15uvEU/DmmFMESsW9eF1nRBvH2vGag
kjWuaoTIDq0ReDAoid5vH18WVamdIPp3b+XHY9otvRUswL3hyZ5PP3ubSflF2WQTLF6qFcxhEaM8
eIVSpF2dZqe/1i5ZKLoon+SSs8GJdAKYTsrPWqej3b1mMfQxbrkPZaKXjeKhCNRqtzWwj+3IPVfO
bBdlCF60Qf0xVb2OD26Z8d3FrWQUg6vVUIMthOggqi/Qr8XQva4sn0jYFY4HFsmD0S2yfMaQuXRS
JuOYjVDePOYCD9Eoio2iDjd7RApZi/gn+E9ooYdwznQVXD7YnTdm+fRvJY/jfeek4gey0dqVBxBj
72o0uK1uTNXQO30sDef3iKUO9pyJgdEhPPKatgsEqT5bIg9stxjGT5mGB3P7h0733NQBAFg+TrKX
u2FpBeUjTEEQ9jVivwk7pPRnTYtlDT49MqxKVDK49kJDc/ZJrRoJaOXOm3zfV38dlCfvrqanEOWC
uYr7lJU3UdHrCVHXoNJBR7kOT/UYlzq4mNOiq6kWarJZfmxF6zmoPCYWGQj1i2y59wKq93QFI94G
dgX+iYKDyDwyK4JAYxshlkzDcaj8LQslRtj/ifdUrnjiAgjMMI6RgYA3fl8Bkloejh6WdD/sHvHe
+o3LvF4CfTHrSAbXPcgNHawYze7riVev0KK+ky83Qe2KJ9ehck0ldOtrGW3XoEoLsL9/7chj6Vsa
a+TacSwtKArjrXtKRV9tq2jy9VMMmc7QyhZKqvlE5Nt/SWpvODpW1KpxJPFG6p/qcF3XyoBi+9Kc
hhwtCUPXkbYGO5L4mrQrc5MmZUdNB4TIs7OsWdZPnqMrkBu97xvGc3o+xxxegKMebNsmrYlInScj
SEk1JC1OU8VARwdx+BVN8hlgiOHmMIPYhNVemVKrUQ+UQx6BUQFq+WE+2qca8NuNSj6iIlLdCtt0
96Ep0k2CemSxyql5Gmoy7Pl5uBN46M4Zz9eFWkaHtxjZA32zLWK2IJJeF86baNP6sJ/IRp/rjOT+
sTFNwmlfM/CYncNC3nY1P7PNcuejz5BBx3VCRcil3h36RobQW98147XMZOuyOPads227Gb9+2hCE
NuXicCrRWSuIx2B3kq2+lMzYfIAY9cEDUY8dBwAspYlNtlxJWk8bRDb1GGGXyeWOltMs1Xm1A55A
JHc+G7qdkOLT4SBLCuVcNGwpXZKJ1I0VFJhiPIbN6xjzNewHIJ6BXvl3NCzioFig0EfF4WQSh+Hx
3WlrzyZIT2ymfciLAFVsO55VAGxAlP3kAPQ5rY7kzydogb2SPv38zOGUnej/rxTqBbkB8aOpR1e1
Cx+YQRjylmk7WfK2rFzoH8Mg1Sc6giz908e8cUtM4uUeqwL0bOUBe2t+8PS3dk/pIzrLHf2sEgvm
UIY4CVKrEV0Dg4wqEmCBNSXYxYbtHUP6dgy0lLjeISyGSwWg1MykFYrv9iw49aAvt8pJeRKI4M1H
7yUAOkwvIX1U6W5v0ZIn/548i3OvNkp3xSQGC9850R7NBvxGTLbWDK+gY1EPYBiynVlsfIZu8EoE
j6AmdmaSoyuojfTBpCVc5ZUBx5jDrmO5vET4VWrFPIuZZ1JcH5AR9iUp8qmvA/ANP9IMk+Z9T83I
OBZjPNeTz2+OJnAE4ZsQ/bhLaFfWFdeaTOdPawRDOgDxp2UNv7j8Y/SeDnIohh+p6ndqiswIHrv+
Hxv/on+JquWGeSUGsHjQzugHP4dQsH6WFHSzispovJvw/zt5eKQmdb7We+S/tjhZXNTK5+tzYkOV
dqAYgz648pj/pvHQJJy+u4ewsv4uT4miH+x+yv4Wl6T0ooWj2dST3HKOCYuyH3JaRvtaBEq6pnec
8DkFDevFoFS7cwHCMtsDLgflpifgBMjf5K5+1/YXsvrz0laR2zi7bosvDCfvE2XHXk6XXY2Sw38R
WoxifNFVHqqQcTEdHUr41VebZ1FYvn17MpcEvRov2fGUPX+v4c1yCa5cvFcrq+2x6xRrd8YUVgFC
HUOP+6Q4BBb8DcZVg37bEC5XNpr6apTOKyTUn/SntNU9uquSFwRwgIb3R9XXG58JtfiGnVMVY0vp
HWpTPIEwUiVpQMEtiWM5Fe1pjoc+STbBar3KtGuC+i7pYzefCbm66rh5yQvbNqQMw9M6BhNMKY6j
yAeFDq6/SCwuVyMzKOskEVC03Rg6Y8S3SbdbRSojvLMKyo5ffAS7IanrGtb54vKhmc4ywVX/oe7Y
co8vpNRj1+jcczIMan5J1RmHeo+o4xZtZQdpanfREdOOmeh1tSZjr5uPi2/lTvQglnAWjohYDzKU
XXak6Hm0vL/SIECxO82IxmS3aPAg4FFgthfckteRN/mzOJMPkOFbkx9ZADr6Tuw3U4E2hoQF/hZL
1k+DISt4rNYP49y5KHqPIPqmiE+Xz3YUMyL90PE3iof2Akhebjg348Y48znVQn3Tx4wP9ol4vlTS
vAwicXIseD1u6kTttSzwPuoAaJnqdw8PDPOBVYngvybYTT9Low6urebLhRFsqo9M8BgJeUe1laWK
cpb+kYwiYVQmpVtmTuQxeXz8XzJWMYR7pQzwbDlsRnirmKpEMNW3a6kOdhQSsBNGNxu8koi6a5ro
KA3rfW4zJwCKBEETl6SsYNu/SFxo6vLq4Wd3VRznQL6VSFj8meP8254s2Nfl+mP5kmbglEYQ42eU
YDbKRmnjhihwMwWPFcWxFBzwrEi76oJfXG4Fw12cXNfYbZBEaVCOx9w6B78r5czjFNcMosi/9bTK
wpNlFo6cqcUUWfJRERHaOmB+1L0EtmoJiOOfNibXq9JzGcLugmjqI3QudWOhosMC+z7MT1dUlff+
buAtVlhS1epH+WqLoTu/eeXuQnn5N4GTD+io/al21bWALXdfo0QK12iweOiJhzdGb4xwLzlDoIgt
XXZiGUtfmWAp/mBTNH1dfeXQ88/xY2LhUfQM/VqBX5CXpTC/DsvM50NKi0XSPW9Ut3Jc9mwfa+cW
g5FifMp623vwzPdsNjsOQsQ04tP4gFubD2xGkxB1jdNy75R5dc+Bjwv94CxH0yPQuj4Gu+QR0EF0
0xW7Z5Dd8Om3S2KQc++ARvnO5/S4lPZf8KtLeZLnbbL1BSm79IPAMQdwaxq296PrmR9edNSau+i/
rhbx2EmksGjaSgiaSGHLizCttxptur5r7xinqXKCypQ0Ny+fLc+Ikzt38VVg/4GSERmOBw5Xhxfg
gigq3zjXcY86eKZwcDMioALV4MFZ8slwLboRFKK6P4oaIetbC8tKKSGsCsdVeMJCcZT9WypSqEoK
p7DQVRp57JmGKDP59jIRg/KkY/Ho+5EZ0aGt7Skgv2pGBR1OapSjVKIUtl5i3QycRX6TnL5O0dFF
LeBP0wdY6Bfzq5p/ety30IlmP43wZWxOt0KYRwPkU3eeho8sgWK2DtuqxGCdaIKWToNBdDxGqmHF
wxRjG7j1ouTg2SUL6k63EIEwd0f1bgE68VKoi1p/CMeJQNBfzcHwC45TQM0FrAAKoJqVGb3ToIa4
BRQ2C2ZfxSYPsHFCMIl8rE8BcZ8lpJpdfBTLUeI9KXY/A/HAT4kgEbXmm+W+2gHRdAFjA9LPp6+Q
/UjMDyrQ72nR8Y9m3E+YKnvTXUBl0h2FiGceit2vzwg8APvDf6Yn+CrmNbghk338KTcyh9Zb/RNO
8dz9DbSIazupEFrEkbCxj8BcsRlNrTdEoQTlbLo8SNGIdwsQtqHiRFg4Gzs6BcXpOt1js/Df/i2f
AUBXddBtpBlltKOQ0Y5UK7LNPOhao+x6+nIZ0vynFINClc70u99Br7hGDCXv9p9YSTxJgtw6bnNw
c68Tp/LdCDO3rkyjj87z8aEdoNH01S4ok0lleDMtrRQFoVEfYyEeMIwH1DK3S5ZoieRGtxQaNwlR
Dpgn1eSulHxRlK76+FOy6Wo9OP8mLH2RzGCVxp211//ed52n93Ef/3YCASMQ+XDE3n3Dd4MnmBrf
pfAvE/1c62kt1p16/TYC3P9bSUZV8hGA4GaW0bkCgPqDFoNKdDKdgpPXG2opQ+ufEOfHtniDVHgT
IpUs6C1QgRRx9cqGlX86a+R4212XrT7kfcnDwLsnonGgD9YuG+W0omWCX0+2b3416r1MHzWCOAap
c4MLYqRh/VhKDJkdp7LttFwy0Hrqz6eB9wBKsl2cZiyRm4iEVffnMU4ov4/yBiUEEfNBzwLhuMff
3jyvYI01YN/IhSoKZCHFJObOd9IeRsSJc5CXv3qRQL8wpr0qQ/IqdvjGVQvc1vnXpPNt67+Bj7ai
AdjPpGTSDMq2L585vmCAr3xjWbbREuynZdRkzoS+jMXLAjR8mCbplFvwogDFE9YFMN3e74QuassH
oLLSlxktSY1ORgFDYPmqnxzEG/SPK1+pUsGxy7NzixhCHj94MbHColKyfmCQ5zKFafm9L5zm3Hvu
D+g2+uodLUWoFIeMJom+UA31raMP78+dwup+D5izgtgj12XcGYbV6Va0TWQw1IamECQ6h/x1H/py
UsKwagZtS6uxQwU5LxbBY0eO+OZ3IOdjrB6bGliVRSiKRxqITRDzlZiIRcfRhrTXZVZ8/sCxkNAf
h/66th3fQBsB+wSmUHVP8SBv0blbnFTiw+iF1qs6jRRM72akJU1DVCOW2cyvTfoJkQ7DilHxjJ1W
YVEw6Hqf99asPc79N4srmIxbsibpCPP0Vo4lIIQ+6F3ALowJ9Z5X3/RjMZV6wfBmnLptJeua2kKk
wu4VIKaglEzATD8wV7TiJ6LyVfAmCKQ2jcZ3EpcoUvZ3TNZmB3/iLynpaDmT8ivzmzNSM7wkSZW7
p6Sw3FTMBR4ISOWEMGH+Aqh89NOtPSi/tnYw5Vn4bjjB0pD5mThGFfpFwKVcmhWB7SwJvQ0UR03G
jaWqO03xHoJ4KMBztk5SbSb2wtKC7R7ct4LoLM0bp1x5D+eEVeoZAC3b5Dz9H1nySgJDg/iKDlO5
dHJKLPFD+Yev76j9lNeeYfBwCHbvgLNjP7enXKiXcuZbJV6fKc4agAJRKpHM8JI3cpr2J+CEquHJ
FVEEVbT2KMt54Xr5R8BKBb1CObuLp0q8RRm6hGgz+lXw+nEpPgrnNffV0EYiqV+v/gvsP9tm8pyq
xLf0zjhkAq6WwqUIqKIpt9Dl1NX1JbXQ34X+a6UwASPWouQ4kxbW3FQR5PF12+gboujbSQG0MRZx
UIXn/f8Ewp4V9Q1W7tN08x4HHq7OA9dVD0yIAVhFGZZUQ82VaTp4bv12IYky5iCnpLNOCWbrqiXP
0hM8W7td5On/vWQjjm0+jKGXxkIfRljaxl6zrZRL6MW17IoW87GtLi9y+qL+AnsHCdMWVTFja6eS
8h4s+CauuoVPW1Y/RU7CcwRv5APzgSIvoGd0WRV3CNOT3m/Mi/NXcbaprDomS5g8M5mDkGO97/WE
WMz9l9c/irwRy6Yt2PrEydEWxBpFR/ithezgnDvVPEwc3jJdooXgiAz1xmgC421tPkvzQk0bdjzh
2exVw/BGgH6OmD9DM0l+12U1HBUmNOUNe+FyaToFP26fNI28XipPmaau6gxhbL9QczkzZmX1wyb7
LijGVH5BHKXQGy1apDnGi04vnF1ueqtPM0IHmbXhN0dgJa9Un8Bf3ZxXEIVCJOcv+IM/veL84asC
Wmeby4PPIyd1isN6ihWMesa9s3LEwCZfXg0x3XvrToGAAy+B22jvD0V0qR66yBx4D0ryzlKfZAoh
MCj4Q/lIKB9AVMXxRentwh5hHKPr5lzsjD+bp5hOzZ2NFikLs+FcPWp92FFaM714PN0xUo3Z58yx
jTNGW2xg3doM3JSsUezL1abc5q3vp9tgbPunx1rg9zRyvcyT1Yn8SCzqgVqSCdmDurNSzCLj9XDh
2xkkJrJC6NYAVLAF0Qb+v67LPxzvCRO6znNbhqfRtsbzawMokqOQO8qd/YPD6aUQvMBrPMe9Nm8a
rbdMXPuJFSe8nFIDxZP4u3xe1nnC/fRX9+XrKUlmcdTJagjehaWA//9gwE1FQroqS6zpvL10OyIK
jasXj+IIJ+ryzWnj4R+Q8+xNHT/yWZqWvScPaTSS9Dzb+Ohconx+hm9nJSpD3ok0LUpYWP3E9VnK
EgkyEek8GS4Zn2Z3FnDMaOwlj3z0u/cWC8BVEd6PJfEjow4E19WKckBn5B7vK95nThZ9u8gqml9+
YqAKCHapD4NMq5uDuEv0nyJIMCHYHWSz3ebYAluvTcLBz7fdzNVj+atkZHHFu1+Ok2xILSXTphQG
xtsmuDPEclQ4bIwA9zLRfADywGWpEavfN61xMYOlqlGMn5FeptnjoDHwQg09IfIJ0ghp8NEHklzv
e7JgTHqHY1Su6kBpPRYIOzXwnGYm03774KOcCWPb1fBET4/ELo3PanVI+Yh5I1OEiJD6SkbunktR
80te9BE5xmYsbi4u1xBS+j4bshdGBlpx/2yzKKsyRR0oz0ETp59USpRKSDbTiR/MJcrHc0qRsXkU
oKlCWEitIM4O4jbGHndMUJmsTzl/sprKQcprjma3H6x1f4XZWUmOKdEynF9rPGAxHDynC8XssSay
ZbsKnu0Tq8gz/j1XkMkZ39Rs7y+gB0l+hPkyVZNPf2O0iEY26TENPPPk19VO24t72E1WCbCQCX54
nmngAG5/s2Mii21smI2npZjzKNBndbcAyq+FdWT5evojXbOmTKIyUCkqPJwKRYR5Aj3ppigE+v1c
DIcZHIeoNVgrc1IZkdVnvCcK4dUFSxIM2B0is5XKvc0W4oA8EAPHNYzlq9j/UEkikS3A2NCppcwj
6vHG8zjTUfxfVx2LUzpeP5EPrerCjb/L/EnhZS4C+kl97kTWolNkYdIYd158yhRUKT+QaQPSEP9F
ZpDEvRZRXC4QtbNlG+Viz2BljtX4cQL9t14V4HfvkhcX/BMVJal0d+KvflnnxHuOS5IBP7QbYG5g
S/ZIr65jPdXORoXkYkPGjEknrqQeUPklWCtPNy7HAJQ4E3ib61sr6JQyhJr3I7jPzGoRq5a2Zq8a
mV0XSTSAgATvYq9+dhYHijeVfGemO3SFreo9X9F0oPX82X/Ld9d+z1tUnuoRL16EyzkSOtHB9WmM
52gUv3WeeSw4/eflQQU4CVgbgTpJBX2NhabVo+nKAshMbadbtL47XUWlps/uogouPkX0+4vfWMyd
k104i5v7ryLtAl8M/3iW4oigpA2XFkt8Fte3hACSqqbZNDvnwMPVFivpasgnDQqNGV+wE9vI6GVD
fxX++hwZQmsX6OgNWaTqY0Dx20NFHiizbgC2AYIORYAPY5bH5o3fHjqsm2G2nzqF3+jFm7hgLoXk
xLwQcJgFuopbzxeBMMqGlva0lYWPjDBDphRNLlEJCmH66Zu6XEHtErbawSp/g1Csdxrt1klo+TrL
LCEoOI4jcdCHLoCKq3zFDpQFF5Q+Jm3mi4ErWUESs74MY1RzZi0+xc+T4sDxilfHZJvK5mM/z7Ga
+cMamHUwA6aBRa9ag+SMVweaVh4heTAsPUIfQO2ZWM55thJ/9PHUdaGS97I5TzzTgmQPhC0sE+nw
9erRZRdbr1pcuQFuxHWBhaNUORlH+aHL0hxarq65Qek8BT55acH5BNFdslnDQnIk1q07IxHuqGDj
+pIoRPwz8XQmMPhqFxvTCjOvu+ClQJyNj6ZRlBh+kILMqEbzrlmQHXdBHlI/KSzjEZUhDdqqM1hb
EGiKxYiAQl9eE9wIOj8Ksrh1B3lTyXI2g+NjFg9xNGdSqeIrRuZf8QEnw3asU2e0kr9EZUau4Hb1
xYichf/cM5Jr3nVJfkojdtjWhPC28/e8TWBeke8VIzwqOul1vAcWOcAfvvijJYstOpP35CAzwUJr
XGsUTW6EXkcQb0r9Vv5CX7F/4f/xKubvoyTgl34QHLhcJc9bJ7XXSdBzaBTYzC5JTkNmaIC59Y6d
YAlc3vKMZg48z6CiNLsbu7Iv8VoxFKGivFV+k96ak40MIFrn9FZl5AihB5H6dFtcxGKn8sPNxWJ6
FYjA7TAlmzrVXfcyHmVLRpm4d+Jz3mcGts0QR2VK/WgFXdYruo00/Vybh+H6kGVVR6TdySUusW/u
keNmMzb2617bKs7zDMBi8Wx1IlLB8wf5PLgdzowaCNQhesQ+f7J3quANPisT2+Q2+UToffx1i8Cz
p+R0miSj0zBgz0jCt6n7TJKbFBYzkLfx20K1FG4vfcGXRo5+rGRnRRLEOqHX/o8sVjGRwuYzK/HQ
PlUBKqN7OxjazPl96bmBnM6Y1kKYTF79xsm0LqxSmlnxfI7Za+qaYWPOzy+DqMVl+/iEvMdwgCWW
AyDgD6q7/oFide5XFPAkUzAGNt5qhKWsgEM6UiEzioSLBGjvwcsJ1fOg/YabVKEVIzZ8k8+Grkjw
zlq/8LPLeiWm7VwBxJpATxaTFMvxuZ0y7fGZhfhRcckhROOfAitI/EOlvvFNYm++unzN7RU72Oti
yjZBZwJzGJCSjmyZ+b4s5MEQX48rI/shz0vogYrNDt9Py1UiKmzep/iJt26eDvsa9J9tiNtyMlVn
GFqvypyzOJJtP1yeJLdYERhzkUEc7RPzFyGiO4SR3whrilGsC/1UFJ55QrsMUgfZQ7BVHS1BZnT2
gr2rEeMSvJI09Mazs8xPz4t6+NwF4bkWOo5chTL3BzzFL+pXoOfoel/1FfucFj/5CFvwV8a/csFN
U5uHF8xmNS8rTioDg91Mh8PKhpLlRzZxRdMZL7ByUnb94enUqYYVwiWQLDStAohOvTCUkLGMFT03
kMwPe6JMDgWuVI8Ys306NbSeU148+91q/az9O/x9S9iSicQ5cXEoFo6uiKq1YdjCXBuLie2vUTlj
3klngkEMVt/1T16QIz1Ghf2WMwbDrTyPogwjQxW0ESgdpSh8zn5OhgK/yEPhuuZiUUKu7mYiLnWI
QhJc4W0XgB67Ka5l4as4z53ocXX1u/k2xJ3gchYU/cV9mn3RPU7HIBYcnufVTyhx+meAOdKqHlVd
xTHuB58UL7vjNwIPmhfdPhhqE/rnLVJzbtS6+XpSS/mRgRFPLG9hMEc6+hKL1o1lMAIrvCMR/GbD
HFfo4lYDoEhtVv6x0QYU3fPx0Yxa6kPktiwqFsf2fXP4fdFvYQABOQSJ15CkiLMXAte9YF96VTqn
GnlBuXenBvSD+fKPkYbMQKscmW81t+d2D3NSBvTYNCALqGnT4AX4JZ+XDz/d/tG++C9S39sAR3mU
LJZuN/CCsUhCgd1+YYzKjtibpA3gKSwpkFD4CKGLu34Jj//ldrtqC0CaHPIjVBb2f0DDVKoisJl8
D3lgTV9bV8M7Qm/zYElHGWDQJzkyTW3GsKsqJtxvkkdwc9tLjJaRL+KNtK9Gbvx03CNYw0jEZpdy
oS7vW8jqj+QAHbo5D6nuUTM0WbdO3DARKmNwjoPjVGdtBB/2HdIkKarJZPl+KEvXtt3KX0qTWpex
hMKGx9NLnUbMrhgrf6cw/TEW1lSiaxhBeX9iPMioqcOgPgKorWdnQ0lsQjee/PJKjDoIynU33t0d
qrsxhEZ4DsCowQ5uJMlnS213fsrP0sVFITyHvGfiPfgvnCHumdCkoVQSj2cuIG+lmuN09vJp1H/a
0WfNITMHnhiaOAVoxAHKJOT4FM4rO0iUI8LEQKvZVSEjqTrKa5noFF0eN1lPNHbojEaVaZ303vu+
Y88mlWY621t8XHEQfs68DpOYDNbrLtICdEEv6yORukFZVjJbeF+mDyjbLAv7lUC5otRPJGqTZCtz
QD3+WelpwLRAsfaxLn6Cg7D9WQp1QOWrua2DbcCNYuERnJuGwuIbmmt5wEdD+Mr5bcf/OCQlVrfV
4FHAfS5V/QgPxczzKVXT7fUP95gaiVt7HUC3J/T1g8sEbz26bhqtL0WJcyzw4AH4rh8sLGMkEZTF
DlbZLGex+jJDCRxo8qZMGRfxu/AHRpf+O0kJSNI9v3acaXP59FckAsmQM1EpD9584kcxKzprPmXJ
W9cMKOhwtwvCxBofFYX+Nk+Ss6+MGu7XNhH4rVriVvNFvBDlFbu2/w/c6nfOQbbGuKM8d+Pi1E+G
k3YOVEdmSizP6oJGLsnIZxo5kb1wzD4NFa9mNsy8N39Y4qlyUMyCnm/k0kw+DOjGd9O7KMDhkw8h
328ytJFXc6Gwi/j35UVLIq6moU2BwFZFPMu8k2NJlkkNFOv2HGTgVqHJaDeSZayu+mZXiGAiak2V
sETUhF/HlMla0dWcvPziltjt28pyvaWdFRCEGQywQMpYsteJRh0IheEsA/Kwg6zTZESpoSM7wpiR
+5tORlO4L/jlyyNT2Ns/r7yPNFc4fhMuOgJqOrFDkNMLYPWlr7GYkmQql94WP2yGF3g5NBrJecKk
7LxWpIfJEXDPBr9DFvIzXm4zQZTCNcB/LG2g0bTOmW11Gz1sR6PT5dj9bgavpd1qev0il6OtUe7w
DMkWZpG2blhvR70kdEJ+JPJkHJdPH6/eNNmdSRu5E5NUM6d9OItxswv141izm9BbmFJBImdbnf4v
NYN5MemIXpScWA5lYd9FkA6b+zi/da/ZdkeFpgC9zAFJi6cHl4eqi3SDynwEhkb8Rqas0I3eY1U5
gwwBZSqVuRmYykEHzaKccEUDAqQPcmsoXtaETGVVpzbvoRQBbT/tp/jVSgqKXK352edS397B6SJS
sx4EfzxC3LeFSS02WXjfDHJhwxYJpkse0R+yNb4/Z/VM1nV7jpskNkKMGdNzW4s8/4jx6/oMVT4A
JsxH4I4NDd+oEpCzidWYE5sCTvvl4wAspVneX3cGJaxanbkDxavQ0NXAHbu+mlq2xfLexeBdYtte
pOoGrc5AxAtBosBiIlFpiv3bcKYeW96VkEGz05i6q1jKWVkdUG56++1rOMBzFQ+Sz/Rn6xPLZRfJ
ZU9DQH2F8Ctu992SWgH6GO5KozRXhvm/dIDsHKI33XJekxoQjcCaAGNn7+2dtJ0+QM37NRLhjs4H
fRoY2rq1z8zAG3hSeQyYVbdwbbLaX7QuuakheRo4DE7vTkKVEcMWkoyRgY+leToxVgigbTI6+F2G
zbeFxhyjpxM4XaEGy/muVNMGlqdGDe5ybPEll3wlKRFq1kQomAn3I7tHe2cAftJfOBUSOqbk0Gc9
+QEu71DCY1rM32TZZV7LSPAHuORV+7W+AzTlLYraovowVxDa/jgcYywFyNiv7XbsTqRi8Cmpuoq+
RYKD4CrjLTC0/r42ccMt5DeqcHXAqU8by3FmetdeGjHoC9um0Lg7jbGO7/FrF+15WDBYmePENk85
Qgq26xM0Bvoo2ePmC4zP/AFcbR7ZhXWyWL5Fp6VoyqTZrdCc+M7KQrOiCRJv62ANXA/D8NVmsDiM
cz4kU60fA5n6+0AmpJpp6IaHRY7hbMi0r/xfRPS1YTMqnxXK1iwLtVhqF8Ayhjq/0EY0Iwi+m5vs
HAiZjR+Zt5yW7H9DU3HI1tcrINO+D9rdxFk8OP5S/JJyMqYcWOoZhm5PQ62MPSyfuDPGmWFWn39f
GA8EVnwZZNDIbHiiEKxq/VYQEuXLmp8Em7svA5vMA0ijdSm6Lsjr1/fKe7U5fzNr1/hdTleoLmgg
qSv6+dnltFrhWkOKWwZcVD/FTglksdexrnOg358xW3oNwC8/NMJNNaM8PiG8Vk7V45gmRefGsX/W
swDhesJrmXu7draxTFhPjZQ5+ptj+gDhv5mCsQuEQQ2pxMRRax0uA3jUjfhdTRnk2x+Azs78DD/E
7gbi3xxQAJD89Vn+ltXJRlomclQ5ObXg8BcYALLtXTfmCCcHmNqOXRieImExDYWGTtcAO1q092Mw
uGnzsmjqySfyFJ8OEJROMLTBOtISy8lThYhDGVeDcbk/yqBhNogzmvas2cgAQNnCacbAwFwko6w8
GWISzBLGcJIB1SIRNIgkMq9P4f3nV5o06FbGPlOq9Ypsk60gOuBYGFKm9fVbLBUsLKpTfEq4rsJD
CsVY6vlxZC9Ohh8sYwA72FVmmUYJGAeI32O2ESsmhxML4lOhU4JY5S4ABybvaD1VvaFY0zd47nSQ
BFX/uv+llfsrG9xMb/LXi+Hj1+UJb0Ze4N1ZbBqm6czyrh+hBdxo4G52JHoZqVJ4i7pam63BLkC/
DXMAdcKUCMM+bzCfXuasqRAqEeWgWIO/BFQzWxNAOqgiN2dPuvzbaWW9BLFECw0Omm4poVX3bqZO
n0Ss7ovuaODNJpkQGZTRfHdGEiFNchrsj5Iqw/uyQYReyr1IJCBBuroJ7ubI9zGFsFWkW+bDnert
B91LOM0+SSkPiGj7WjZ770al/eBu+c4ddMPpGoBeYt5qEIh9uWHYCGDMg0pjD1KQDI/6KpKYBfJk
jMmHSu3mCNJIJCqm6EM0FhoY4bGAPYzP40mU4akopWa+qzFgC8CaWRokSJOhD3fCTsPVaKbU6eY9
+/IFUXHNs49gTsmOzycne6UvHDGVJeI5Z4nq51jlDSe7p8L686U/5E4v2v6CwJ7Z005+gyrkAilX
WMe9s5/2vcVhDHhBItDaN8XbnxdtoxrNYxJ1W8NdWywuDjJrNtyHsQgAnS09ndzktKKsMGmIaJ2j
QVfW1Fbe7Wfq1uRh2AwjhFVI4zFBpGoyP9TXwhMzEYsFopKN+Rr+riMZpnyyo/oOSqgU1g6o6LAv
x3hFzoqzHd4GLxJF5iY42Xr6FLprdrTcjuqyt5BaJScFATOZ/cHDDQlBzigT2g8WChko5avITRT6
dbQu8hpu52CKC1HkmaGKlvg7QTR2fACP6D9Thg8Wukno9OTclQytDLbJ9tStMwT74mh/Bhda/b2I
/xp+0/9uqhDOc3AIFZbHKPPWQpQugRk9jcms44a13W50G+4eA/XmqP09F/Wc3soI1AE3PqbliIVY
SzA0KJ20FFP+PSpWh0tk7ntQwucFN7S00y6MvxvRgUmyr2l5l0ebe5fGumINcDMw3tpdVPIN4Ir9
lPT4s9E8RoEy+I0mcLTR2bf2RKH0IPfftHi/64jAsKVT9+UFB0pmW0cQX2WtmihQd1k1mO87AhhV
Xu7mH5baK9nCLPdnZw/6mvHO31kue7DYXEJOOYP9ZJo7WC7YTJ03htIgrC0Kt3fTQjS/vH+8W9ij
vN50Sp77MjCM5I4Ujx6yVT5V2NCoIiflG/Us7Frp8wGxlYhPsM5LZbl/08i2s75AHAf66dDz6iyf
0maUP+RhiCxWaMxggjg0IDNq07mW+Mk5dnP0lJhp9W2P+XEuurCKgzaY7WAx4VOd42HYPuq/2n1K
Kbl0fXcH4dTljtmeCefsk6NmYdLPLiksWctSvMSaoHziUhnyp4s5gLpzwjhvYkpivhwd/27MvIja
SsOeV/fSFx4LUejSsbnpPzSVM9MoQGcrXHLPMRME3RA5n7GI0mVMZpUjBQ9246QVWFOQK+o84NC7
Y6FLx7vJKoJOUy/XcpBDSA9ZRHKOiJTeFMFMA/NZR8aoTwbkOaLwIrk+GDzUxHt9Cx1imc0h9bgG
yeW1KOD0F97j+qudDImV6z0KZJcutx8fa00PWmqYe9nmc33kkePsZDtjufdjkp+DoXr2ppr6f049
F1CAj01Mk0kSPCDgr82gBoh7zbzExEUZScn6mAymp+mYGAM98bkv9ELg3aJBNxFGFU7X7oSb44rq
GwktUnPlq6vIVdtiemnC2Ct3fGlvSBPFA/1JpIOkRIooSQvFzyeZY5u3trvDNOKuTz6Pm9wS1shq
QsroU9j27OdbTGZukXHcDp45uuzWrpAdxJQ+hA0fSdlCECf6F/HGZRpAdU1LU8iOib0FWw2mBqFG
iUd7+lI4xIx1ramOlMgvAoSVPXJoNQx9PBjk+iGXtrDH668sGtzwoDyI/bNvoS5mS9n4ZDTUcgvq
O3TW1aG2RPQzqa5pKxKGr22MJuts9Lb2ZJG7H+MHRMEN19B7HZj898cubXc6QAye0A42cglS0ud0
LY/Micx1Hj53qKNlS3r3QCra6DDXW34+4Xqbd7J9sn4nGqRlOVMZRYMhKvrJ/gHni3fihEHz11vn
cbPejWLI2BFyCsDj6KDVVs7nrdGXBQiCge48stlA0PCkNV5GAb6JlIob1barM3qNjDlyiuhPK3G4
Vd+RGMkEZyHbF2794pY/mFMCVCBarPKL6cStee/0bISl0fZppELsnpuH5ZBw7WoqCED/MsO0c/no
4xSVnfQ9WqladxipqiZO25OW8jOXUv6n0RNsoB7CflQJ/jPiM61Z0tSW36p8pCD0GokiNVTJvGIz
k8lcKeHod3vbLP54ku4wI8sljUI8kg9M3lxz6IKtii4Vr0Xj3JN50AHRxbWQOpNs5sL/QMCbUatR
EjYeYHXSEVlsf32aPLVcJH804YHH73QmSxxHeD881Ae0ZaCrZEWN2muigYDbViYxANZQNdTgkrIe
FZq/kPZuGHi16NpmDJxNMi7cEmX1XiFTqluXzVxGEhA3OJv180RXsprF9108bBBwTkxS3LQEap7e
6BVtQuGzu3/cdY/f6khQGgNNpSuxaaPwv8IVJ9iGfQSzFzmJvkpFN5sO0OQYpPFj/bIay8kAVjmE
d87xpclmxHr4cDSx5ZquMk04qBibO9wCbfazLbdxNvqFAdcQAb7sojkBO1pUXeFXRoy5UyCuLUsc
S6eggHZW8brzG+1wagG+MENbXQwsu0BAP6UYRmXI8wMOBmfO8LJ1c/3ZG4h3fC8nK0uEcrVT/eZn
dlg/hMLulFGNziUvX0rf8y91SFd2DRTAQL4OA4tTCEprbCkyX0qTyDPUAw3ocF2r5RBz3ATqpm1Y
aT89cSbID1/z1Eii9NUEdiSw6rZRSxIruG4NTz8nEiXfTg+GfiIYn1tg3zzO8quk3Xj+3PCe/JKj
V7FYAy03Efnsv8nk+26bztEzLQFb8ErlFpXl4XWOB6NMkSXYkhvC0nRfoI5D7VEvl/yxdrt3KQUQ
7yTG++JMhu/IoBndveDIVFR/X4ArdadRQgsrDXNvoVAQyHxPDKOYkmnui3rZlv/jTEtAaJlx5PcD
fXdO/2nE8YymEY/QxhmL5Rb/Ng1xAe+Cfc9FE0qa7klNmwVoWV0hAUvsX0Q8UABrJCjDdHKKncmV
mL8g8zCwikV1543mk+jbO+gooPnapj9YaQ5IU46VLEZhVbGh0jGIq5jU78HVy2mPUWb+zRla87Gi
foL5J/Qb+Z48pPg9q40XYDVo89ULV/kUpwCvQtWPntFPBgzitbZbiYmDzfbsewJY11j68VsHiN5k
E/FbjfNMn0CAF8c/K0Z2oTYDis8O/qf+yc9NRkPBtM0bjDcdvX7bXe7fjWoZfxGs5zLa0KDt2Ijp
7ojm3XUhrEJCzjDbX9BMmYD21rP8Fkuon/FcLH+Q14No7uHl+1nr/yEp6HtTFmCKT4QaFd90yhdD
3zUGWHLnYRFCqE5Lvve01T9rMtSeKjZy6K/IokwuUMp04ikNg6KSMErCDWXylvCWUJe55vqVEJlu
LGH5QXQiNM6S+inIeMgd6yZQCyjZ9BnXfTdc6Z5iG02Df9v3vptfLwIboMGx/OUk2kcWLKRX/wJW
wEzsRmiXUoovgf7x3Ea3j+yxXuoTePmCN5Nx/lPQFsit+Kt1fbO+w9DJNKBCX6gttchfo1ALsD/f
c9sxDDt67Z5ScWlCCerx1hDXeqnjTktYaekM8N9irzhDyiOEj3svpHZwh4ZxCVKJDlvc5qpP6ioc
cV3ID7R5XH5PswAX7SUXkgL0wh6SOWOlOd9rwbP4DArC2KvHQGyzLbuMqrbe0ihoUFQiMXMVh4H4
5D7mRSBHNhRLleV4mVmIgXZMGVejhhOJx+3WjkE6IPIg6u0QLWzkCbV5HvIcbuSg6MP4KgeS0OLP
NFx+D5cMnW2ytxqCYDSnzoN7S5od0OWqBzpG87DEf0BukscAzSzQplXz6YCoNBTMGnpFpnuht0pi
jyFWPJ66UM04F0crYZSiHZHf3KKkMu+pRuaxE4SqkXvuHCpBQmyxlh2/yjdcLQphhrS02Aai6wVk
Do0TRnh+g0xR5d+IMW7W9W3f70AOT3v4uHkRew2/l6Kg8NKDWqyLQ4yEo9vRRl5xewu9ylHJnAeC
JKFEzupR9MvL7I4/bjXIInMfwbpRTsdJrmZr6p6GuaXMMTG5NYwwMVe+ix6xb8xejWHz+YJiiv9a
L3/6cxVaP8aic5P9dZpKlLUqE44cruYjAIVJh9+66MOkMCZZzG/4UTPPaMRXJpLT/k5QJuXQl6B4
mugxXDq00+oTfr7g1f5uuAsz31Rej0hN5BefjMCgv7JSq/i8xx/Ghb22tap+hmh1sCGxGzMESeEB
r86rzDG45hQ9yFTC4FH9uCC9yyJAYI/XSkyr9cEzUUFDyf+JEQtUjfHbWHhtc2ukJaTtEBGOwXtM
9mGFouyGiRI4d+RQ3LMkhx6PEISKWvRMU3rWIkx1QZOjFNgAFhpEBJJcSBoM3YFzHdv3BbymuI5M
oDWWffH0JLaw3YaFXNypQ5aKpZWBoNVEBP6fzBua2IcVD0vZ0oOGVBqIq4/GQVRltwyzaZfwOnZ4
0nqTugCSq1B1GoheCZPr++zzYkhzJU9PPVuUi4dZsJihLyPIwFzWA3yLr9B8PxtS+jyrWz4IEVCf
A0Ew5uTkxPANIDi1S6HFVc56vpchaewMi3ZeNl/lB20g9JxueRTY9Khg39UZkWYDYwhzYvZ3npIf
JLSwKvpZWF4yftq2aEerckvBqx908qrZyeZyY9Woq03Rn6En+cSwTfmzwedAjsBcSgbStKDzTutY
jjqZi2a8d+4IhzoO+Kyv6Bd8Gv3lZHGVGuqNjJEP1aD0Zh0iIDxGfz+bEeuXApHpAKqhG3As+Yer
0XRquqc7AV6hI7CK2VXiE/nyZ0xm3aXjtsBd1oi3/6p1LMAV+EKCVAFQ/jMCKhlGtWrxiyM1hiRm
jah+i9pU/IdcshXlNySgQstPsBzqm6rlc9J2XpMSpOX2IBiCZOzHdsYMjiKHLSop1B+95jjDep6W
AwXjfMhrN/Z/ZqgpKdU61ovSUYicj95Yi6DuBAbm1vCWhgckWJJ9nJb5laSKRznU4Wd2gxA4m0r1
EUEbhiNp/98JTBPpNDxiBlWIVzEXZfXXZpbOLFY00AOhu0TH70lN+UoPW3+ni+CblzX7xeEMpE8i
hOwaGdrvxNRqmA5zUfVzy5krm1uAMOcBcdoJH/ThOdB5EnNcqxLPjhdQdvIm+hE/odzXVxxox79A
qgvSPkqeTg689Huye7gwLhn2PAdZgBjdKwiFeCSVivh4K3RcmLeZiuoSvzV0w9P7FG0bJhHenM0a
Ao2FFDcdqLdmQMlQ+KnhCm/TEunAlr0lkVrdkm4HPjDzbsFL0K8dxFoc1SDh+xfzt/D1VbqG0UNa
dY9QIF4efT/MJVUsTnFGHtQz7nVwrW9KYhqFkS/GGaLfyNNL82IdJJhPMqfyJRa5S4egru8dMuAM
x2l4OYkE5SCLQr+0ZCbwBd770tMD+FAhiOlDRFAyg+rUBhtdkorqz65dASQFseky92vCC/dzri8Y
dSNnGIqKlo9mPdFE9Sjevj74DsNKcX9maftLN2ME5sx8fAFxeWbfMWqLKyR8BASpBXJkC/VzKVJk
k/LGAFKhDorMmeviToJSezBy3jgOwURyTCe/X5G6gid/dV1jtAPUaEYygZiK4HM1Y+RimjCU4ExF
PL1mZDU4U1YgCBxrQYUm7o6q1t/+HgJWn1DdhclZNur73mjzZ0vqZlH7tfyGo44xP7t8k9oaeLI8
7hWl3obcOlElFcQMJN2Zruj+x6ZGFdTNhUTiBtCzz9xW7/pzpXMMp6OqoPVEXZS9PNHhAbRmv6V0
NXRiXbV6MZaFc50CjdPtfyYmcwFbyM4iZrhFw1fhKQSda4jvl5G4riuhMvYY0YleJFf+TULMtA/h
m0E2TX2csLkLSHA7JXoU9q4EY0hGizHdp0UMUVLXe9DlRIYlVW3r3pbSjkLhpPSaVn9JWr4fq+ti
B/4ou8KXsJfEe3vN1PnsFlHkdeWlu4xwdMpdjrbycF9ThXn1utqrO0dizByLVuYJ5Qm/uQJ75c2V
/3goNhlNc77cjJa+eYOATn5BJZjOPYWV75EsIqjELuIPwrb3NyCLyNjLRuJYb0o9e4/GGBGDYFQu
EQ03g/hMCOlSASNQtNq+CgJWDxiwUgy7FCdIrPVK+NDpkUOZStw4lJtBkSdw5VJTJzZrhLmFKBd0
fAZny6E0FQWjDQjkZvhx9LKDMiM1vDfUE404XPkISPU8oWyN0X9LRxzHWWmWlhPTtjzyAWTQWFED
TK5naua/Hvn7MTyQ36i1h2b81EkaEqLBE4sIdsDSLq+Gw4jatxQMuUCxi6EkqzeAxVHzKD8yRffz
rX7VFp5K62t+y1h0DZrMxUnM7x0IGQSgD/CySZTOcAJrd282F4LWtNYJqxONHwFVu3JLjc5XWw77
xQWMCK5n6oh1sHDS0vzSPCEpHEInuBPkKmnsXGjrnZIp9RK9SnMKqoJE28J23opkBtEbcAEtS3ps
WIogogFDyahaUNoHovctDS/AyqvfcLuCwprHYkfX0sWmXKF//pnPrBFkSNzcIm+H+QuUUU+Ka1fi
j0A2HCg58CzuUUN5poyZ8H1THysmpGWjx9BnGym+rJTUaw2SIF5ERL7phdaYAjNO9GbC/rpu8Leq
9D4i4QXKoSDkeCj6Qxu8PNWipfdvMX2D2O73F5FBwhI7tjR9rFJ6t9FBp3Io07aKdX7vkRdq38od
/uBzI7O/LH/RIEjorFEU3KexjB+Nf/KeKHHei7pHtfHpZcg8kXXP/GJIMqwQagOnJ8iYfHvgf3HD
3NQPNcacOmXMxaQPDySKiaAXcMzyIzzSS0FVAxeFwJhAYH2j72nmokFcALjzXTVH3szTbd5SmYWr
mFxc9J9JxFZxf+vFfy/kFuNXD41jm1qvzzr+ZdlgMbg0v9/uIdBU0eLhAf3e/6uPmzD0Vxmg+iHv
UU3atR0K8ETXdVs/gDlJkwbkog4UdGo5Fr2XERFC1RW300VBbPiKDhqHdtJ0/GQqlJ7SKFFQEgRn
Uv7CawfPGn1PnIceh0UFb/S/wtJZQnzoMdGjznbCgbUrpz9Qvr8RTPUI8tM+QZtSlgXvo669pJhC
lk7+Cb3DEze4gNqlw9JVKqxU013BQW8L6i4CQDsJ0nstdFsZ4eO0ww6JOPl0Cu8pMsQx2ACB5RFy
lDvDJ4ua+bx1cuwMnyg/jq/oe18hOTyl1g3oB03CjFcf245Db79HVEULhqq+y/vsrq2csuW7IHBV
Sk+YjUGSo92cKUlH665CJk5RR7yJsb6GGMuVRh1JT4LCIZaUWJCwFaEa/6dByExWynt/HJ/E49LU
YPlt7jdwG9V4Mb+4iuKeUkX7Ab/EjOg2LB1ugalXcaBBwHs9x32ijjT6bczv64QbxXW9nXdnMD77
v8LvIp45PdlQcg4kq1IWQlDfrrcptyXmQkyYlD6agiwOnQq3cWG0fbEXw3l9TIdAHm7u1i+dBaCV
li3v1FrLRNII1nZ0yZ4TqukjnnGn6s73u0773zb3SaMJ5cSK4THkKK1uLe8Nd8djA4g9zHhTfYiG
UxZ2U8nIxFLHnYZeJCiYhh7avepuIaZue4pQUdaEqHXhLULiY6Lzy8m9pZZ2+Ww+C9nDaVAB5f5m
XLs/SY8vn9DnexdKmOpt1ZAJxC6Y0OAja3I4klHjpykejoZyinLDkP6pvTzt6IuyQLf3LEEIYbkG
Xk12w/U+f/nWuwpIxOPWNkLe2pZnd5+B3Alukuc+3JXYgqcN/ZgL9Kdo9s+rlr6FtAunOhpdVVcY
GMOU5ScCuO/fD+eRvG8uHJrNBvOwsqOGjFVgCVUMLMFeee724B2OUWHFIrLG0MpfDDZlrB4xzuwG
PWhrUvZqLz/J5FGwV4fuNbJhU2ceYfvS+yhBPZGEuOx4vfEMUWY/cPD0SHx15ypkOVBkDlmXR0mo
eXZILsbv7I4NIiM2ThTCLxEdqo6H9dD+JujrI+PoKXX0J8JnhXAqCv520DsVHh4tpnWx3lj7czy7
zrlZQ+8Ukp7o1V0T7JS/4iAV3AX6lVRAjuBYHZm3jcbXPffPlj1FRxdC8O5gtKWc6rW//WM/Hqrc
vTzNqOvWPLNrX5yLc9Zo40myza+xIUmMMc58DTHngxMWiqo/dTI6VSAR4SYyFwUDMbk9ULsEmFBO
IHJ0clxdApy5d5RZWGDNtQ0TCR8DGgTvc1IfnI5AQuV2M6JmjvuYVwBNNoyjYRtR+dTfXUtKZnsP
XXQrGI1mCWBFQm6127tg37XiiZSq+Xuvv4Nda2oqQsTmL4aWv6g4DoApuyMapfDoe4EcXfZa5heE
43EKE/PjA37wmefzjY0osYJl/67QDr/obAgiaAj6kp5yfmSUZc3zmg+SxNJa9GLT+7+jqaLysvo/
+skD+vaYjUBXgjoWYKzynDYASLO615w/43h1hmOzxYZR5RYSh/rXocZ2dnaee+vIU2GmjdzBEy6q
Nx2Xwc8SHxyezwb43dSGFu22/ugxO3Ijn9xbS/UYOjTvNnlYE+6osn/Y7wM7SPk/3oIhHdus5T+n
+YDpM9naRrm6F1CMa/02d0wDq5MHzmKJHTON2et6GbRwXUeKVLzk9dv/xlIg9JvvTAM1ajtfmMdv
HZoJ2HQ7XA7hYFV3lHYXuYYajU55dND1Z2Zh3g4qZVqJU1TzZZJIqFRup/NUaFOpJUgF/qlvYgOc
eM87TRcLa6VixACpXZ7wzPYgu28NybvQnMD9Up7g/iGeXCyA4CuIAH5JBMVZ+VoKGi53RwBGquH8
YauowebKM11GYSuCqWBLw7dR7VWJcuwuxAFaNbSU6T1ZckWvlqw8RNH9sdNHvjUI1BpbfzRx3EYq
qky4HUzPesN6zv8qAXJHlg8Ilj/vDCwdHDZ7sSltaANKX3l6PX29WDTeob7PP9Ag1Q2bwUp9cTVo
cr0pcd4i0b6OXjZSv+jN1AiWJDe6E3w4A99xE5rDaXtk27A6IoQOMNINr4+UndOVwrPg/e5Y/7cd
gCZTf4Se0r0x+R4pP0kDC8faQLQIpWcRggcLUZZXIg2R1Q+PS7/2+J6w7H1RV6J0iJcVSukoy8X+
PacCFuPLfgOoNmi2m8i4qtDpCIkjxO+4jZEfHfho7szivJjY0hL4ZNjtvlAV3YzpAQfYApWJaIkX
iGfEbMLfLaaSEoWp18+Z4Bj0qbHwrl5n4UcIbxHhPC/kh3AxA5Ca8F89BMIsdE5n0sBDK95P59Up
omPg6iJwcoVrrepgFeMIzG/4F5sci0aFd6pbqoRmhDmaJghviM/FN7VLIJqv/hf7u6I450eopT3r
VjUqqsrU113eZvk6XbctXexDZRL5DI5YJZ6ZSDz937oE+B7dYCROROa9i3A4REHbfZTELHSTRr6u
NCiHBnW4k3ww1HkMak3NG/Z/RBhcxAiDMk4Mp9oqklRNyCeNXfwb0nGptlvtTj2U+Z77SQr32uXM
OE+3Ok3TXi8wmfeM6e2KOlM+UORw7dDfF0hZpK1CogX38rs4khSGqc7lJweqHxsWz/KfJkvvhh+B
ZSoxOhmeBdU8aHKUM+W5lQHWvLXaIuew4SzI/tlNCtZpWok9v3I0aYQixDnN7L4liYqU/IThzZL2
xuCm41Cohofu1g+sMgnvtzW9xH39Xy22aNrnSW5EoMR7PzQKTwOC65rXbpfvysh03HHVeoE1t5lH
6Qcqhwp6cmftVrnh5rJU0VwkKTjiczd/YUPPmgvEkWeIXwBJSwqEb8g0Ix4qvJ3dLWQoNWl4Emr8
dKErwLhZkgMlLuC8MFruqNz2kLSJmL9PlBH5twnEcRXM82/wnJ7mREJ5kmPO0aGMlFePHFgfanGt
fjHueM0I+9nDiAGlPPRgKkLNbQXpUiVbDc7bc0nH1yklplFjEuOFvi/xPn9At0FE1rDV8MHQhhEY
Id58O0LdUIAqCCeoyVt5pD4S9W+dOOkUWLjBSNbRFu8m/BJ+PdTjijydKN0Yhol8OSb8wBlR3BIK
c9g65Ysq5jZ3V6ghW5O5xZ+NfD6t3vEnlbUcmcJP77BtziK9Lm8g51WMO7ylR7i1Y2jWRNZEHUi8
lLbChGdtdTINzsH4nI7hk8g804lZZPv/dVfuZLjTHlJIXNmV0UhwoCSNzhcEK1oQOE510n9B++U/
el00+pWp4CjkgXBeOXVyWdkSURVLAHmxqsLisy1PiIW2R0iSJYUZcexhoFplN2o3rVyk8oUI4OYx
ZXcrLZc3brzDMgr0LukLAnRny9xoA/TVNWn8sqky4rSXj1qj0QSLJQAvmdzI8N/d9oo7xoQdwHGk
s2OrDVk4X4Woi3/cH2SqPXPCEBCR8pjFK4Pw5dBv4p31RVOy7AH168aStx2N79KC4f+jMkYNJZ44
GacINoEBwtES+COxPEGqdkW8RxFHY6/19W5snlIBLyiKYaO9B5MyR1RC1ivUOdyE02CopiuZ2gNM
xR2kTCQ7zP/FcM0iJ/l+MquokaD5F142gVmyUywzJ1EoRQccHvdo3qGjBceJgiE0llGDdw5UcUQp
Du3wOjM5ojbGPmjWVu1/EvppeaZ4yxyJBw4Ti49UKxLHKkyMcb8q9yhcEgHsBjuQuCgblgTKORRY
X//xavSxyveePq2s0brZ35ouLGhq0AzPMPYrqzIIgXcM1s0Iflsqk/yBpZEJxLcu3iAbS81qFq67
39ZgrWKnYRioZwkYpxH78GssTyVVBc2Immd5syzl7K8RMJm/uqOeThak5SepsnCo5N7YJbV0C6ol
+MN8sQjnA3xBfdrJPjL0DdyRgkKnuzLq2hGNdjyhawbWcO05OHl9/I64m9odcXhcxVE6t20QSvFH
WwmCKHO0/0zJvaHvEctSBN2UHHj1x+Y5BLeB7ilE9a7cdgTAmCI+djAZEKtmcwTT9NDzo0nn3zhK
WeSAppcgJ9zZMlUvK3RJ9MIAlLO1/CIMvu3+7PUeTxQQ4RfbCbjPVpFJwT3uQR6C40Em8KuEPMuV
W5XRjA2eK+n8zIgv7+AJdOO2oyuEU0cgm6m3OnqSSmZv3CI3h+Qn0yQ14eF3wLPmhzvuVkKmovMA
73vPFN0LIniRfvo5/Hm+u8Nb/6AmlQCNU9Q/oaXqqXxbjCSVaVD4irxusbz1Iavid8l/TJjNqICN
wpvBwyrdCS7tU3rbaoVp0DgpQ/eL9sLMD56xolbHcrGYsF8yC5wV+Ls+0eF0n2LiTUE/Ti0R8+9W
jadtmJJu4OZTofjESzg21DFap2RfFqxBwCIbl3JyeyFXaua8rAhdCD+lGf1LGsVV9f+uVpBodXhW
xuZtezwQVxMPlr0Gvl8qmc7IUO8L13kXCB9/Sr4DTz3IjeWZYYpKZ/wNXOfK19VCnhmRyqzV//KH
0MBC0+hn1B/rl46b/giGlK4+u+ek8xEv5E0iAVbrRoPgI0mSx1TfrH7Xjwu0VycKv+d0jG8D4Zcl
ytom1Aoa9VFm40ICwYpmsi8Wl2ZEhiyPzDeFRSUpFrY4tjtuEOLkIY4Sl6df2L1ApmE8/gaYSzCs
3bhHu/EC5MCJpnyjcdo2NFkeTYLuZJs6ypCwHWhGWJ26grxMxrcBfXgXD8odAwP5nUHyc4cViHE+
lHyYxy+wv1XAQ/mTmM375fLcHg+UgpVtIc2TZWMn1jCpISvQ7Hf2fxwhEwvL/vuZNzEH6pax48H+
/xPKui0xS6ovIuWsZEcPYEnwm8Bz15VGt+Uy0Hnfvd8NmAwcVvBDDEAaluRPv7dPEripcNvormHv
yPNx4fT97scDBcbhZiMXWuVBmgKHHaCDdXaoIagX4c3YSpo1NNakCoz9ur/1OdWfrPSsP+t0oau/
TDkM04G1YqNAh/sUcCx9n1u5XVQYRq2fmbEKxKFdOdmrZR7kZpWMCf+FTArRy6khVXgzzzNxcCPc
4HnMtbh9j0twF4XpphfrtonkAaY79nkBcUtf+xby+yqYQ1NcrhUURM00pb0NT6N6YxiVLcuVUh+2
kxuGurPQxWO8/ciFyKJROzw+dd9MukGls3YZEXTZ2c2G+Ogk6DonlfTkMf7NVaqTpSjjLjBMjLmE
iX51J1Y5HVBivx+ce2os80iSnBu0GT6dJevd3ATbh8iSEY7NzTS5oZP3mytGD+zqsVOmjiUxl/6W
ANUa5r9ZKcTHetlNejkNabHm+lIKupPizdIutlDAuHzsnvR5XGSBKInY4bSqMsblc0UvzPNQ63w5
VUMQeZhzR711FKx2XYsoab62UJ34CftA3mRHj6504znfszk0WuvEMBz396f5lNV80oN16AOIoQqp
fcgM5FMN36Nu6crSqocDSIuvZ6snvGFAbPNpE4iGQUNg+9fOzaCOsio4M8DIR5DIFDi84CdZlcSX
PJL5LZZ4JDLWH0mBDXgxXYDsUkg/FU2oc6RKCI7Gqb0TY5Nz/KU1uPNgxZlvrEjl3RCBsotCX35q
8uzr3VBj2bOpRDyHlmn7BuORC54N00Nuk/PaWkfSdVUodK4GSTeEsa9qR0To8xRm+7tkL170Bv7r
cgWUjX9YsIHsJ4Hsifgt8rbCSigbSXJV876MjwP4HF0ogpQseYFs7X159Ynq1tS8XwT+5LcuYemO
iiA0SmJbhQhQytU4Av4xuH+SlMzEj96r9fvFxW6ajhP3Py3KGWphdPhCGec/RjU00Rrg3qQ7ovbf
HGu4+2GQP9mL6fkUVw3jGBCzOQKobrJa45TRVkP438Xwk+Sd4UX8nCZNOxw8sneEr4Xy/Z5Pv7CE
/94sDiYpwrB4HlXGD85WUNK0XOgilWAYYtHR2yyZ8xS/5+T7X58zlF/miV8NnMgDJIv8xlBcZ2Ri
25PhfgJKtb0YHM2vJJXOH+W72yxHTVcwuGMoAjbfI0isHuw0EPXzlSbKEZnLbiUsKB2OX3wiiJBv
JlrAXJ2qzFq3QYw+SHnhPBLG4NIhRyMgsUY53Ne/c2oqowVj3Fqkob/JzUdEj/SSjvGMuruPxnTX
7OUC0bOijP+LMd19fJvrbbEg4yp44mELSAYFX8uDZzeHrLOC5GBifyzU3YdQaFKWNOJNXTO3lHuN
BwvEe5TiPjmTydzX5tNoJlj3zlATxgK/AwYAa30ciZTUJKfVO+Gp/V3J0s5VKBFwvvja5DJy+7M+
qDKXl/Tt3GSnn8XWwa7RD6IvJMdJNuSWsKeyd2PVWxjx+c9He6/Rsu72ePsxSXzt1362XRlVQ0RT
fKQjuxog9HRu1anJ3L5oshBSZ5/pXsMP3yLsQJH4DbwN/Z6Vur1/KhnLuoo7GiPTc4waW5d+wPJV
ozFufGKJdMki8waP24ugs2/OrrOStiz6GRUMPuGfHodH5CbmqJndOPQF2hFtKWEynn7ysXwMPOBW
XqB7QSgexaQ8nm8gK+lWt2n3dg1GdLBXMHcM7/eujMVahxTU2lfKjrcI8+vchHmh7rRWRmk3A8hh
8womEk1IKiiHeqpvbxRY61ep2FIX+P97o47rBP42h+IQaaG8xZfVSfXDJAYC9YDpwiWzEaGGWzFY
DHQ6CsrugrvO39S2Ao5zAmeMIy9tng/+0PLK8kNYZ0YrF2bf2EIn/85vufzyvriQYqpb/Gv3McZO
1Q4twFRBxszuVRxh+CYEu6iF/tcGIqDwdR2hEqr3zbHzOKN8KGpWUgZsIicDHL/C099nuf8bjLP6
JpY8Z0kyMqFYkAkRqhpJtGm2CEPb+YNUi5Q2kKW4mSgc/V0+OBPImalDZbR56ZBba5xb7pJ5gJVF
rzyiImtDBfUoqOp+iwcjItb0sg0sw31zK7VMo8S8Do3/SmmYLB428qCdOYpln5fvvcH+S4ff5xki
vt16/3vcknQnowgKl79Iq8vbawxrrYoJEH9noPPqUHxFCMlM643SzhapcPnEMMKq+NYsKUsrX3Ci
/xhcVxukBjjvnxDZBwrAbNXmF9hmbjq1pG96M7HYzlosm5NsNEtWgVgSzVm9Wx9cy2/chpT+wEws
1PmOBlVlcQhbPhGd3S+6W2btPDUu77ZLWdQkL9VnJa7AdR6Uyj1kQFfTdgy9ua56uI5ocPdHYr9i
ZDHw685YU4wguRVjjtH3+SkdiaEVbJ0sMZhsmN8k6Zk3fh1XslKlKEAAXQMyzZtJDaG7QxlRhpL5
DFlkL5oUJ4zpzw0LCB7gktjJYxWJWKFAzl61PsoCV+Re5YCwvKf19Z8wkSfFyH+Zox0u3f1scj9E
HR1l6jrX0CXgNGnCTFQwGUoFqCHzDFcVbJTjxLZh411XZpQJWdgg7j50q7D46xqx3Zg0WOxKxS8P
g1yiZnDhQi0syPjrPNHVUY1KRhum+R7yiZCMBVS+No8SypQFIXjiCggeBzoRkp5RKbN2oMitWpVh
dSv7Ew3W/Hu+3NL8cmCaib2EfYCgZb1k3GsnS/sen7Amg8P2mHynInbAABFwP4vyvLwFPg3twyAN
Uu/SCXpBHqm7ne3wuxo7OfNGmngqVy5THnMl0XrAQJN4fz25/BJ7UULznyCfJ1NbLFTfyKFlz+zS
G4wT7QRcHR/5Hle8g1S755+0mJfmTV2MvuaL+yQdkQbd3267vjvXUtnmQDs3W6Y7oIRNJffMiHSq
6u6S2fjY7d+w0+jlr4b9ajEkR2aBtWDsGeLSHP9xr8Zmj90hnGj4Dq1rXVxGBL+BuvTnhrv9NqqI
6G3Kf7XVieVG/6SOwTOV08z0uxHAgiMmWiaq5JBsc5pbsnfWdC6GEMjUKUnj4cmuUXejCQqQvnU+
loTBwD/AOe7YpUk259dggCUVlqwIhXMsXk5XNnuSdudUt1kDB+0HEM87RBXXIIv1WemR+b0vtMYd
Ok7xXL41s8c8iaChh+ATShx0Y0xoTREOamNL7PFE3ufweUNoPJ5NgXyPpbSRYl4c8T1EQ2KoUPCW
WW5n9OQsiLjn9sjldU+GhEHFUVVQ7Zkt8s1gn+CchxYdQHxoyx5l33/McbBiFnRdCzzQCENU/Asf
Ql0U1Ef2lHhjvt+0Rr6+qUAbhu9B7H2g8yZfXvSseL6TQdShzbjXzaq0Bv+sKE4QpPQgngtncgLq
PZRBrk86OaV4qHm0s9n1VTsyffJI2ZBPXcKR34M/NzliYDNPGSyhIoeQ7gu5dHNDONyszcaNxRb8
YIBpZThO7les2CkFQNx3601IldV4K+mM8cwt0msmHW3+C5ELqHb5FRetmD7Srj8EflxiIkeO9Wj1
uFNRdrWRyJg83uRHKlfXRVj2lcV70KfyjMesM727ucbkV5oXuib8k/1NL1TLAa50egUS/XkulK5z
nOfpabs6J3HDR4vATzbUcwKYO5DiSpz0QQ2WmMxcYWxtqY58Rx1E9FEcLH9ss/KF69+oHuGGvw4k
YQGn1mc9GS2l/BzoA2q4HHNxX/1Ur3UubFEnIQ9F0j9CvJurDEQYDlPihvzc0sk1aTrPjpVnUqWb
92dgpfPm5kjv//mCercWYFhY4p8X8vfTDFUkiZomlXl5kGQ2su5K2V/Bz1GPoKpi6fqUceh9IKHW
b7+yRadJt2re6eqlxEdj0CutVHzeTu6ijNDC/tNxWEw0/qcBiXtRuYum5deJ1GqbWaqm0fJBqMRz
GyQStml2rBUZsi1A1vaCrltO/XLKDzKmFWs/I25YM7CUV9QVGUfohc23HL5rtm4Y6UQ8jJDpcMHR
6tHksCF1zLMiIFZc8dlb0m4n2mBuzyKXs6/kdkiWU/etFV8eWy54m8LzMEBxp0r/5TF5YqnzoTVU
y7z738otb5jTDnvH2RRT1DPCRCzbh6Ib71vyGL+PkIhKbysduIulRjCQhOYQrfo8suI3xMEt0l4T
cyB26Jr0M3sg5xWHzE/pjs1gpdmdFSHdrPw2gGYdtaJL+SvVvHIhZttdHWynK2DGvr2Nni50OJhn
HTtTJ349YTOcaj7Zi5/mGpO2/iyCacUGSoKdacRzNBJH64nSX3h9RYPvt+o5I7jTIiAF8X97CVvZ
45lbCBANDtMrRe6z5mXOD2rfk6yMoPTfZadmXlHruNLub95vbpIuHAAcwF6Dc1YvTIqXs6kN19Dn
zwQO7AyaJGrSp6sPtZn6KY0Fjy8/N9eGsxZ22iKG15naLV5O2HTiS5pAuCdXU1srZ+AS09KhpC+6
kXn3TxUy3o2aee4nBcGpsVRtdMH4DD1Ffi9Ode491ummGkw1DjwgcYQpl7oOLhLx0yDbw4UpGXaR
7x0amUMrYhX8fa4p1ckEj/Svlay52k3O5hIDfXauSKqZuqDWQ7rxtdKqD8mUbU1VVS2ZZNSqGcXo
AYK/SQrORifpjt8Y7+HnVP0IvhGfuYOZ8+3MPCdGWZWwjo6G1VfJPalydlh1w+pMch2bBv1qputi
xfdKleupTiopQE5eGQobW4SPzL4tDF8rmgk8idGuIglIMLgfiU8CIAhBjYEIQ5eON5PrDUUyParp
ak2um6NMP6c+XlDOuIYRx7vSZDMHUwPIJLE1SypUHz0/s7QSDvDomJv03b69zUiJfbZlsdKAm1KM
UT4EICS5x7lgltXuthiNHT55OYL/soUhMZxLhlqq7pzReNcWbb6O6aglzUHxQ760nuVeNcJs1ymP
FHhfzRtLEK1eW+oynMC2GVcp+S23uiGJRnfX4W+oB/TfKSkBmGKYg/H5c7V0qDwpmP0y3Fy3sz85
QQZJQrhtSKSre60HeyEOu6EcoSCXv2+jyz02M+fdQPcVcljZXbV2iWCC1PMGMKdTHbiHu30sjWIr
JVVPA7zjlLX/+8z/P76v0NQPL6Y3WaMzaqNwNLUbrJYt8QDzf9oChY1HFAQC/zfLrW8VPm+cbTJP
6Lmb5Lzd93taBSRuhf35LY2600opOo+aRzI4Qq+M/IM2+dnP2BkrowFXwpyfjqqBC9cCAscw2Vi2
1kQY+vL5R9jI3QSpmzNBunfTeown8V5AlLMo8+X/U2X5K/j84HXuHE3yRl5YuYjHp3l6AzSlT425
A28fUQkiAqjvLox6b05O8t5E8uwZHZ7hYoDiBcPeJkwLczCYIyalRE2kYsZos7hWbj3C7xT8dKZ6
wdhxxpRFFodW3vBlsb7yGipa3rHpoyE2P4B2JEipgWu8yuLFZKw7srhzYNlJ8MVF+JX9bHyEnTRy
9o+pTHp4krOWer0sBsmpuKaaT8IdGMMYdHGdoTFTberab+JkcJ3q9jlGGanVL0rTk5pRDSwYyRiB
1zip3EOlqg8AjVAI+2Or/j7jt5/ODOF++x9qrTZWTCyZTsbbXnFrW1KWOK3dLTZxIJmqCY2cmNaV
hiH+MpTX/qMZDVLn3pHMMWxXQuEIkXtjRVyyX2welC23h5arofpIdJkkmOkT/FAvNRNkHPJKR55W
k5QqzoSg3ACZI0uMcLNMsiz7n59/lsfUpKqK9X4Tlno9he2hSsdEc85rISi8IB7NsZZTG18mg/oH
OM7ySqA3D/59XwLnVaEOvW/eOyBO9YPD+62k3aOSbO47AU967pvgkUqkD8Mx2w/Y4PJTt7gLIyfn
r5qUXDco0DSmqJSVKWLVUDX3e76VIaF4avstNA04X4RF3OdznikS0PQeodOM+UqZfvBrzZjRJITO
O5qEaLr0ZAbO7t5o+XZqzy6NfyF3FSpF41xkMHF5swHfkCdjgxFzqgYIKIr0CR33HYhPcvAAtKkn
oRnsnHIMHFfMBFdDKacYC7HHfiavxDEqO5W2Ft1CjNOTtiqDJpM5Wma5+lxeErs37nirOcJvtsu0
bln2uevOJ1YoYTxuQzN6WjsQVXbp5yIJuwEKQjdhUpmRsI9kyhAddE2ENo4M5ZBVYw/7DpeKmENB
NF3Te9yf6Sr+IrseqBuvnlTQZ1sO4xkbJT82ZPGIrVUgN3EnEZ3PdmD+BjY7GUiy6T3I0FTj7Qo7
WAqpTfqOm9fG4GGWgkIoO2l1xLgQTs7wBdLN2jq/cvtOBiKObdDC8gC7UoFWPCG2dRb3ks7RW64R
PY1gZ4tuCaRk3DdATeTFcjCYvl68n7Im7wzxmhJR6aXzS8ycLq1oTnxHxeKkuT0BU1yLRxByNm5Z
EHwrTzaXjLqMdxAujw5sUPVOpjcj/MuCwfodjzcsWVBAmjFvnrnjKAS52/MFC/E2fUQLuxcOrQJQ
6WmOa45Uwu9gcYQSApMvQ5OVoJk1dqDyg4fKigtf1Ua+eO9WTkFQPp4UeCSbtRYaudNvppzPjHmt
uDsAjR+8XMub+Wvk82ZSHQJ2OGWMoHJyhO3QHJDcJqVXP8aw1whcoVho1BLROII64qM0WDrVK/GM
wjMkKvsu3LKsoZ8pY1xUll9awhRZHn7fFNdER9B/3hO+SPtJ/cXt+ujJgpveM6WC8rGCYvpCmoAn
vAHsuwhWM7VyVQBoFciuTu8MQvulP0jZJuP8D/QrTUX8QMfxYX9EZYCXp4vAe09y+v90Tcqyw1Ql
iCuLQjzbyXAO9OdE6GgOckyHWQCH6WBkAzynOFfI5VK+RY71rEwMB9VJ3D6IZZ1xfGV4eNwaPlz2
IFw06u/wm7gwjNsUAyd4EmUYfCW/xFcQDXhf3Js2a1aZnD3fXXiVrKo6be+MGgYzNLZmb83N8iQc
QtuN/70jjhnQ+3IS8BK/MJYOsXMabWTvHvqpHAnKHRFzimNIqCqez9jUD0ARoeXbPXxTxtKhrnkh
QDm7fGgieonIJt2TbB7wxJiSh21Zz1SEdULjRHgpg8BjTmzWbzumqHgt/Nl8IoAOr/qvCu0PHrQr
qnrnIU7vPoptIQU1jCl/uwaAaQluApqaIiapxeFFMl0WNXUQj8z/fc5/0lwZ1CK7g3zHeRPCpvyE
929BAXIIE5s0E1tdPLQ/wkKRJfzJLBwZ6lka3C7/zIUZLhirTNFr9JfoNOUb+LeYxS177ELT7KKV
GalS+iHxpdt7847f8xZ97GG6NLrIfGTM4O5EuhjFPkDEIxJAjqy0e3uaCBIq8CAd++F1JDLTEJNB
iPQfWhA1U1pjReB0/t57OxnR4mIuMvctWwXYdu15ccXlBCIbCK9n1rTnJgbwdQOtH/yt9aSYyRE1
NWLS9fNxAp4qg9Bd9laWIcigrOCf4FxrnLhtVwzp4bmrxfZRvRzXHvhhVBgy85SkbLStIKp+zg9r
AROS462wi43aEls+sCfqrK9sm5sSTC4UiImEKzPdLw7gJeQEEa4FgiT0M5a4fERL6FE4OA/Hwsc2
ipXMCKernyRE+JKwByXBk5bslOgV2SHhwd68OemFAhC+lVod8re1Cj/WeoI5i6GqrIOrveL8BdDX
SBRF+ohReHxyb0D4ci3H8GkNPCArvPN4IlKEJvX7wwSXW7yR9TngtYasj/v5YgKApS7tx5skCwVE
cq18jZN22T79vzXkmVN/41glOA6ejoCxpSbYOigR5O9BvAnNrm7c8cpzIpLKzD35vyie1ZVVRjLY
E425HwotF+yez8XeOuVmm2EYh6zJrq9nc8u+u0jrWYpKJ+sqYFJkaFIQX5CKiPbsS2C10/QKbb9E
m8Qi2DZBlthanlHcRMuIuFI8FjDQGtaOjVnZQ/wqAPSuRlT41d8MzTlK2SQOKJ6jXWqIwMkR/DqZ
kvdY31tXlWOYQa0I9KiW0fzSF0wKokU+Js8PIsTd9sRY855D5Lpfx6ijy8FFb5HSjv8GPPi9AcjC
YxApRP0g7vgPSKnoaOoQVwevCSJs7kY9Giw5r5lNlLfskwq/2U6hc3TZlHh0VQYfh8p4D10rs9Eb
kVB6VXOeT3dN5vwxSAh3OosDA/QwWEzF1GDMr6LdbVIyJXS1I5gcqssACf2500T2g4lwWhHfCZSC
aEUwISKZZW/S44yJVRqGwotE1AJt1hDnLmBKD+fchDoOicu0YecDIqnQcP/QTgilgoA2sqOXY7Df
TL/2Nbr0M1Dh5VQzzF6Sw8KGD5MTHJgrNJQi/eCkKxoAolTdamO8ot7oT2+XAygEbkbSj7Mmol04
Q7mO3nPi5H+/bJP4uavH+bkIEwbgNKda5Ho3LjA+KOVUtKgnMuao7iJeq8s7LsU85yW7XgujfUZc
G+EvSUVW/VnGsVTTtnpZ/uB+erpFNkfaoBcwr5X3wgL4J8GKhuNR5a28yB96QWW7GDl/lbqlrxRU
Jtj/LqSj1et1Arlzzt9/TMvTFzX92r38tuF+7uwA5vgi1Peoc8suOIch14Q6WuWrGn008P4+DvQh
D0glI2E3iVLqT3EHBd2q+UUbGW7g2FsqoOHokjyKXvB7NwY4dfb/P5uCvVHEzqEa4/BwVeoJ6szM
yxkJteaEjyDywW62/rEbdnYu9g/pUKuiU+LtgO8wT3CE9g1jOT7QfSatbbfFbMGJF9osHSjKklfL
kc2S0M4GqAzzRmS+13/AYFJs0EeUdw3sHs+JZOgsN1LFuuCf+ByUeiDDcdHo/yrFuTDOsygMui3Y
JbmBaTIg57Y0lW0QclH32msd1JgJZwzX9FCwgiyx0rz7Zc6J5cy7VVsRrtUeQtRYxmK0Aj/TGg+k
Tswt13R3L2bIXkZpzEB2EAmiH3aXReSC/C2GPKLXlKAe1KexjNHLB8vKSP4Pzb9+ZIHG+yxfvf9K
wexQ1uxKzxOyNLv9Ob93JMsBL6eyhPebFem6PCX5fFWQ1DKnrSFOQrDfwckKAoHRNNltGen/6OqN
FqpCiei1A7TdWOmHBYLqb037TqS5aDTiMu5c+BgF2qEOmZBAfoMlvto9Fv05UFmJ/pDjwpXii5Kb
KbQfC7IDTWB0ob6Yy+aeFt2rMom3u8s0yYJo3k4aqC9z3ZaoJxSH+kvfSYJbdUbNyH/m5xpclRaG
Ac4sTxV2prhFtv/TVPuDNfLn5NA6yoKPzUc2+CD0DLGYX3DxUoHj3tMdt85h50frobMwaW/44wp1
ZuK7VbSw8DeCnjQCNTOxbfvE81DOmniCPD0MRUfegKW6h+mS9ZmQM1RAda5WIcHilkMkpfcVZTDf
B/UqEI5FMCI/vaNYngpP+01d8SmIGXN7Ljgli2dcgGmkUax7mmJl9J25F5ZXZMVy/sE6MhFqsLo+
Yvo345wtuDBfJ+2tVv0pAoNT7jz8EqIiXX3cyG3H6H5KUONRnaK8dVx8alh0/xX+9hRnTjMYRY5X
hSVsYinGP+nvB5MNq7cZVmiePCtoWir+bTv6BBYzTjRYTDsnwJfUSDu4eLXaShwK0YzzOUERh9ss
RmpGz32NhPLEuJlHiR9i4L5p7LeZR9IhWejE73vji1B5XOMq+wHJ2B0aLU4T8BZV1s5KeS/8H2dM
83hGOR8gJTAgqJKmjBw+Zii7CXdhPSl2wR5mW5NXAgDDX0hFRXqHwW4rKMRqP+LcIQf6D9niyjbV
Sma4K+EVbKq0QEB+E2ISI7F3vsJYkMxEks/dnCuhe26SAbjxzsyh+MHswCIvDhUjfhMTtjsldrp1
QcZqAy8PcvzVRckCvVkBA2wRLg6uViPnF45/s/gaJrfFfRIGl9S9Kvr1ItMfRgrnasOAzwD4NNts
K4ZeVf18hVQ8Pj9UygSVPF6MrKqJmcEolzYNhHtWZli12KYT8Z60ktzabwnGym9o1JGy6Hjbwn0I
6Zm026rkIL4iGC537RonNxfNukN1C3zDl/MUxBnY6ZmBWZGKsGLn32rzjycksmTQV5A+L6+5qfpF
KWberlruAw0OvImeCpgoycPzmrcAgranYJKdoGOGzvS4Jt9NLjWlPe/dOv8TeNvo9ZyrhOKNq8Z8
7h7gThzFL7XSgsYnifyWajpNUQCSYTI2FtwqA4qF5UnySsSx7TTPw6eefxzs1DTA2wA9AHP06BlI
YZLFgg1kZ5HeekypIw43AHGe03i+DF1vtycOhUzxJgp7rjfn3L2dCKRYv4Uv4Hl6rSJX79+eOb/M
YRMe9PiXnyRN3hHW240hPfAQ1xlw/M4Rh9H6Jy3mzUt8kfyIk4FYNYj57UZpX9/svuMc+8uQVkAw
u3gx7ofAat0tpotHonmNx9KhKizRBlWiI7afIydbJkIabJi7WqN9gimtgoM2wXiZaFXWYT2V0Xdh
W1qURQ3L++0ODVNdmr4Mf3GlASs90lD27neEc2ILKZ0QHgT/qg8mcD08lsOpj/XQdrupAxocDOiz
bNEHlZhuipb89X/o5DP8aw1q+5SRZ47fBi3D5gypOblV/JS/z7oShdcKZnR9Cuak/tqjIBpBMstT
YEd1wO3ELYZW3alwHVp8LXNJpPNZ0mvMGK9a22c+w06oL5eo9GdGIX2sGlEo+/3h5VnBiJRqFSbm
E4411H4YUiEOKGRyDlOI5rQob8l3c7XB9RMlmN9gcA3ECbGsCeUFTht8DqLT3PTHVnsJ7/X0o/FX
Jo5KNW24FdI3Tvu2k8pGaKuuQByXxUU5RcR/etWr6h0Cfn4I6bmr0+jpfLqa9wBMkhD6Or2/dAqi
sHiqbgB3biRDySxjx3SbjBoKJo8Dc2M9PavASHIF4s384Vc2EYLnZa4T+/n0caJHfgrTG2sUVfl2
k/JOpltbwL3s35hq/fmASoT5w0PQq3l08D8OAD1pcIrNWu7MEoE7Vyyfzq2wBNlpS4J7BA39OJek
VzdsjecEUqEBD2eaiFvcAVS+TtI+5y2WYeQj/UbXzPNVmAZImMi3ObhJ/qVAnK0RpCkEsWXIr01g
5AnRceStrX7KhadAPT5raremNJ9eTlLRRXdgwaPo7BQ7Wkk6VNayH/bBs480ZXfvqqoTBr6j/m7P
+/rfLTHOJQqwCRgQtkPBx2tdC+P01DXnALM0CET14O1bh4afa1rn/4Lx8xp+UT1aBPo8VkeDZb9K
FZyY7rZ6scnFEwcWJ62CcxMkOsyrDl1v+8xA3BpduQyHoOn/F7WUIfc9NJYPKWsyoAljMVqR49m5
qx/frSqWMN0KKecx/1BgG8ft8aR4CoT7+RxM8aNwa4oTm6oi53TQcEbnJQn67UUnX4e90rC90pfJ
IFQ6ocQF+A0IqLgSBtS2i7vTSUkzE2TeSu5p+iwvLHnm/FqIEdemZgUb/XrEeB+AbJWMl3A/NJep
MTAZr4xi5KgWjduwK0VbxhZtg+dQFEiOtrrwhGf/GVmGxoEEK0YFBmDnM37R1Gce5r0Xu9zK6Puu
ah60ILhTtnnMhYO1/POWsp4WdPdHbZiHjcCCnoacrLqEMXFyhnw3BO/D9vRte8D4/VQQ59YKY2ZL
hdHoua7siANLPXMtHxh59C3zVP5baneB25Sn68zEKf0PbaqFJr4bvPoznpLSkzoixLxKdfjCaEBN
Ud+cxSeNSDhfuKNcirujeqD4qL7MbxvanwmFsM4czRDe/CU046zls9UXMoaLR5ftm3X5f9zRD3Q4
bwitV5ZgTHWyY7EnkcSOpDBlE98XsBnjl9aSfXHkS8NDdDDcm4AkZfQH1FTFhYQfhyDC9w8zLGdr
wCE7BMBU6oEQecyEK3Om+V1sasuq10pIZl9QBd1/z1dXS5cZm/f4XzJ9vRXUocrFwt2wcOn3VTyB
/c7gTdAZ0xZPk98LxdGz2pg5xqcZb+uPN9bMHMoNe6Q5+Y7245bdFvDlJ+MzmkRperZKfYhduqRf
Qb8dr3xg7vWSiEBq0Vm+UriHzv68O205rzG5rELXcvVEr+xqpyQSgflX2g5hbaH07qVdBuZdxSwL
76BjVrjPA3H3fZnRRIaGk7uCIWg8yishfsSOTUQ6OwsxlYsIEz5cX8poq2HsddmrvV3siYzYs73v
sllnBhzgbd0y7ngL0yDLcxc2yARMAIypWQyYvI+drpUKHkLrqropsXuZq8H/H0mnREbLVNENCe6x
vjuwYf7uklBUI5bBjVbQAvezGE1go8EKai15+LrxyGI6EvRHgPN7VU8MqxDRteUgBzQD/Ujk5fIz
m04h5rTEUfzjFQEHimUAcSqHrBguAH7frylxhH+0YNQvVJJEwynWCh+w7sQwCsW6nveCvBOHGvef
CVRQrmsGGHbIFvc6GPqoQ9b/4Fo564CUrD8/rYztDC/7AH0dnkriyYv1zEfO8FCNJZw5PsBrTjd+
n8k51Hr2xD0MtsosgiOwA+XED32wwe1uktTg5eoPfnpfPqMOeLBXsGvGjqMy0KMpdlctOJLe/pkr
ZpvBzqx1bA2CPcqRgdeBDKwvuQLuFZFVStdx4mbMbEui5kJoEP1Txy0GahsE0hHQKei1PvvETtqO
pQKot2PRhTdsg+987tkVPf+1Kdk75y5ygwrcJuMGqlY4OShIBxvMHMuVWSVGgM9KuO7mcLunUOrQ
YmlEisHtNf6l3WXb+Kp0AoGo+XcFbyCiFxgKa0Zgms433yfY/qjPVFEi9r/PXJRYeln3DcnzGntQ
RHJD5WOEJlIEn6uykhCn+W8X3W4HQpO2NtPV2R8yH3fnjyazu/UCi6uoGuYEFNaWIFtjK9QQ1G/y
JuH+M2SAQTIO1Ojct/F6Fz3oXEiLkPgI5ISsnej2WAKkfYe8QppErJPTMAFqOFulStHeqCvEbA/5
K0qCk8rRt4QH60qvAP4yX6eo9lgogA07SJWeNWvrhrliWW2dXDw+BaDyEB7zLUjnLvLsH3XRYvgA
DwP3hV3I9Cxw8PSA6BaBtl+w5H0aGM4wKCGZast7vBhh4rqmLnz0Q4dUNIWgsiLZ6ISLHzfyFvZ9
9QqxfB/st/Av8xv0nfV82nHPgesQmuRAXwWAG/YWPNGrWb7+e38dmIam9FWQvhdF1CxRUj+UMfbI
AePJz60gT3s/tXz+BbOcgF8P6a4RVQcNACs8CuBdS2nHlltr/SyMHzUcHQh9CY5fKUpT7QmL5K+3
63mXVXhHSwFRZU+7IB7em+M40BMOOluXjl7trkCkP2gc6t8XQuuyabP4YjEIOdWa4SxWnGWfC8eO
JwAyL3eKNUolbXt0E+XeMbqFzRXdHNbFxz5PFQscGFec+UkLoKOmXiTvHoD1bTP5Gt3QOCD61n9T
yXFE9t+/ZXOTApxq/1LFoaizIGU3BAD4OW9msDr3znDRrU/LXKtXMcYyrJM+oCj8spTgal9f4mIh
3wHKRBOJD7+DtcvwfItn3bjgw21bhe9hRnB9RguTigEA/qP9b6NkDEn4WuRn1ImKLdnFTFAt4z0t
veDgsp0KnFnfh4+CjmJ+aj/NU+EZQXaXdrbcBjcvBoT3CnQxCt+LZyeFQQURfY9BmBRGL87Yyrln
hzLYst0qqy2pG0Wf0vOZVc3qGtP91NOfIv5urin/TOgjfGyO6SAZFkvQFw7gR1WTThGujeqS8ZkJ
ngqK5UgcbU8UvLwCLDtOyUeXGEyfYAIn2Z7SpP5RGFb2Gdj1IQrhBKFq5T/0TulD6UCsH7k/fJqZ
1/yzr/xea8Bg7319G5zOBYSLmcayBOXWv41/I2kMlFT2ZjIJnRdu+5dDsV4dytOxcC4ffMGuj4Y2
6Nm6fHb5u0fVt04AHXkB+9/V28HtTbQxQVilTz9JUWYEQ4u8UL6AhBRn7TRImE9PLZWvPb13oBOm
UUdvrQAG4hGuT1PxbwtB5u4kzazwipLrT6FUc4B6AWM7W62gtb1NuYGYqK8RpryZA0Mn4ogkE0Q0
dUxemdsTtUcvyQgmhjftoO90PT9hR7+Q/TzMn9yC3z9xSOdi8p5TCsJF59SIufghSXIJCxDZA0gj
xah9ZwyiZfbobYtUQ3WIUTk95KA93+tjTQzLNBrxzdyb6k82mAEyHRCEs3Wi/JD3QMxrebyQY6nc
bWHkAGXhLodyUX/wPGN3wRBYg7R1chnBdQVk4iWfQjn1CH8+aCbnjtzYe2dozTjvTH8s2OS7ZcaV
uUYBQXAj17jnyKHjcbxxpG1fL6Z48hXGCeDrfgaNulZHT4qqW+RHPv7PcaL+WCTu0jYevX4jkKQn
VjbklYZtfxQBj4CsDE/xWazMZ4QqTCxy2LuJ9dm6dL+OXWbiPGpPE3UoRg7c2myMRN8b40HG7u1k
VK2QHlyJINlej7YcjuNt+SDusXTm6ujoiLSy/u5B+I4nn/0CgglCk4CUDqjk2DDViFZaXy5IYPg6
/s5Nmv7MzSfhsk9m7ftZhNwA4eqzjZBIgFnONhekYVwvFerGDLtK1j7x6zH4OBMR/GzocYLuIgLq
IGLKiBa6gNyQEHK2M+SsUtCryb6bhr4I9blxkCs806N5mcGRjYam2vXodBAUD/ZD5nOMuzjeDDes
d3/Oy0OFtuKuIjEOBjwSgQcm6c9Qgh4XAiCxmjI4v2qhpZ0ts6tWNhwGnsPWIE0olGWSdeYHyfCN
f2IVeSEH+YnWpGsJvp1LLozREfut946psfdllEC9chvdAEyFbFY67IEIGdY5royuODhQW3NYGEYN
hwS7jzA1/gAOyWtei5tRYMAO5UOJdHqNCojHfUINj55EdxywaiSTGeEkxd3mqhTfUhNPdVHapU85
rjiiAoHNWROtdw2j101Li8MiAqQRGpiws+mypb0rx8AJA4ISSwyKGXaQRh7mUneUMeagyRvgLjWh
YvoKHnwI1EltvO8x4eMSoUE2MRTH3bFYnkUIjtD0KydU51qGwjyeHa4/Owvt4r6AagOBKfwh0oRi
YpHWmQ0LJaOLCNapq5Qc3xrEtaa0nwZORTtkgemMSXWJOiS810NT36G+eXzL7bbv5CHNFWIpAhW4
qUkhbT/0LtniOVR2OMAonsVFTPDO/7U2v7TKv4WeL5/wKN51Mf7IQDW3ed1+K0I0n8fzBNROhMbL
C4ArTgdq/ZzJkuxs+9RX+eqI5HWi18CMflJtCCI8HaqeLj7MS9+5TVkI/F8C3eN2WQ3vI6zOMA9u
v269rqKd/zv5bwiJvMZIaumOK+NSskuyGjbFIHAplqorEd9amqJRrjQd3CGW8WlbYVJKijtn8HfR
kEd2AqaMn5De2aIUnKKrNuv4UUqA0bhaGEvk4Jy7gS1O6wsWaBd6GrlFCSG9FwAEQmQxbeOTcbCC
xDRa2YtlsfyNGbOiMPBBh0IKofKDSjG0jK/kUrJr4KzY9ugsLnZV6jYPEkAPSd6VXOK4o2o4J3dp
z3nVN8vSgS0PSnIWEYflphYV3WtMyc5IWUo/WDlZ4QQlw6RgirFgaZ2bqpLSC3BTBGM2i/srdIAm
4IfKQPLjRw6ZQ21hYa9m1h3qiog2gwZQYcZdkgnmJmXNjXeBNB6Ia74Svfd5MPttAzLP4Vawx4lT
fv8fqd1tJNnnpw08xRda9rYA8AqVKkkzxSbr8TIYevmn1AwEMrCKhpdF5RqLXFGXV3dgcJtsVxfh
olGaQrLdnCwC6BYwjBFWGtqEVy7MzktCeFq4AT0qoxZhaaGODRsUe7jeMh5xymphzAp1dY/iZeVW
dxt6yqzYsL7GSvelIQUyTSVez3F8hu6ghbBdZcZ7qDaBHZPekepKt1kYnl+ERjNsUQNZfg9/+bDT
snxYWX2gk+iEVUKaLzb2zgX6Xc9B4IH5JEC2t5nitCBuyV1ovJzkAKoC+eEu4uSMe3trRnomvSUB
84cFMnRCYAJbRwtFq4f8vAgGAXKtsD9VPQTGdk9PjS0LpQZ96ZnbSILnYjpXqnQAd14YV7JDtmdT
o9BbaAGRMhdTKwc5YVUgf7LesXxe8jT6spAsNuNJIC1RyIiqf8PcSfQJzIwB67QXdW2P63n6Hfh7
Ba7ptntM5Tw8Pgog0P5sdAr1RsfgdYEo8ZcYRgQLJM55EMFKjz7f40I1Vq9U9TkwI+8VObH+88Jz
ObSocj/VIvi/2+PbdBjPvTAtvA4SjHp3/zaMfSuhEBNlGM7UndWMuHgV6jMYXQr5yeq2fO58dy7G
0khXxi/kKhFVpQ6XjuRja5bJhfjgyLY+U7H9Bhra9uYoh1pvoHjg2YvRfJRenv9ROTCekshjHCgB
3RGd8bI/Eqr0VI7EBrZtBq9U3mYSW85fUw6dXlQkx9RhwvlZNhacl7GkqffM1cwlX4nLmkP4TGg6
ybcLGRU/iWC+OC8R1Nj5fwzWjJEBWqQjY6zXu0BbU+yj21+pfphrWODuM5aE4j3eaZBSzMyMyexP
wNFSqL2kfpycD+s76N8Q3h9NrXloojGUwVlRafOE+44SXZLgT1j2O7NoYhAH3UbSC8i6jAB6NgRi
UGV2LEeEyNi6MOdDOHt1bedZrjzcVuEhMv7O2O0xQOgO8M2Fc5l/DGq5Ykt/NiooL+hnLUn3NHIL
z3qel3hzZcgvcE3wREEuqfFDmP9LaqvMArsDZmPgn6gZVLS6IbU6DkjCR1fTNi8152KPy8LljLXm
1FphbmvQeWfkZyKSLIK6qbg5ZPtQDy8ARXfXuROFcIcQ+V63eDYD3zWAD+aKyxCZk7puPnSFbpoe
aGCS9jsz7S+njyH39uw4BkYSlFocYiXZ/Mnb1GOwQzVTNRDQFbc7hiRbVoAtYF2kSodsyzavBYoC
AKPVYov2UC/CXNWlXELzRw7CEgfwby4u1VjhaI4AgQ5S6AyoUIE+NNcYRDFr8XTffynOgKAZIOYl
FHllF49PRH4YFZvmfXdb2X77Gd7B6Dh1TB68+g8a3ciA4hhGF6aYgmJR/y/Ax0ScLClE8B+pTqpz
OPbdPV6DPP2kWv4BUNsv+Fm/r0b61gz0iGIKRb0jVvnUrwq1MWHN8xkleLYGncoeNzDcZcc1xWe3
T7tTPzZl2KPhig/g9Ud1nsrKtcMFYTia5m+I9s8BcsRYV1ieFe9VUJ1QueOWusRcFQbq51qLnE8r
QEOvR2RkkBk0PL7iEJqepO24dWpnPTT3s+35HSUBFxYgAd66/p5k3cj2X2UQlz58k8+OZH6PQoQO
6GrQd4WiU4dtE01QyxbgBbNhJ2AC5PobkvIYhH4SoLXdrVe0v8PQnxbt/YahA8+NKYqTNfyhjKbz
GgLJXdjB+trHS42xy+kBlMZWbGSpR51Ebv/2T9NxyOy322Vb8Joh62hgs9ORcQmj/MKIZy0T5wrY
W2AH4dnrjb2LUKPaF2NbyplU7r+Fx9kGZbO6aHcLPVkPMjhQX4KpVaLtjxHP7UTS8ZgmofEEWjNV
U/jV5+TP8cyLV0e/hQW3Dd2qyAseIfVZ2KRArzdbfjsowNbvH7SVEP2kgc9fAbCvidUuZYTjkVOZ
TmR3H3pwnNQqpW6WjF3EkhNx7dsxj+dU7aPctL4CKvtfE0fGud4dYkxVcSDoTOiVkpPozTfdTdDi
XLc4KXc41rW855+E2uwQ6YYCkEdp0QwK2D/I6q2zGEGa99WlSD4AIfMtE9MT6w8ddy5L1uiHI3b+
iXKNP0Q3d9soRdr8Zc5CMb8KbqPuZ5fD0YrTURw3sQ23bQM9V3JjZOxjE1H8Q/3Jd0JykWfc8umP
MPQ1X/ouQcgEXXvMjqzdnfo59y3uiSTovf+OaCb5ey+inL7FFXjg6o4MJcJEHUY3599YJ2wWpJP6
0IIPP9XwT1AnqnNQauhINb8qAAlyKgJs/NzQJO4fpLXMMHypuiBY5tB16A+Bwv9kzKSsWEGB9Z+U
BAtCLIsMykVgXkJXYe3V4z8WVuqSr6FiuNjsuAvK4f2mJDh0ZQQ201vjaAoeqmW3sm1d+UwknDV7
8yOn5Mnmigc1V+tUbZ0uoT0CpScTaaVxTHP6lQtDh6lM+vTbsmS5VBz563PKvcXdsLZGz9PRh8kA
w1Q7Nd5mD4hsLwPk+zXhWK3YKHd4U+0tFnMlJ1LSHop0IfhWxtv1FixuhTByYqHp9SxBqmMvxTf0
xwEJlfnYKg2dvmFa+LZJf/ifWYx+P5e4oM8/HYkyNJSz5LUCd5b+WXhEv9dzEDXlNkokZ3UGmBwa
+vtxdWTZVKltrk0gyrnZipc4PiWFjed8+iJpFLPanKfXZrXq/OU/4N3vARiMsZ5ugc3xIrUAI/3U
3yu3sYXv4y2clyMAoel4rRvuHZgkizP3w7L8lo7g2FtBhXX2ocTdg+cLO/JSNxVQ6tDo4uYxJGGz
7O/YAwnIUuHFj8xb8RHf+9G2T2UpzKpcBCGY2SaAmyG5Px8s2VfLFryNwxK2+wLIp4+4dPD+1a3r
Nn1aznXNqbVOOiQEwcczwpP7OPtxk1vVJOabZNmWQXCRF3zwJVEY4BB5jLgXFDj4BDwX31dB5Vde
OLm1yebH0MpJY/rWSjHbrHu9tv54IAzi3KhnbBcXhK6iE+T+7yYF/RBanJjn0PJa3cvf7ccUmrY6
5PSSONqnRuOx9I2O8wW2i1ZW+SjNPUvK4QJD2EGVEykk+lYL6UI21Jgft1CIMJ7gJLFmne8lZ1pd
LHXX6pLvcrjaS+1b3j/+8IkgeigDkOYB8Sm3WTgtXtj7CGWT6Q8jLLOSjQroJsl9naz9reNh7UCc
PYGG/LvVCv9rWfSaRfeqOyWfhBjGKAvGBZecv8PfkISdO3bgzidY9QCSR+baykTeiUX8WBHJMMR0
sVXJg250Ptz4A2zU9DtbUToJ3eZ3PgdPXU3lepj/hn9rrbfP0O6Sx5uFUB8AFs/q/xvNGNqUeL3q
rx3MLVaklw04iyqqUAX1DV6THT7YieQqY4YavJW3FT15fHePPWW0CROg5MQ0nUKtF1msPaUbX+Xw
nFTBUB6paMgYY5+B/F/3zIJS5rDEaODifBfZA2OVXap/xLv4ooL0NO2h8w/BPob56pBhPPyFZeYG
sEjdb3ObVHDs9b4iUPtgumly33yjfIp4gNMpZtm5JT1lz27WltPMvxERnE6TfvoOozDHzHrmx5P2
VY906W4z6PdnKjAnzDgEQKLKr3iAKaWmrIYVQ/AlrJJM8rSY63+qcaPNrJjV4MW/MlS/E3swru7w
sveK6sInEol1IsLosUS/LSRmCHm9fUd9nTiQxpH61F3ks2NVvn70YbvsN/g1AVtNWlR/XoUSTx8z
dYzdnI06xpB0MjTXMGUPRSgHSRdQ8a8WUNEOoSsJwLYrHj+fbdqp3Oq9NBEIwPqI4EwUp98wYTUy
uXcUFmrZpB9sI0LLoyH6J2xaVFKSF+RPG+c7aLaZXVc1sZuJhCtKZ17JPLI2zBhEYE7xIWfo24Qc
bSVyx76wbcIbSlEe1uIHSwJDj+4eapota1Dsk1XoXGMG7AtTpVw9SA0PVnqJY+XHeavZ3Ss4u3VN
ZtTtrKWeGNLMP0IWTgakE9ftJEg6w5X6HSff/x1MW49RYexorikyK6cj9mcn5FEwCjn/UVsQhKzK
q88UiwRsNfcFdN9iHBTWor0lW4lYd1lFnEumFM0ylMTpGU2qFGcNSAAnzswPBvQae9rrD0ODxnUB
IFzHJ0GcXCywNxcES+1SFqK8Q4zBeXtQcRa4iH3qdhtLgE/u85TrNYBSqAP+rPDE3xaU0W9Py+Bq
pd9pW25fumxQ9EVgD/bktyH+6Ly/EpxhYz2kwHjNcyEGeFXYUhneMJJliDJju/ljqKL/Me11sgzx
IFNiXrU4noAPw68HtP9CCAft5M8hyj8dbAYOk+slaK2OiDnNT8NWMjA91m68jovE+eyIkUfC9PKu
P/04vUSRY5g/4Vo998523b7lQn8jaKtc7r894zFeWJJOhSqbndQZqFUe44m5blFczcTan3aCJG8m
2P62oVpMRxYrXGOjkN9UIZrlrbFlN7e0u1H4xXESUSHPgKGGzeqTiE2WsEQ53SZSzLUvCjxXwKO1
+2SatHGCNGVZve0pT02cBA0R2Ai67ed8hZrikJO3m8TZyh93SbIqmhXJLXeUWOs/7buZj90CFpLB
wjfdTmC+O0g+Nq/05zwCKL9cKw/2itnznWNmqrrA2/XCVJo5dIQUKtb95LMVvLXLtoFpMNoDWD1C
Ed8BZ4LsyQDcVO7iMyN75GyXPGVnGhEGT09MQcFncnob751GHwxPE7ZMlLq8gnC/vEXZ+iS1ONqF
EAIkKt1Ry9WgzztLPL6EzQ3dffqlWJd02AT4gtZyoMi/z1afQl/c/ic6ts51ct3FX9wyMbJAeXnz
Ij8v3ET3qfG04Z+ng/JKr7F0mrC8BMzmuibUtHU+ZO597Okj/eXXslJ+uVFpc6DtstzrzoCy7nuo
me0O0SPUvUs0PvYWOp0zperHAKze0AgzGLzNatNprW/0N8RfXe3JqhsAsF/zkT6O+za7sOUbJoUh
Vgg0bLD2470toNkZz/cpbDLz2wvSYEkMXgCLsqwIcCofFAMAb3IEHWK3bPgq+yLHoFOOXbi4Rist
5iW2b8jPgBZHNVSDUebBN5ofdIWA+mGzUohCV09XJWON5W7Qo1w2ha/rIFPxD/Umof15ItbasMml
9B88tdeaAXNIcgOWiAhSqBXGxA4yTzYnwAKEiGPQ7CqdQImTsc+Fd79V628YMZovuqkwLraW4j4G
UhtGHQf1sFReuHS/KTz947GYsZt2zOTjoxigXYdQCqecJexIRrFlaUVeEVDLuYQ0Lwz8HUdL6nqQ
4itm78sofUfQ54ojmREYWPPh97KrsYqsRZBjApzrZw82JtscLOMip0rXxRLGILWJNSs4K2kUZkkH
GBmZdccaJQNiOt538PDU0cs81fwb24UnU8DzkRdexanMTPbjzP5UPEuFspJf87GS8bZrQfdvl97k
66F4ynvdTH5Rvg59a7W76H7mg4W8n5mHupu/ThCo4IfuSQDa8Ownpwn7LeJYYW+5OXYM/yP23tje
0hnUBM5Ys+MnRHRkC/qaj12WxDqT9t2Alt9bz6siQI9f3TPJKTZX1PY11MlHH/irF/lNJ74+iA6S
eVujnkCsWDwBEpOslHDvcED4yKcyX0ksRq99+B7dhWi42ui99WGBeN4//tT7aImmSkvTPs1i3iru
SrRAKPdsqNFSQCVT5SS7jWSBlzsLEQTmewg+Rb0oGiyPO2MbzYZgk4MDqjn8wcJIQcxMEd1nYYIb
zA3tRqcEZEZmB+4A9Ksba1/dloGl4zH4g3FLgn/HgYYkX4/bf0vgod3czdbBMqW6k+nDTaoMRd85
ioeOvOi/tXgON6CCg43bd1EXJCQ9tJ8OL4gMz5+Gs/UXeYfcfB1EQ2cCFvVivfmzgvH7duCVdv9N
A33UXEG5VimkPzwF7f7CbppCzyi6MeG9Kh6M96zY1tQmTB/KWNF+J4ChllP3+djvxgA438AczQs+
+0DbCWqByKZKxszlZm+rPG0BfHQGdYwTWt4/pB/XHMri2My5VGgwqBn2154MfKDDhn0WHXfRD9ER
MIcMSQI0qdnaOaBY3ASRB2Orx/JvdUL9aqmkX8fdmwjAp6/dKVUyAtp0lK18lhuEXxXqGs6p35GG
tGVLkxh381sn74TptaZ40gYVXDTAfYvfNLC/SKAOFXPuVyUDmziU28MLYJgqkvdmXDJJt2EZgh6Y
S+W8TOXmfwwfFJH0sFnBy5pWgNa2VaZMZe+1grGRt68+lWQk0hP+Xcyn8rp97+Az0vHRhlIF7n0+
kaKGPfn7SwaRlnKttPl4RtrQQB4Rwwz0jqW8iQMn/S55U6oMoYDROmiHPVOrrMTC1uctnoVbkXRS
rUy37WcMl4FZ7r9TLH+rAXv3aAGKbhVM0/HY7JrRoUBvpJc1hUnm8Zd3auHC9RTqS0tJyg5/vGwz
a6NajV+GjH6TS3angd7lWyPzGnhHZ1V4dYdICfjHzu+BnljYmCns9qV028f68C4UaNiivOij1ctq
ezpvg7VMw7khtg16aNeFfJ2tH/Asa0TPNHDRpCsPGJFR000MC4vm99AfVr+Jw5EItWvErETDwd7d
kZFN4/eQeRhbB47kPaAm5+FH8/w4vArfNYa1TM2XlzV6Q5VJNLFxmwRYzfccdUiUBPnd7UIBK4D6
mAGuCzWZXVaQxylmegM/ksqXdyux3LsBEgmBps4ltxTpWOsXPL9jLK0oaJElMRIKAx8HXKGRrtIn
AbhUUMrGP4bOS46Hq732fiNyqPngCM2tWxFZuZKrWhumKzXZm/uvzc67IdEAXISkq7UIajagwjKU
09ANNsIPpH36xS1qPYxIestlp84WTOrfXJ+QMnHmgz+2UlORUQPM34D8/7l6Vi5Y/zRLi4mHE2mw
17DKYB6k6juEMEy5pCMczAp/Uy6NHnG4NYePmbNMaDRIsOO/ZJRHYiZ5uyO5qVKWtE9y1ydGGXyF
+B8JYcu8acwgm2ZLHfog7Z5X8yhocZb1JCgj6uTeflPHmdCXvJk2tTkip8aQuVv/RTTfH3QZRosu
6jLlp9poNv/TgUGkQjN7WBQzscYS+Tj9sX2RA2KxQregbXyp78UgtvScF0Y+xZ3QV0VH/j46HBpY
yknO6nQPATu41DvC67/z2lSy+VVGZAMzGpBNpCcbvqdG2Nijvd/F31mUXmla9Dpk4s9PYFZHrd7h
fTF9TJEzE1MIQAEJff5wlreIbDOrhmkEuvOO+s2jr/WG1t6dQJFEBFntxrcpr7E47mD7tdZ6alJf
CGBGLnqfGpEzdup3DLLOd8/JZMzXXuKXYkfHnwJnsiUHejFrhLGirk1yvYVJxiSQQBfuCxsmbckw
8/1HcuZOCiiA3jW1uWzvNQhHaiZn8L6Dj4qY+HEltExEbYpclwkYO4GO6cLM0XMnw4vBh/9lc1+D
wYaT8+sApXLdiyVCzI+SabAKElvAnRZKpfHggKba7j5mkrPpQ5m22GB7RGt4h+6wPQ9Zxe/F6nrk
okNpa5xmn7C6qC0sOcasxyNhaI1aENsMt6cQOauoz9y7tTQM46B2ZkfC+iaLeXiasqqlozXgGI26
wiausCMWu9Gt4uCZ7dbb1SRvcakCuYt3PNH7z7Mn6IOQAOzpUeQdMOuARrEMoyMd8hONVLZyXCSE
Zenj/NAkNWVVH5kF/PaOGHHdgklK2zds3dSpa6FRzvcIzlponduLrCpwArQ/WlikHcBOmehISrsF
8h7T9y0mPa00WMYNbiDD4rgNXz5IGUhLNhFhJv4ZAk5fAklGCXeq92/eJw12dZXiTxypq8EOuemE
Qqo5am/nhS6Gzzd07ldr7bwux5oQd7aTP7H7QdXcM33f/m5C5g4kGDlEODg8bBf9tHZYmcoKAXcM
/kV5gZIHgbWaEaj0MpB/PGGDodFBxYFMHYjjpyM2MOqQnwfhFjBBCaeTm/hhxzoQ07S+X5Y04Z4A
/Tt5Npmz1VkDGHPrhbngKW5/8cZkwe9PH1XQ+6CeMuDQq3evDORI9wuZAOGbr3Y+Gu6tqf+eE6OT
W6HCMDUr5cHVuC11sJgdff+vbC2iPZLvz3AZpoIdxAOIs+AytKC2BzGk6obCVTmXEbSG/vGG3jtP
ZFdPWe7VEk9b0ckutjkG5BmjiJ5BNTjEfDq41Bs9dUKuWCzsH/UTQEc6XlMrw5zmiEcRNvjhT9yx
8FOFryD/F5v97Y3kuiTmOIPTXU+k9TUt9b9Z8kfDBHbrh2IjtnTemUxC/xepfDxjGYZt9U+tu8tF
NG4oL2+P8pN/BOUM/3FGybpYbUUnC4UzVDO5ztSbyBnfYSPhsGY/hbXgo27cI2/XcrkjpbI82sOM
mf5me7OdM7x2cOjaCvnX6MoB5ihugYC0ZfbUEgKlyTFD98tURz8OlYMsy+fJRgziVaYkdsuWd94n
oJ7vAd2eezKOO3kroc2Qw76HCpfKn7r9oSzd5Z39Uk97THLXoYx31T55Ei7QSw6eQAy6RNLENGGS
l8t13WbJp/6hJk/b82jJ6OHZdjkXQ+btrnCcPKJHDAGjTOYmpLTqr2Bt1FhxJgLBsyXbsKN4V19V
wC6qJx6Tbo3au283IjQms85fMB5qb4eOSCOnShpLmBQE6/RkASXIcbW7SAmwbqr25ewterG3AeIc
Ufj2Qg6Rw6JKAayP4XpVIVJuGJpB6rAihKoEQMZfP7HMk2ZYc0ScxQvSuFW5VkStUUWHJh8TN0B/
PxIzThIHyN7OHwtDifwH3F8C3Z6vEcuJAkqul1r2yBcei8rTlSgILYiKBtlSBPvAiHX3BIsNznoc
E5pifb0PLV9YZJOa0mHk0PCdQTNUom96RBYNBg+McbjKLNao3Mp/UspxNq4pHWYBV88ggjJbufdY
nM7ci47cdStnUWiTPudqDPWL4+6yCK0DVfEtAPnR/Kur3iG2p/j4+VqclWRg7wbWOUQtOtdMDlw3
pqM/3DxzOPhxAskQhujEE43IWFEAHeOFfadqY2pmgVG7XIuDgfEzrCc4GPSg2RtLGg5ecjB+Xajv
mMySP2bAa0ohKaF4f5h+Ox+mhQYM7zsJhM+UiMGAjyud93BwbWCXmXBubGacMIcCAEPdhCkgqJ4r
GZp/IpB9fj182fUx4qD6JvneE3475a4HkNSru8B+AmMCm9k4anOGcWV/9I67+f/Fy4b9YrdtdZdU
XUzHa5ED1atcD9MosIXiTGPxSkrk9eWt0U13u4sfJ0ROf2MOcaS7ogLpz2FAYOiIf0I8bAmD78r2
ZaDmnTn7zpg7O+OLjKCISX1ve430FH3J0ymOd9NbPkI6vl9p8oA80lB2dKcV8cNrvfxZA9oKtiNu
xXRF8xL2E2W6U5JFXtG3PLNTbd/ko1b4GekEAuS5GUeGI3WfUtmg25lPGq4d7DyqqaortuIYoIAp
uBNIhpxdGOvRLogM6N3gNrcCK++ctXy81WKOv/mJPAg/XKImEXCu4q+ETLa3X/4+RX34n9nKUp31
NhXExWgr/qjvMm7BCMdWonCDyObqi+irSzJDvIWhXRLuUzir3qN/p4OVrc4ELC0xBVYiQ5LgaqZp
STJzEho0KDupRmOynV7+BSeDKOCfqk7RL8vDqmZKwTYIPtHWB9fzh7Z6xhAf1/fVRzfMaOl7vFma
4hmL59lTdXqfhq43mVVUpfBU0DPUVmjSvlDzanE7g/yzI8xUs72VTfBH24EUcBvTGQe4ibRryC9y
Eu/q+rsTR/iOJPLGA0jvy6NCV16z9+amTEJkxs8lWgiiPjlM0VvBULQDj/l09+zdQoxqUX4OoS2I
x5LSuPiLnXQiyZVzVCzA7xRgDfaAVT3ePrWs/WltIY9YBVgMk/WVDNkGDxMWk8L9zYkHrt4a2/YJ
oet0Rmnn22dGmOmcKMa/22eNoqh7lxCvMAc8H7hWuTxLmCugeAU4tYU07dmMQ08waHoTcex8k64R
EafbWpRq9w9s9OsJesTy5G/UdkAUiBISADV+WUa1USIDmwj1Ky5h7QTBnsMOXqCdCrVd3+E228iS
CJs+2ZLwcb46Iy9Pl3QiqCYTWqZmDig6LuBZ3IlhRFHAPxleuw21IsnM6CD3NHtLSNycLoMj3+6u
4nju5LUM8A6w/Z9eDo6eez/2OGuatInHIXUQWbvnW+jg/S8d22Wiv3i64CYjgBHF6uR9T47gwMfj
buS6cjrpSmW2ASxBCUPb9IE115TwjD37KdBqMKJGIKVtvVoFYu25i6lVFzADuP0I2BWqMFGW4O4R
ERFiqqcF2MIqDUHIoncciUQmygBpp6GatV1rLT5HLdydgvLwnUgmoxlv/YEQHFlCb6n2cE3pGZrn
jtvJysISGvR0gDWGnxhJAHvlxqwCcF/KwRz4QF4Ywy/vDYSUIX0qAolgSY29GBPmZYgKDylo/OuC
xJvoZcQ+stS576u/tpLr70l1Te5MUE1zOdiA/J1Fk4w/2FeKmrbJIr9/CTllSvK1F0p4tWDhMJnH
mvL7SSPcjYbaWEH0nKz5f5WAc21Awra/1Rutg3CYboPjRU0IFN8ktHFYKSiVbYO40o7MJayBnBOC
SzaV1sus6wW5RLMxuY5vmdVDYk/YawIY5QyjnJp84bH+cx699SAcNEXFFvakjiYHxZIbywKjYYXx
aUnE9zBUcZJTxxTyHP7nH7ezt9XY5gCUTURGeNYaAEUUXipuFdiTdYUnHTHKd3uQ5vkeo0AAkRlA
LQMz25XzUplps/vlCOod7my3lf0PZoe2EYY3KsmbHRvM8SLsuuvdmsEWqXk/8SqHUAI3G36C+rxd
k30HkFQx8V7fjUpOZzVt4R3+5Vixjwlni1qUM3mCKNY6Bun+J/DLM9FuCBpwZugjJ04P8ak9dHW/
LHsky+6p8/KnzOWcoSd4ekbFvpQjuROOxKp3ILuVTXXY4vtX6sagfCeMFdADW+iu1bwRle60644H
ZVmK6JyQd3Bf1UpxgxSstfOdu4IO4mTSKOwFZ2FJRcCPDMr4apO6OPDdxykn+PZjrOdd6/+IhBkh
rYgoYhPWu1T4KWMaQUmtpCQLLdEfDSrPyTvj+9cDXANq8mL2BlRW1Mu6Ahaheu8XTB0UTH9gc52n
cPo/TiG8SpPoellWo/CJ0T+MxxTE0tawRglPf7UnFsQBowrgH7fmBL9fQ0k6D0MzBxnEn0z7L2FE
zQvBXz33sCbZTNSC4/7A5e7DYNSnxzJDt0PKg5vJreiqPe2++vcHikYM5UCrY5Egthhm3iJ+UmZD
3V1Pe78t27VhQTNo9qm6aFwWUmJmMYtBv6cnw4JmgNFo19WkrJtJVWRYZBD5Sky7NnfY61FI5yFw
SEckWqTgz48bOZwvmQ2axLFQgwrVbcVaLCJFldmTnM4jU7Pqk9jM3+5c/uygXgkesv9qwJFR0Oxc
BxbIymuprf0ZYkUjeRq6ocGx3UzU//QIEl9h0OdEdhCHHP/eatrA033rd+qgYKQK/xqq7E0EsFCP
Si++yxqjhrwF513UQhZloCJFSGAAHPAKcLJmeWkM76gnO2G+gRwIk08YcV8MWJXPUgDftNqCnPd1
lV6TyzwiNT8chtLE7Xu+BpQXPNK0iK3xK+jMbH0yUsDb33WKzQUbIPXYKgPXD37/s/9S6MDAl4La
SUXYl+EO+D+apG+aW1Mhwq68SDR9dsTdQoPtV3Po3ewyxvFpZY74Ml1pRC1Go36xyQRsDT94PBhT
Ytz9QHKBLfK6GfUDkz44lIXp1vwfEL4F2NsdZe7TTV+Bg3D8Jw97XtWnxAvFGrlRI09GVKD0daFa
5ahYpdE9kaiOH1r6EeO8EoI+5yI33FzXCL+iPUdY3KWtfsI6baBzyumP3GY6OpxYmtZd/JSKYU8H
I9q5sGu8Gr1cw47mvjikmIxKHFLriCG0pXgQaqedcdHqo7uD++U9Yjq0kT90pCR1fyzsgwqoEjVR
rbXNQR5roBKcDAUiSC4vbZtTn0FcM9Xj555+/+7wyPga82gV2nNJzsa6iZIIiL0U6bWLwKRd2wxn
74XT8MCh/9bmuvdNsFlD2gkBIkWUHvARnuH7NVSs7ovXCYsE5dOpwgdVWUsWfkOI43aMVdYe2TgX
U47vlQNTDGX4XAx2XFwCRT82pfuxJiFUXoAAtf3EAZULB7+W4KEQptWXphg0tvRDtN8U9hxt/BRj
zjcZ0RR2o09vaXa9U3tjVIVxa3scwZXNRHB/Z8s+02dhhrqJD6n4DAwFeJqWenLoPSITVk4ZCefd
wXcewZGbr7Vhd7NBw9oTzNWZl4bJewV0EsBAcray7tCYooj0/uXu3YwO2eLcfv6wi2x9kPxSP+0Y
W6NJ4Z/fTNgJFz1KO47lTcAQFB+7vgZArfi/biSprYxzBAE+6GLLU1E73UGAOIL9mQFSJr9yT5qi
/HbjD5DCQ4n3xbARR3qy61qNVdOgT87Q3e4/YG+AQT/9Bmpnx7GWi7y7pJb6Gat/2FYwV36VmE13
WGR8ovC0qKwTkOtTc0hrowXXEm4bVBtbSe/y+WE8YzKLvgN1hXJx8DT8PjJI6aub0MoS2EKqpR/e
tOFb4a8Q2AiJJ1/e95d9o5ce+JEfO0zdl9h96cfqLzSnDZvHjpwR01Js24Km7WUhD+ql3uKKF5a5
os7GflUs/mXKef5kp75uFo9XdXI6w4MVUjnSvK367CGKFRsG45gy3S0i3uQcytGwbbwEmTht6a2O
6prPo8VZsKF/lmBUsJ9WRZ4nRRUpaN//aI5QBVK+a1aVRYAej7cfrYtWCGW2H0kLmb+TdioQKjMw
GN0uA2OfWbFEIJlY2t/pMsGYhj5rqvBL+HlXqlHtvg6j9GQA6qJraTM5nCMVu2ih66I5zGbKNkMB
IEqV2M0Naldn6G0d9NPH+FUv9FqmbiZVoCre+Y3Ya6F4inpCHhHM/nV73Wqcgh8nJj7tXYMLsWdA
iveo4EW7NqAuM58VFDyL8FDdpRPKwMgU5/cosxbXU+m7+RET+ZiNlH5lN0M1iV/hRi6wpJu3vHID
T0omKWA85xPF1jzH4/G0yFoYli1cLiROT4aZ0/ZkMUMyCu/A1GMHpZhEYEu6H11wB/gXom+O/lxr
5BLtreNL+Dpk5dT+GrSlS5J7Kiw7ruWV9PBbMygvSrDsefJTlrxHFyBLWF9wL467TIrMiSkbRNl6
yblHsTr7SVJUw7Nlmtkj9bGrUztYfD/nkTPf1Wcbd7jQAe+yk9bual8F6eZ4vDR7rbYcncWvOa0X
4vLIngJyb+ZvgNx/yC6GCDuZ2XXN45ip4hzGHSEqno//evs73dAUe6S5ty5bi8oNP02CdDOiauGS
ddr7NTeHO1S/Q5ndxe7caMLlIMtJmhOPGu5NfW2eckcGcWAYAqI1Jb4ho1VJ2d5REI6jvl9TBtyJ
1S6xRAQBjI9jntS13+rFGCELwv7gij8rjXKuWrdPt4f2EpEircLDMKQcIG/Ay1EmNEsn8290hOcs
TpasULkf1ZNMWKFboUB3MAijbbQGru5E0gei479Gf5DM7ciYsjkFLjbauATsgFdnNFkJkaL0cAwe
kxy7a3H3n012ybQtcYuMl584ANg6lJ7+OzC2Gmm6J2fow/a1giWm5YYQK4KlZSqVFL2SdSRU4qTo
hp8izLePwWY83+dOBzLurc2MYwWa1rlCFCIf4VznkPJd23UTQj0m0JEYT2ufG+JhObf8YBYNlvnw
Q6ZUt7LzsCbIAkVcbboorGvAditXyDHJ+EQOFZlvQFxtd78YeObb2dSxGDTwtL06S8APMBuQJJfE
hN/XGmMqwdazDCPZ6mInWQWZvGqqFztWMbo3sIu9siBGg6uNAEPFqPdRxOPC4wkXHRxUv2C5jhje
tNC71jrhV4Go4HTAoet80WID+wNdyqhFSe8ELuQ7N1uD/yUChankPSKMOoeUIBCgUc/QBNc1FsBw
0BR/tRu6T0+kO6MQ7kAl04xTAOpPlFd/ZyBmHh+nNeMat024rubyKvx8MTp59Ck3ucUtWHD4jmlE
+KVMrgxRC/fmz5NwgnoZVfs0bBCRNeUaWQtsosb3jnl8bcawnC17qReYXetg4H/Djd2ApGFVuRAL
7w2jXCRtQkIZ7WZAWCxfPyed75TvtEaJclG0KBsqr5IRWi4MUWoMnM+SKKV9RJ/hnR35dgg3Ltq/
rFN4Cx2enk0yuWR5jl/vrXOAPKPAdEL/9K5ZWluNVTc7gBT0VV7XAPgtSxmPXDXDQRjtpOeRU+AD
WlFAijnG7u8oEC+TqTiR6m66DTpBFscWVxPeQJdLOANezA2zQjTrEeYRRiS/6tVZqQi/Mw0d56hb
ZcU4TToXCuzfURaenw3GQiZ4EcMhGH8VFSYNEJzS+Wk3qRh2URGcEbkB5+ykZ/RnUbMUmHyhVk+c
hPsPaaFQuNhmGSBQFYap1JhuLQ1Epb10wkXzk/hCQK0gCQL8Jpf7tDJWA0UArFPnQIiXV3JrU5rZ
DOaK3OTk6i2n8ILpNPigfM6AtTCzbGoWK/InjqAlc3UCcS8McYyofECYX0ckBJY1R3oDZIzh5/eQ
6tI4CCNWC8BcHAVJJtSl1a7Yen8ct5pfsmBGmbuz1s4ifDeiGsrQ8jX5qG1Qj0sC4qBWTwpyzGur
/UhGI8ELOJ9xfPrWXU9Y5W+FRPTUgYWUtsVv3uSqEUQ7uOlknzyG3K5OZvfiduJGZiB5oYNLjzZG
/H+Pjz7+9P6DaYWM20qhYs+NxgW0qBOwiPBUn1nFFni4s81YPJiTE78gcBm62rHfwaeqMi+37v4S
Me9XVdPOa04ZJU1l0FqCwYxoi4+BCn5tFYJkSajzs3+Op3do6sfPj5Tb2HYzKt66rPzFhdhI3Vf9
zJGipDJFqX+IRTTM74r0LTLE2uU2RmRLevabJAQvbceSiTE+IhLZVHFh/UaFLuakug5SKBirzX47
S8+car2UluMx/Obz98ENn91q7s5aYLGBY65hm+fXNfa1oCXdXa8kLns7uxgWcC4cusrmRJXd4SMt
Rnz6PDF3gInxqlrdjwshtPhaaolN0uZHs+NOwsjKGM1CTMJo5tyyyZWGGULA2tr29X32OIoNE/JI
L4ICYQwb5hBw9TeQ+cOAMb1MFXSfgPzvTlfkeLglAhra/H+tdsQg3kRGWtwH7kppzz2R0cxajseZ
BwemK1xGYo7HCkeE9HyW/HI0gar4aB9D50nc1Vy6qK1UxC5UlaMFSKEMUyrKn/DrdTGpPoLA4gbB
1zHv/VXviW7pKI17EEEj6qkYBzOXPcTh0dRj7e9BkQuL0ePxQJG8KuDXejV9RcTy4Foeg1OM29Ns
08jOPs5sOu1h4DN8mNvQox8KPXjdQ9vTkJA+Qsl98MPzOgjzqeDNFw++aBI9D8ooSrugYTnExvUU
dBrgagqE4ZQ9py0QDJjnho1qsF+GfVMycxf2DSZ/JFXiTMJvWU/nBZuNpFNOOJmWSHR5YJ+uQ4FL
YqIJD3BvhzZlwsAibWL6Kqg17+QPb5jkkXTdrstx/7lfRHMAJHXtw2AP8g1JJvu+KTYYiEniNea+
Yo8R+uSw12POEdFZPQOrs4R/8iNq+xCxd6fmrROlhfaWNJkX4eDCaJK0k4yM5Im4+siK11a9paVU
aI6kc+D1uQV1iMeQ8HaCijOZix6oo5mnaIefLY/Xq2sHIo9DoJXhjvYjLotep6RnjUCRT+/QHYvV
Ei4hnMimBQ8q8/Ar4oYlRNRAxbi6I3qvd4rYMCQQ+JdGWyWjFpz8+3Dq0C3VNYB3YLhMgzeVFRV7
gQ6/5eLzokpgMRM2Au+8AVr1ewy8TkzbAj1ackAsseTjPhf1Rjd3mjjPGBMfxIWVilZV4Vt/E+MJ
pNDbIirjdLIYdqtYDgbjw2HswXYGu8nHpOAcCnfDSIVfCbrh0LlaAqmKb6SenH0WqkSs3925Ud7c
i1Aavp4W0bxHzzNqfagjFXMhI9+PJS4eqXk019q9ijgVYhXxIxSS7MTFogIAF0vEabNusBGnazhw
0mvDfzzEUmb5aXxbcuW41Jy42tv5qiZM1Si/AW667+5vpFn6R85Va7T72l0qYamo0Fci4Xt12OQ3
9Cw6mkbNAACSPyFTmU5H083kADsuPqyJfLFMCPwsYSclIt2Do3MNghBXJ59ovfKiQE0gtUbnnfaS
cTAEV+amCYF82dy5LVnv7GV+Babg4gIDmFsZHPRd6/8HIiw4UgARyVY5lqLqhAT0LzYI8GtxzXvv
2rjiJR+Z6s7hKx2omoSM3BZaHBbgcUG4b1OouRBKgKfpT6ZgxzabxE0FUKzFBShL1O2dhqwoWH1T
M9SxLO/Kcfx8dRDG6QoEWnBXP4z1lilSYIO4LUtE1B0xt8BRoS2dzLt91MC7euAh5jeeoQEag2g5
R27UfmJ/8N4G2TMRnoKq0HaTI1T9q2L8D1CyvMHnPHx+4ffbuVInWAYdwg9+BTU7jJyEB9oRSOAp
CVcKiQtBKIlow0/XbD+5ux+w5vO2yuEWPCbTALcPtOcdlDLg2bjN0xlrGnQx3i0U52/rdesMso2x
KpH7gRBSciUQUn3tM17qtWxAmchgbuyC7pEBeL5c2gyoupTux15XZLvMGH4tFNBO9iFA5NJFR92Q
lk/TKkbQAQyzGhvDBw+oCrIHUge3PpA8SNBeaFb320r9W4lkgzFMXaWKNcTYogife2JRWWm7w2vh
EKKlOYRhA7o9DdG3eRiPYj2ZSm0QhYRi+JOMClz3FYYDkRQm7VeQjfNL3oXmYbcFkhBkZ/P8WWRZ
eo/da5zChclBM6AY7DzxUkoiHqyp8xLVj9W6ELwereZz13B25Q9KY+fcgO6SEl8JGR3RK9QlVFOZ
LdPbQYqqq/sKIgyG+aPLx9rT79H6FLOi5zJbqAkRV6waf1pUfyvmc0WzHEteCbfmC8P/Wwv3gox4
AKteyFN8AJfeWpIiyPFOvW4nDcvgBYeNBRQXC5cxN9qlnug0f36mCFz0+hSJfnD/3mNDnTUFqD7e
9aKSOHo/oSgmj9yTMcMgsVGKvhwYVzGv1zmbF0VnfLTzlD2NeWWgy2LaBRkbHIR74DPqhYahw71B
kTi9qufpviUHzRH4rpkqZlss/NsFf9aujLSHyiEZLi8xLXGdPL+xrQAouxtka9ikubnlVBW+htsI
xwAIXS01S8D4lCUAJdDlsJF2RNyrII2KBEBu+GQSN6suIwamZ1ghdfZ6NBBcl9alrRcYzfaeCkzI
/ZPgPgx8Ki63x9y5eCUqdVuJN2+VUpma08NrU20yJzHF7YxkKEiBF72KBHo0LHlSISREFngvMuI2
qIyT1iePHXNRxeiUAGZH6Y2xHgjAB8hNwCEJPmcF04sUbD08Xl/FuRC5+WsgXmhxmPYCo8s8yo/j
Ws7pIBUqooou+7VWYkxSyo/uyRU9YC8OAYB1ATEY2wiU6yBNieSUmWS7kCm/dAA9j5LqbrBIEmzZ
noeVGRwf1Hsl1VVLnbxn/k1bOHQ6yn2DduWXOb6u+I5cuHPEz5sxbMoh/oY2wp/+MUkwBidJIlXX
Hf/B5I8Ekp3rNy/T7Tyh7yQCci+4Lga24xqnYF5wxj0eQtS6X+3nZvAJnjP8bNlsWRBvAmKTYfe7
gJIRRY/mPtpFJNOdr+XG/ZfdQsyWQPzuUlMrVLJ6HmPTd/Yq6CO2UycMmklnK76AuSEqoQL/XXaQ
1886YqSd/U2B7elWKEFZLc0rj6CxMMny2GIiWlmXkrxu9JVuy+5w7hwMhfZH3IRgBSXdOjKQ3r/y
eoxYzYyAc4luhBBlLrko7/+5K0+TdXbUV0lLV5Gr/3fsf8Gz30ZSIbx5GkWu0MXAaTALlPnZE8Mo
u8/1hi+tTm1y2RBtUrJvViaHsykHOnk97R2dEKcS3QTGvKiPPdB4XzfciyXyWJKUp+jB3gQFU6zF
MrwgRDB8jD73TvlQ9ifdlprF39NVAxP3gfJNdIMmCC7SI+vc44dfPFoPWVtX1O2TSkpmm7N256f3
LKprwb8gQTu0msIIhGXHP9nNfz5lIg5CpD9oG4eE6Lc4pkGLuTtksO6XDKUwfP/FOM4cEuiRum3I
u0WiHODh3m6n+3C6GdgTXiNz4SZnf6LiXmEVvALBLbTlqD12UXxviubwu8KFJ3r630etc2B5UgR6
3zoz2Muj+CxvvZf5FDlPCRPdhAc9Nx9A1A29rbHRZxDlXOvze4fHvH5yesC2DAreFZ4xWHpJMmnX
A9qiomZParoSyIpFgGqjDeAhfpvqa5OY3uJMCKQ/Bb6RIu4tuNzFoss0rn5SHtpMY/yUQzn1fjSj
YJF1OjESiAipUC9h6Sh6W/bMvTRUjYKTSL1DsVXTxdiy3hQFRb4oOxXiEJqrFcMmXPnNQXFDJaws
qR+P0pAMQTW2C5+WCaWMNc1OyHTXJFNWQHfA/EG1Z9vKCaWWQQKu1bRFXgQR1+jWIeBkF28XH8NE
DI+8Mcf1ZqqT8ItDMDHEHo38XFo9sH5N0bby5uozWJje/+zFjUPHg6rKttZlV4pzJGBxPaC7eUTJ
C7noskKsjHM7NqhWt/hl7MkHIUn8avuNHLaD9d8rKLPLX4pbPCG7JD5Knbx7Z1Al5Up0pVMN7q+n
bIn7QS47Ksg2rv2c/i7HjZ1P1Ku3GMpZyBOYP54PAdsOtQ3XT3V60V6BvEDApfp5cky4xlzpGTcp
wLplLCskxdAv+2q75XaW+WE2A1NPEGJGXP5Ar9FR9CLMgQQTaTTDiRzPdeOhtX2UpqSILvg2YYtT
1W2zjYgKwUVgyDvYeBYihuva47/0HTrr9kuwA3WZspljHS8hA1mm8RXbR5xUsgBBpspckMDmtJRE
kXdKQSDWMCtXpIGI+L5zwgkP5nszgdNsuoSknK9JDlR094z7TRxTo5uAoBDLJdRzQrUBIYa3mZX2
nGknA1dzdiQ7m94hq02S1QtR8iBmbn6+CAZeM6Yh1UuRSUzSl3rwBvD3PUh61z3Fj71u+IrVY6zV
8cE5G5NZgKuoM97a84gRf8BwCEZpBNhfZNyc2aqO44lLzQu6t6dYKVLCzw29uvQMylCKW5qGSO8a
DL+1CfZYH3tWUFvBurfNO8QkLK2CDs4svtltjVmrtN8EErdvlAo+QbPeSJaKZ//WJjtcs2YwcMVq
NCI2d0MvsjZGacDpTU6hDJ40VQ9C1MKZ5OvO+sBFP+zjjRgHISabTDM/Hic+glmFE8/55lSAx+HZ
WN0jtpLioAaxrYfS8tb+5jF6y9kk3+Y7nvZ2sjttPtsj5u8Do8dVw+Y8QOO2/nnUVx81CK01gvXj
RPeHuON4HNjCX+qG0qUZEJgUhz7jNroLRWL771zCZBtlfxQreC6mYW4eQbbnnZ9uDHb6/evt2Hi+
b6dVDOi2Xb8k0tx0sZgfyCWLgMGpLyZbOfn37JhpP2TRmJLiu1mdu4AwmkBj7b2j3Ffge3oMseno
pr4wpQN7/iczNMpplxIeTVptZh6cTLrg8+CqfCN0/9e5iW04UtdBKaFBx+xvanmaKx+iDdglZUWB
9F+D9YMvR4MkAYiqmHm+ebVTOHrJ6yBF4H8VhpAQCXPt45+5xZYBsIR+gY1+NieSyLOU0uMV7Bms
Hzrqrtpld6EKkxrsViWDOQfX4KirpKblOyyfoo7c8megBGPte9Uj7vi8DfpzEIjjj89DErABtI+F
ZQ2Fn1aXh5w0abKEsugoF0Be5GC649tQ1EPnWYf6eAnXhBN48qSAlMXxO+HDwC2kPgebBIMVwnoD
NKm+jf/NnfD63cDPBXKQygFhZ/Dgerc37M8PmwZvOdsYUm1khsVCI9eKNyQjfJT4wiGpgbnF9TsU
+/0gWyYKDz/YFEN97pwB1z6Mgit0kvdJotwnWUj6hLJkaf4evU3PpXMhUKtrikdu6Lysl5t/dJWn
nOcxcO5vAWaCT5mCg0obPAnEsDzrVT4Yfj23FSLXKY0YA/dDywlVxL+I0OJsS2bOTguhk7nEryZF
i31s9HkT537ie5G/oh0KG7E0WyTpTvYbVJxLGJ2E1nShRjI03xs3HCGnspYl8QZbEhg3zDQu5ReJ
k0eaPOD1+yHP6rgMjbI+ieD7QhTV8wQyqcbCKHpBXxXHCa0epeuGkKu++pU3SnXPh5fdTqNt8T9Y
SUHp3wrEaqyrVZhlIpKt8Pu5PPXX+BHoP1vKdnkpApX156ZRz6kLlUN/1eWNOunorXmYRzbFuBbG
pFGmT4giGS4GqYe6/6H5QQxyUj2Hlt6t/2zJAEGWY1h09nVu2g1XokTP6Rye9/AZYbm4syjFBK2Y
sqin+aM5zfNrmchs67CAmDbqnonzfEvZWEI/rlbECOlDK9Pw6rp0TiqesDPbrgbBl+IQbE5HPDRb
K/yi9IKNyezX1QsefU1L/xItYp3KF8ZLnWaZz4YajDv47tZFZm/XffX1NraMj8DPfjWFiuGih5fQ
ca5Nceq3Zjr+JPF2nYFl4gJMn/IJqX7kzY7DBM/JrNE5K6kDY2ZkGDwn1qMCad5+3Sx0gJvhUUzo
bcMTaJKViMolW3nplMuvdf7mZmglSHcMJekuZjnqC5hkBB75bC2LHoTJcZQJPmMe+ZYChuU6xMlm
ykNCHj+mLKJPGHgjjOryrSmjBiYX/R5/HCRLUfIdsN8kEli2+wri/IHuFIYMUYjXMa195LLLQ4lh
VlNndHXQYiu+VDLfHYJgOwJ9zuGlvFUiYRSK9nGvOUsZK+aNiSOsxFVTrMgTmCr24hnrlSSOHj1A
gI2jNvsBac/gDst6Go3qmpRpNJsyRpCD4Qm4HaW+nhAy77l64FELG11xPAR/ljFVkJsv+eEdrArN
aTvKuiz8QiaFQa+HHaGS14sQz+4pGFsq90ZiPG73Xg6YAJmgJkSVxBQsHis5y2L0vilWSrwvTdtv
H4vzL14ZsVDlg8JWuKNpyBN30RAgOEZhOqvJZUXvldxitcjQO8x25an1unyR/Zfmjis4xpkNBa6Y
XMC6K/K+6XjhNC/xYgUHpy23QoI3vt28GOJhEYDyYIIn7IeadSsZukijuyJcsb6uOEbmtga860fL
uon73/sCRWY7BuESrec/T+mjSCdjhE8imjmcpyo8cnAeNGjJ5/NJEu7Yxcv+Lg/yq3Nmm5o1p8xz
QrcPYUWvc9ytc1NsT/l+SXp/Qq6uKkGUgY7nyzDKZQcaF0uvCGaSqMT44CwQvlOq1ejllbC7Gr9h
tknCowQs46edO/c4MJecE8bvhdLz+ScBw3UUxDSrC1aAbYIGnz7qJdvdTlqIEw45yOP/YD048xaw
jO4I3M+SI9IIIUT4HvR9ev5IM+6A077y14Mt/K9M6YNV8q7f8dd4IkFB0sguOjiabiqsGfkZeUAo
Mli1lSuD2nvq4CEKi2g9aQIwXL0iHYX4a7vRxezOUQPlDRuC2oamxR9YzXpD1nqi0aO1Fvu1jvAb
BKAMUqXdomWOVkecu05Qx1Nm0enjgXnAkS775QGRpZLxw6BNjoioTvn+MArJf/EtzX/rDVs5FBXH
Sown5KTcoZyT0JMmFjGfvXGyIScvioixgllH5kUHCagi1qw830qD7GXjXs1Inbi9EAONxwpFHAIC
xMi4M+Vx5PGH3X9xa3tfJ+qUHhDEv6ilKbcSLMvPdQhDaPmCa6sq/+RORDCrJJ0EbqOTsbcz2DTW
lQJGI21YUFezySKa6//ExyamHBUifosUd6OLRWp5R+WwZmmx5xpRglgFo97/t8dY4RAfdW45AFmm
KS57umF7A5JMKSuZuhMFnZGmGbIauzdyV952bsD0jmKZEY1jLH+gpOaErKgRxF/tUP6wp0SYZLN4
7KALdWR0+oz8dzvYp+d0zlyEQyFWk9dLiWBePMxZnR5wIJw9w4SvAc+w1MXLafaorn02np7+Lksu
NUvdS5hsDV4F3Kpx3eo5ESlb5nKTwBTCRoUjBKKdRM4PNR37hqQhtdleJwqouyLSz9QiouKUh9pm
CSq6d9IqGAhvsApYjI6EkeeE+l1H7UAhdmti8RZA8ltT3Pk68yWJtaUqXBEHmgURIHlMKboI55XO
yNJzvjUTh3klf6q+78eIdcgXtl7T02iHRnH+l5pVRwKP98aTK0FVtRQ8Yx3k+ZbHOKP4eIeWwpQy
uISvqnNfYAcU/4SiFOiyLodo2v3otD1S1pu7pJKcbDyx/p21C8FeG/4uQF/vsR1vT3wDU3D8gdI5
aOeISPeYVh/VJgaO69r2E+pw9YkzzyUYZ6ixe+IQH4GepcMvxSwxCcgWc1qpIsGcldUb4+3h5ful
vp7OVNJJXFQe5x8KtbTbrKmmA7AOyOhtkLf1xzsU7CyQXF5FX1qPu5/7m5Sy3/5XSD3+AXnrNo+s
3/jWknTqK3YBdCyWllijZ74qBh5696Bejdeyp8tsJU1K2uk3W2vcEyz6JO5Lj86PcFpe6J5NejbS
nqOLgbE9hAYSW/GRDvo3Vsawcuw8knV0xuTLc9u9HuucUKMtERt9LevFQNstqDXZCrzM57NPG/lI
E4S+rnI7X13KRuN5toUeIMS2V85QcCRI0CZdH1zPvcLr1NZctUqzDNdd5kn+6oy0wbW2/UF7QnPB
5kg+7P+366FysZTWLXSo+SXKv/5g/AkA4BWf/Cys7iaWo7YGCnBlmdLn5o2uIoJ0RxYuKLhkWuNm
Sb+BhhdZOohbKI6txdu6r+23r1G62FN/tujZmRG/2dFlBIN/v1/WRh+kxvDc4oOKxXs3hSnHvWRl
xU2fXu9aAsfRZ9x4Wwc8L7GWnZxTVpTJ8QzV9u5QVuqqvX48FWQWzAA320TXBYEdSr/FSIFUC3G0
bYx7KdpB2LuFoeY2QAirr/GjthpOgbTrbU1BhMZXr+SMw49rDZluGiAF/Z2tOKzqOQWbihww+8NA
hhTpI8hCg6xuXuaI9Ej2RobbSHxuteXoxQI8ISp7sNG3yFose7HuvnLCJOnMtJfExq5NQtx3uvWT
XLNf5g/0WKb+jCHCP7D+NO2FQ3Mu/CszQPJY1g+gzAFO2tqFA7Vw5+xJS4UBWDMxAcEH4/DUE/Xz
3SzsdFp8fH5ADmD2i7WzCBX155GiwQ4+luLCgzTtixZx8W/tNJVE0zq6T/cTuk9IMhLpntAl4XxS
dlrtBHMbrDzPHb3bwN9lrtwc9rneJd8BhkXN/CwetaPXlgLz8QtJ9Hh5UdzsWPw5IK6QJu5S6vkt
yTtBLu+KQ1zIrzASe6DQo7wiV5aCiOMcF9PoXhqSPTpPqpjYhqeqhFqh+Sb+iqPU5MAFfiG34EdZ
ZvklCPWGGQsH1wa8hEcEwx2Sp0Q+TSy0XHtqlPnF98JImu0V0hwffOZ3bivns+MyKNve+V0/bexo
23ZCNZxijL8qxkSinkDdtX3359okUjq1nZ3G1gqw8YGclwj2IQEKAdQ8Ifhsji/Q+GPFi4zjr5Ni
pHmKgJXD6EiaFNOMlhVgjr0+P3uVhGlzZ/Pp8PtsGXX+4XS/HvY+nXWlKVJ87kQUCtiYtV4M0lLZ
80fAXH3/I+Scb9BbzCLbFuxDjjKz6hY8frE2EnDR4uN7z/UAXFR7zPqpgT+vV6+T6m6F4629syI3
0ow1p7CCyXwkFjOIy52c8Vk3wNTtSJ0dRc0CW4Ccu+XeHRj/V8/Suo2ksTFOD5zlSIyunAd6ioTe
byhCI7d7lqiP+mNMFcD1VnAR9JL6t/8ETvompmSSRuNJUU1y7eb28+WwXvsKfYqSHEcIMxuvvXyK
UEfomrZQO+6YuM85q3pwmvQT6gQwSZKSHseQrxX+ZL5GxzN9ue/DWUDn2aSZmUpgK6Bej2+elKMu
U71w2z/GM13joS4A/bFaOxNelgcxJdY8AYzfqrEgXv5AV6B54i4JOgBsiI95+1DwHaktbBV2h5ZH
7b0xOSQoArBxjf9kcJdEc6gWBjtFDdjEbYi2oj1ozq7wqhLDm+PpXoMVZc/18PMN2qVQ4PQxY0OF
xDZoSJw5lLGAvkxLxzdx0kGTPQ/XP3Fqv6JZCcZxwAWzXsJFfVZteT/BzQsPmvZBJXAiyP5Ktt/b
khOH6kWZGGVdxoZUFWLAtH2LkCPrVAD4/d40DbRvWVfC47ZtIFLHyqF91fgVhP9oANy2cFYW38ko
TEV3+klbiqQyqk+t4HVpfJ1MLoqgL9cnCmqpHm0hMGqIVoplJR/JEBdc7tbQ2yiDkbHQvC7NZa+h
aSBtWYOGgcN1a9NE/mSH5Vj5uMGZll3BnyKDarD2Oh5smmccNWOq239a8jG5tszgr1+K8t7fk+Qd
yAGWSipFXpWXT9SIa9Xg2HtbKAiWPIjJTgbdF6j2DhDZPSneXzNfNu7L0AY2rKKGuoIRo5EMugDj
Ml/yx3A9zto0pFxpvybJ7q6y3q0ZzkOiX3zzKnF7azxYXjlZTWaqK4FyxWlmXxKHUR6HD7B8WmV7
mUuEeNeG82qbnpcpArivorKhU30rk/HblNeL2SBnvO6lhSyx3nDHOZIJu1bSdcOjkI99NcbG1M2K
z1Iei5KvFywP/KIVplxJJLPZfC81klmB5OLlNkUZ1IfMMfsgtRwc/eyYNJGxFdHzaGBYvrkLxrrQ
QqN0F/qLefVrONhboTs3rB5OFGCM1efGoYJXU19oovRddXR6RdMSxiInxgej/N4p3h/WSd45IbY9
nGgiHM68AFTTzmJYKUDqRF7Ebod/4vd8yyRXvdVJEtBrVvFf95hcgc/XpqvH5pSC0aMGEm5hYKJn
x2jLg6f0I8adlOBIp29pbL6k5XLFSGFR2FrPrszH0xTDgycggREnTPFUQkhCINLy8cpu/xGOg0PH
KANGDrZagJywJkpc7IdpJO8DCpSmaulKejLupz25dHnDoAY65FsaKa+5w4zkGWmCgaJYi74u4AVZ
WbpuPCXTzR/cF86TH6AJIyW25KeKF5NBhSu5J87t0eNeAvEb2jNFh6g3sMtVYbylwtbYdd/z3Bjs
F+738AZkUPiNlU/Ir8/+6MlG3c9aAxPItnafT00tJPkCKiiZwkugZpcYKFHNKEovdLofEwYb70/l
oXr2D4CyoiKcHYgFyDtTDyNg4NubZ7HAKX0bKyVZA95/yqVjUpy6mttgQTmjsZ3h7up9RJ0jmUCG
Svl7lq74GpkPCtgJexStoQAQoVFRHxlaXDDj0WHwGLjfXB/YHZYUgR78tur2ek0XgGGIhUf6BwVX
uhqqWHhI2501YScnvWDOQ8vHfnOiF+YdJyIXp5ZYvsa+OPY36n+GejtrT6i8EX/YOkQhdOt2ROaA
1PpnGJvelWpjGDM55r3wvNcsNlHIMn461EMBuYUIRnqiI9kAlWlbVHyDVzr/rjYJwBjV+J3FZAnC
HmUOQpPdICD93NDRu7PopICq3YKqVleeVwcPHIS2rVVoZAeEYSC2THns19XnAf9XZBnZzoOVDUUe
49vn9yLdYCT36XI6Q7/u8WXwB3WbFJ2b+Vh5WLbZOOEaVdG1Q/IvDLaJMcYYwwb0LkEoAPww7DtL
EIlR0uV5SLUEfRaJrGUUXLQmCAQRXV0EDXpizpZQySA4wA19MrCrdI0FWSiGjfaTPlv9jgvSixq1
icR7mw5iR+kNMU6QZopvKaAJLNJ2lttV0kLkbS6p18pNa9bD996jEG8qPKUiuR1zc3C3RQec1H3J
LhdpYj0soWgzdJIexo1U5A0c/Q72UIkBZ/wLs5DcHWcMv8d5nfid6Gn2KX7pwTjMf3T9ORNrOwAU
+uldzpwAQv40yu2tlyalxxPMa4PdRZR96/xB07/DslX01RGnfwri7MsZ1AA+bx1brTkymkdMf8Mj
R68ljIKjHw/3Z6Z72c8D/ZFEgvCUmvZwboQnUTybcfX+Zj4ZEF7xkx6oXRIpJauPFbuciToglqcB
IhSVcK0yyovOhFmU5ueiizTKv3zbkKPVTMWdNSeUFwn4AjSHxfDe2e5AE7XkBLijgbZwgaEiFeLd
Q6ZfWNNmSoik9G4tLMo7kTUdj7fM3RSYNddvpmz2C1dQgFuQ7ZTLZm+z/xacwpI9vpTAtoW3xUFb
bDHaREO1KhGKp3dc+fsCtT5FaGqwDMrDwiOWNlAjADaoomwFywoiuZsXzYm9SwC7vtgcE8XFu5mQ
UYjEb/PqcUcUSwOcAxKY/lWEvYLbj0PzIMAa7S+XMLOswU5M25ZIUTO7AGfZiyNlWU9OEpfArFpt
bx+07sqnyrkOM7PK+XfSlz9oBjUlpibo6SEXotDUE7F5cCEvVGuwwmxmBAecOQ8HdKCP8OpBR7KE
TkvHHzP8i4f296OhQU9JWllGD8Qi6YscbTsVIBZX39/ylvU/YuGBmrVZ+3+tzvtmkEMUFho3c2lf
k5/46v9MWyoap6UHOFJ54uahQa53NgBGR/0015hdeAGvYsXd5FnyXe/Sh2YDfxrWId0NULj/to6v
ikkZfgSdqw0N/89gHRaMNCsi+FSKZ05LfalawNAOw6evMhWBYwnHIi/pbYbrKxcgyWqyuyNT3ZXR
fvAb2Us/RAXLFZzr22WAJ7dgkXw6Urubkg5+97Vr01gEhWh60jzveR49xadyoNk9QwzIQCi9OLsl
7PAbpvRJDgYsVkBEVzJJlKXFYBOTy5XJy6jxD08679y1Z05tLOSlOBWnWSG1fZh7a5zxHq1TFBFg
YQdM4BzQEDlkAUH/xjoP7M1ffqOCwOFZsSeQIyXJntgN6nDn1lxQM4Ah8CwBLbG6w+WLjA80o3A+
hHS5TqohwSuP0Rz9xAVtknQGk+IvWYL1WbmFm8yJu3b3KYcF8XSjP2ANOaxQJCnAc4bKMgXr2SSy
6zg2iZdqG1YLzlasBgTHt0nDByja0GeCyK2xIjmCBrNymUTE+4dQuzK1X+X/25BDMJ89w/UKGVY0
mkQwuOhHGY/GEDTY2zcU4pCyoJI9lZExo5z0rbbFCgfFoJZlgyAzdhj0XSbZ8pph/SWLa/u6d2lN
6KxOJrBWIKUlZg91xm8yi8s3mb+kjoBRDVhkMPJQqpCpcb/hOScyfzIEsLNX2O+675FnRUHuMyrG
S8fqSOTMKwjwPJG3nBB1BRzlnYnd/CO5rlulvVI1MpkO4KsNgP5caJKhwjDVxvj2tWPoxEEuLEiv
zpz5SzyjBym9YdwEOvXjQmUGhuf0THCqQYnqibLi6ObNr2LIxuLOqVLEYWgsqu0DEmmO48E9NAqi
aIbcj1MSNP9T1HgHCy6WB9eOqq/ztqV5O0FLJHiE6z+98OhU69OO3BbwsNCWM+ZCYP6TZ1XuNt1c
BLWcNAGIlOMmtmQER8jKRuOfJlCc46fWMLMfveyPzG01RxBO9asChZoE7ntiYCCtACoYZu+Ee+BD
Fq/0fKk11QL8mx6pl3gHMEYcmHeQJSlN8ICmlzH0r/DmlFS9ryKUAUbnEaYbvWgggo7aZ0LEa18/
rkf9PMUUhIeSX3JuodxscTv3kz6LZpmYBFi7k21LjXBBHHmD4IbdV6WkSwE4Xfa4vpSfgtcWsU4K
g50fN54zk7iI94TugFLwpZ2ZBpaU/fs42V/sHLZ7LmsiNSxW02u1uIESR3n84kcixTFaChRF5HBe
RNssMmdTWzu8weEBWk1kCJK0E4Ux6uNKICFgoV2gTWY1HHXzB/U5RmRr90soJeb5//S0il6gqdFd
1N3QCsaPROk6sh3JnCp1ETmQKPe9f6/2i69wtOgHLl+y1Uy0w20UoS2yM+1bc+fCV93yn1NOX2y0
7p7JOeALr5W8CyyNQ1a74Mh8LfFLHwdKEVsP2NdkqCxzj72T52gWCqQ88vGCDDeSdw23eU261l19
eqEiEDz3zSLBnMZRRssmGGqwh12k4LYaQWoPDgwnyvdc2O1Rw1sVphdJxLHpKOxTflifVAbje94p
B2Wu1wCRubAHl5vRoL1My5Vky0u8C7tY4wgSGio2Qg+En+RtltXPjNJ4dFmy6FiUu6NumQmpW/wj
GBvQh2k6m/54QQmmpnNv1infkvrTkU/k85EZBn4rqpsyYq08A2OODmwov2zbYkOjTOJ65Pa/p9PT
UV2QcEHJ+FjEK+vkZHboWt24LTeoG4D7N0e4JMfGlJPiFG7ElHKeM7O0aNa58KdvIHimRLKLLq8M
DCj0ddye9rlml1DziZRUTPuFEa6+G9vRhgqoU17nV4NDk3WrUgvxRRhBeJN4CtV8KA0vpIgbAkdj
wzSCWp2s9Agqyex4s8guALtbflHVJp/6F17FBCfjdmCqqlTT9ftyujwGCNGrRjdkEWE/mxRkBrdh
4BbwBXuICVxK6BEA4G/ApBKaMosnVO9r/jgNymiwXGQC0+6sA70DQJA21yUflRO9xnkXKznUPgMh
RGrqG3S0HGq+RdyhyQPI4j/EpaRArplhhZDcvgaaF90p615/va/LwMCZHbcwYnUHuPSxgGOQT5M3
nZMYKE1ajhCpDnFCIrswoxaBwUGLZcG9iKTeTGvcFzEQojuO2bK6RPeDAGHBJPJfAggHf2pUY/1p
7O7yVb9ikI3wUU2vheItvqsz63PTobphbQGMD7dQO/8We1QIUYsChFSyCY+Fp4nnSsdBD9jo+fxY
iV9T2UYvh8FWfCR/019BobY5x6wtUWkaDPCW+Z0zH9e1qoQB4j14hpgcWumlSK6zzFpOUrsk6wNO
7xrVmbkNUlT+t1v6DPBxqo6t8VccEplvuLK4eMDVjcAyOnLNJeYJRChTtBftH9xX81bh2eTOZAOq
uuDdofQi0L14KVH3tKaK8/TcXEUPmHm4ik9FKpbHrA1wec+7AzCyDQcaCcF+ljMKePdOxDLf7qlQ
jgNTDEbBsgAG6u5fcmWLNsw/pB+Vy/sDv2zTM1WRnfHfOFSUbIBk7xDujIRs6S4Qfmc+YdaOfC+L
GKNd+LCKiLfOYmfmHBIcdZshB5xDiftujpcg6c8+ignk5KGFAQP+lEML67WevefPLiJcBcmBVPMD
Y9jgdAxWj7NwIPVvdt/0XyHnZDlAYyn2lscxHThqfCJfovgErjesD0rNTlWLyzQ1L5AL2al/c5NK
ONr0mG/q2bxD/+KOlnVtnOC/zhDKdkzdc/0FnYYUWf0JlOnTW1mXNY2+jeHBI+X7j8V6j5h3qP4/
jewTzf5w315REqjz7dWfhbB1YnJ9d/cyKpiobx6fBVU1HDpJMOEBYJQC9BdKgNoJEeU9UyaHakJ9
J/OddOjkllGBeh4AnewR2aDm+pHpefpFkQzyMJRwpitjJ8ZEqhroRb952MQ2Okm+szr5oJKHiOlW
HWo9r3nc54E8Zaq991U2Nis708Mq/utMZwaZikUI273Khe2a3Gtz8a/BMtxULUTSfoinxvEuX2MN
cCXpyIrVLObJ6CdIskcBOcppe/OEgKkXfHGTT2dDZ59H4zWw4IQgHIlKiMvskS5lcnmk78cnZrG8
8PtIIjLi9SweBiEwDsXDEoaOx9ZcQ3K8ok7JFIrcvcGhsfhXlvqRWGq4YCe00aWZ978jDj3Np+bU
qbNPFqAzsZKJre1ZoxMcg0jkybMof+ykFZqEHCNzECU2mBrd4Dr26uCLLX2/mkdWaWN6LuoZ93yY
B/5TN2b9AHYGyEYbLTynuZUNWHsPPBeNk6D5u10qobSZNg0DlLG8ijCl2yDxH5IVU0uh9rTMZrs5
JeOvQwcGIWA+59H0xmocBN8K47WEmRSmEZslRp8GvN1jMKluZtER6Y5sJNxRWWWmh5wSoGWEIFZ2
deAmwgqB4DZjy/+fKli9DTC2gSXGEPP2xCRnLkbyIvd6uNnn2QcraDEonhQwk1rCETwh/Oy2xMA6
/gq131UA1vhW7XKhT/Jwr6canQeu0TMMgN2MDNFLgi29r/YrOFK7L+eWfDnTKyJaDgQ1Dy2RICut
kvdGFEaIn/fPi6fAlEzP/NlYZv9TPcyPOhCNKSfEFSDct4kRKE1qlhRuIMJJoC3/hu6Zx66EhWX+
RApqTa/aXdpKei6y9S2pESdYIN1a9XMBjAax4R7eqwR1y+BbUilq8mxZwsHqgdS3psd+QjMo9TdI
4/k6ftOj2kOeQit4T6bdd2tjuBwvjQSrptJardprHxTkllocYNaWS1kt+NvlrbA12789frDdVnY1
MYxOshG1PdMkJy7CgOJFf6idcCkG36YuVNSCmoRKy4UENgCt5bygGEQOMjt71vOMhYbOnqaxLgaq
3x9VIsWTrELZU4bFERhVE++8N4+x8K8dxhkV3dAUNSZ3szxDyaiBPYySRHkrdmMl91xhooRGatDq
JAoZxA9tAo3YHE5DB7JFA7/JfzTsAipak6f7p8v3VZZMCa41YF4hvXNLtKpeAFAjtiNx/4wxoxZ9
f/bNcg7PwUn6Iw41C3DhJh+sj96US9rBzfK8Nx9Axm9RtbXcfkWQiDGN9lbexdDGYHhf1IRZcB59
oTbcGACl6F+gFCv/3JDIe8/pB8+GSb04pEcgCM7EBRAHaW/8fDGyo5q4/VY7Shf4bbtUJKNnrYaF
/aHi2hp9kmKe8Nbcemejrb7iH14XVvAakIJLBL8ykdL4ue4uBZBWA/Mo2/cDmkfPxFuAOiiP0D3L
0UZ8FaCBpS1hk62Oi24bbNa47BdcldyFAa7NpOVL47mD1UWU5pCWi6BBYIt2NonecvzlokEzy2fv
v9sFNb2yLQxNCqkxCXGaC/nMMYxtZQd77dJOYRW9OiGzu/J0dtTOTYFpQp24AVrYY1PbwxhQBCRR
hlCH7DdabwQv3AqYU2bvIHAM53qtpl0Lo+kvHYYcpkPDAmpcFA3Ik/5uZrrzq0T50FtzX/Y+mAQd
iI1abtE65BuvaIf598fbe50CsE2j+DFbNdty53Y3lI9OhY0tahI3FMZkQPl57rls9852+ONNcLLH
2qFpgSbVygHm0JfoPlf9tYbaJ53XQyoiX9msMn/vKP+qUTz36YccfDex0Inh52mfvkWGaNRvSeT/
BUkX6rL5+Ujkxq4N154mv5U2oGl5RCb0GwTABY/4cjZFkeLncfHCNl+wa4KrY1axkwolTBlnR4cQ
UpUJ9nWhCiPzxUyXxbdLhZgPxofueEJBTE60p6Afew8KhYt9ks8mtDxtBN7GCavHLV4P8yIMMBDf
jfLiKhzLtuT2DNknzvjxegZwh79re4wOOplCmuGDDv8y15x4xkX6w99pylaW/iYzQlFEhFr79/Ra
iTG3JKN6gtVx5H+h5QyD0ynxPGKe+Wpk8VxOuZuVgSDMk8u3dQnSJ22GO3zEGvpNpLdWYobqJOVI
18FbewiFZdR6TUwHEyH03l6zuopGiCyFSZPdOun90BHOgnhluAlIPSV+diOhoZBm/Nz3hYQ42MPw
mOaHJfUDVWI0OoR17Rxa+9dv8BBzC6eRCQdKelJCL7HzKnlRMrvD7ZIXkILg94M15A8A1+MGUfkR
rHPsOB9T+OogdNiXyN0nP5rB6m7YY1cDnFvmJjLQPL7oZxSd9GBFKFAKTN5vZN9qS0buSsZ1OetP
xE6RMJMfAeCSnNpxGVkd2h/lzLxoXYI2E6GdwjDdSoPFwX5nFsUxoy+BJ7WgoXsJlEr3F+uz6QCr
9x0i/5YDiiJ4oqNCLAIZH60VnzOxPZcT+pAw1jDU7xkJX4wxLM/F8V/7qe8PzzoH9brQFRjrMpRD
hy6eqkL9feSPD4trNXiIpZ76kP77d3SNCOS5NeuOTbdjhjw8Zq1mjVwtD1HHJcMd2R3Ba+3jEqAe
ZrT21PVGMGyUAz8+Qh+hgp9jCyjV0C+9GV4EOOQnBaQD/z+XqXMRuDZn2v21w4/Ra+bY208TdXyj
RFS7a7ssCxIq3OeTjU5p7ll6e+exADevpXseaBh3ju0zUf3zEq++kY/Y67nh0Ey/2Gru+s/+OX0P
XtU+aBfq943Pq2d3jrcbkIpjsqqL9XzobhGHEj/fKwkVS130m4Y08/jV4PdIMDSEU8yxVl7NShxB
hc9pb3w6DBWhpUXMKZJ9cs/yQzqAmtTlp3tfNMMxWOr4WkW+NTGTa31GkePS2YYm5RWuNuyPUUq8
Fu7tEEHxcAHUGMuvCacNbtxLDZmDgxFwFsgf7MmpGzPI+jWLEMEMvd1MsiHvD+pF+CS/iFynWFWw
suVDq8BuH8r847249Nez6ipEnAvVJQWB8HsTDYw1pNekuu85/QXfI6VQ8l0moSLcOcvJd6YkwvoY
1Q1Jiqwu2UnGZXtje0VUgAIR6Jeu1vlQN4lG591Yl+usrxKLyoIBNhbDPM+kcQj0bomrqNdX34aT
NUTuxUgC0uJ+8FpyD6QrIIwPxcQ47QK+ZfoN5iSrmRCb7oxxtIrHTMolkqGu9eZNdY0jc1bD7zPZ
kOcMW4dQAfOYdLk3JpbsmxuyEPWmffrJA4K8Cv4f45byKywfaF11+MWo3OL343sg2BRS4qT+InAu
MFXfF9HAMOtPczqozpCk+ZwlBtijNpnp4gvqdXV9jGyE5qmGpQzuYNjeyHh3qS5uCF0IrOHgz0aw
qHsFl8jFFmR4pMh76wAfOnGGntz9w3MW+fmJICJU6bXKSmtsWjRNzeLfWgwEdrzB9L9XIjVOOZgN
RvO7gH+5g4Ucsn5fFzJ+lnAxJJ1hrtAkuXiwLBTLxM+Z/Zd0CEO+2Z6JBghbHF5tRJ382z2GVRFE
euJk7MlMBo0j0oDHP0YU5aEGckXOwLbbLp/qUUu3QZ4NYK6jPlPUg5EYbnrDnnr1+TXRvhw0MQiH
Y4p5rPfQghicT6tJsfYj6RdzC7KqbzWzurQKvloXx/RYjZXUvfGTZr0MMt+at9AfE3JVrHfTxR5M
bjpUMiDInVBqdCsZJ/Z/hmNZbuDV6wcJ/TljO0XsoJFH7yO1+MRPFfM5E9LwsRkX653sdc5ErvW1
k/LQBKWnZjSeKSbBNolgMQRuSTKK1rBPgGF81dxvXlZf4fjWKfzVtXVpHFa7ZMJMQMv0dlO/j1OW
teyx1aokXoWp1aFlE6HVBwhYlQyYpX8v22GW+ugvE6uUZTBjKhWduQC6O44BADjXIPlU5/Rszt54
dn86oZzD+PenyT5EtwUBlD7idDbGAnJt7Mtj0Srwp79/DL8Equrz5ruOtYoo20rqM4614dyjl7yT
0dCA63SsftvOU+TIytaZaR5MxfXnHh+QunvjxirwsPLGLyHR8AQ8CUkz+aL1VXY4bvurLlkdccYc
0qacPxDSYbVzmqS2XLCX30DlsXnaxfa/BuQ/MiGlGS1ftVRx19Xq6Zi1zZV656uqw5cXJK1FgotU
o2wbsK4cAUiHb8+/aoX637XTuS7tsuFoJpJSfmKsv2kXYmVkzDc14tpkOyB+01z/4JkhnJ2ceivt
7o47IzaymSp/CQi5cexWvYJ3mabHHTzBNSLrDp7caeKxlpgQcAui7P3nYhdSGpl2TX8zyFsO5plT
veVTuUT4EEO11+4fWZnsqJUxdAz6zpGxjYeg/I+a6nM8cOBvuzRaEGl4QCv/Khfi4KRIL7QN+5p/
j1AGA1BI1qNK3cuVwPsRRKu5LSx1XOhxg1W8R4xo2WgPU1B+9JLUpIBaeBGMXDczvGizqGbzDnSH
o4iT/E3bdUoVUIrEokYCQs/NpZlbB6kfthnHVBfxSqFTusVPxEG1ko3LXGiwWggIIeSzQY3seC85
IhjBqc1UsMFSB+A1zD2rKPiXVtYaHbc9Z7gM99kEje5AatUOVJLjPVI72Dx5aKhf40P5nga8EgGJ
5H8uZOgtcdtYXBAe4uNqqB9ke+vF0fOczE5Jefc0XKkyIGOowtTuccYCPquiFvqqOC9bBQ8pSiCB
9FLDmszjOAYZeWqrGXCWFwyT0gkNAVueA6yfPFAXUAagLYND97G1n8cLqYcDI2I9o6jX4BHizdvT
rV7YH1cEyoNMl88WL7v56R8EZ7dLEw4iSaDrhILXGVqa3OxvAcc1UrIpm6LxcNbeAzzCKJyehIbN
RP4Vuz9ZXexrZKt4JnBmbCjtPGskqmx21UFZ08r6G0jNaAXn/0ZJJHqRa3OpLmCB8gJHBM8LRNTg
AUrIk/Eo3mFotnsUDPUHQO5FLsx7AxXJ1sNJHMIFQ8HdBfay8lUwTKtQEaMFX7VsYus2/RL8YliG
KncM2V+6iCrmvB6BcRFPxRd2DakFi/Acb57x/eBsanyP3bT32kssu1fg/EDQFqGxyX1cZ1erkMEW
+wbZTxI1hwdR/0WBB+E/Nt7QnJ672STCylpnjLn11lX4xuFVmxdPU3kzRXVYFf8jL+hVRdo0pqSE
d58Mbrzal1Z5W7YaKh8Y9/N1NfcDzkbunWeFnubgrF5M8lNG96s+wKpEaCRYPlfnfmq7qfFqf79m
X7con1GDtAWmypxHqpp8LJ4UUIsOO94ru4l4lLj0x/GwiP89X59MBYhiYhkVSjjJcET0OJ2nf5SC
idF+D9VlnCKqS9Eb22a0Pm8XXJHK+RNHJ8mdRMIAnvwTFgaBD0jK+u9kQZRmsbPBKxswmfRcALLt
vVWk32SqQMRufIgRaixXLpQtWEnJ6s32hLxnrbz4xg2CDvp7oY3J4hvqjEnwQ9htn6KRENDTQE1h
QwfuUvs9FMx5uaqR/IkQa9PqqBxDHCoy63fFkb/9HZo+Xrn4hv/xkmxh5i8goU44ezYkhmlUGQ8G
FBdzlV5Cx8xRhibUhUo2uWDy/ZOMsHRoeTbzQZm6AaL+Mnn+UpdA6qtCXWEDejqsKY0M3t3EwEWx
nB7npMtS/p0NJso9rJ2dIaWdOUTrk7cJWT5BvU2yKTCSScXZN5aEwJlQ2LdJ/U6ak52zFmIqPvxA
MTdn8m1DQj406fYmd2gPY6tQwZbIgH4R2hCUEIse/RlGwGws5vFzIaLMZ1VnFVPQcnlav9lpPSeJ
4XVWxOmWs5YlSDXT6XOTpITwv+3/bo6jPUNdvWU/pAL3vVR6DLRKPvTOV+lHCH+dE6qIt+OC10si
Qp/H1cymcyuj+nZhG/na7VR4bVaCrIyYAsdYVSNzRct97ExiZ8mBrvTA+sAOV53ic6F7FItv2n7P
6WQyGO4y7No9Ta0M0cR1ayQmHMPVR8WrPs5aJVUr1StDV83kpaDuOGZ+8M2w6PzHE7w2rHDnjTTs
hsJx3y2J6A5OckdFnYduj186m6vndOcN8VWoXA4G8/SLKQNM36h5NMVmHIl5WylNSB0/dXDB/2u7
3kK3oGUQAtfVFCBZKgyOWuNm/JaExsQiRLrPb4h/0GNmuLsUrTl66iGQFt3ip2tb8Nq4cgZnAB4G
1OGCe0W9r/6FY73DyAqQhUCmuwOSedu7PvHdzom2NWRUn8A2GHqOR9933MSYLUkVblq1LK31WbRh
CiGPo0xERuJ2Ie1QSxFO0Ma0eiMhbgiOYGJiNAnmbrgNx5X3d3ZMlzBFSRN4ePfpl5Gh9d6rV4Xx
jYF5eqgtOkGuNJx129wNB+yEzXnQe92NCvVqCwldaZrLRnNa4mT7I8XjSVbCBbuUPtDxngn19SDz
VpvekMmlz6LFvIA2BBFLjslbPYzvAGTFMzxvETtCJ9nmBSunOtzL1vnUD2XKF9CAUBcMyCsAph6m
GAw9lxcoMzZZnOYbZzS1oOMMGmG0CFPtSc6N1HYh7jFtJQ2EtYEMmxMyaFzEQM2CAhWQItStMNCY
TtLQ8XeBHwGxxh1rFcci8bjjY0f2lLKt6uv0748va/1oLFLYgGZR6wVo21qmqF7rd9lKgGPB7+O8
QbruYNofIaLFcnwaeeWCJYWKt/PhBd2N9/xHMVs/1qK/IGpYjWkCRaUFNDxEQU9+K0FaYdYwBw38
6ucZcoYlE+AF3P6IdE9eVUHu+yKSrOY1YJFX+55A1kASbFFBZ6fRUmJpBf9g/QC9zbEdO8bGmQlI
U6zmFIgwVn22bhSy1hXGqAV0DKSlYKzuOMp/rjKef2Ujbrnp3riPXdPeutAv69kqX6oHZ1+vmDBV
hsI1Ykaq515A/EKKJLhyeufT/m2P7GjD6SMtpxHLmXzDVQp1tIXxGzzrX1sPiGgELjbkWzioDZO3
orKUheb1HEmjlztUetPXIHr0oGk4RHzcVnu0PlZ/8S1Ts4DV1EG81E18UWO9f5qK9v50ZV3/8sFt
/VDOVra5qYxLN9S2ow3iIs7IdeFI4WSmEVdZymYAHUSz9vW2qMV/kTnzsmqx3oe2R67r8bXKoHBE
hTrvxGMLWrMt19PFZ0cBQVjTQqxKED3w+ZoDiMGF8yA+X4lXCdgzgtBcnmXKwmqFTHn6elB8i/td
/YaAQ9rWGgMkY8EW5+aXsCUAjtu41CJXJAkhkfvPLpF54811kY8JcXjzZF9HOMULazhYcEAcX0Ef
ht5t9Yh0wLdcu4dw+q6CGZqUoAeiB5+wyRClmqOJNBqAFPBTVTwfw2tUwjKrbCga+CX7I7seLSEL
INkWDK54g5OLnD0muRfqQsSLwday1fR/5du4A4If+SFFlFm46uu+ZmHwClMbX0boV0K5v2EKasi2
aVkcvsEv4bDsFlrJpflrvfsEvI5ig1zUW2YcIDPpC5ROS18y4+WsERbCdNiA7JxjUPsO1B5uasmq
yC+8gIrb+YhULsf2eUIyYpUuV5Nbv9Ir0Eu/7upStjC5pX39inoXTn/zoNrOLC15c9llmb2yVCh6
ScEFBHuFy1Mav5mnxTXR8/KxZ/xnKzO6LA0cROlRVrHbS6WDVndabGwFPqCC8EVrrM4W9/ZYyFqp
loNsEb9F5mJvPVp0zBGKiqSdpG8iMnmJ/4tqaIjEGTdSw4dIoDkJclEsieb2/L8kzr3rLIUW/vlQ
R214l2fpDU8pjuRsL2+uyHDUbsXvfIOj9Vl5TS9mfaxitlJuXeevx2SqNFtjDgJyRbH65fTl8YN5
rVz8UZOXAsm1DY0Rrf4ipmp8J9LThB1dSKRvXi813ioIUW0yn92ztbk2TETGhD6SEgicyigaJRav
DAekK1moeJReNbCRUGZZD9Et6WsK2at0U7YqYOpsQQzDFpMxQOQ3qqAHhFo1peTWCzThkDcLZe0c
XbNjda+3BMyJZ6tMI7FnW7mK/eTMjS3Fp+FoLmEsKMl3CJ0mxdNSA65c/FeG1UUJyaRG7On/HZQf
AHm211LBKwzZIlMGxGjIyqS2kgeYhQd4OU5JnurdBak5mp0SCRyqzUjQ34y39GfUX8HZIoMEhGH7
QkA1bK72fQEBfdjn8rfGLQIp2ub9sItPFhg77bRVQG1aech5I5odo9w9UNo0JR+95/DPbetGBBKG
1AlrpeJ52cPXCj5phIAq3M4hU806fn+VxeFN2vC2rmjqpPdTAJcnNGqAChRssTuDPVMwtQJcRSlZ
adNT9+wW06Ea5trSCwq46IeqnBuZImX5Ixs+UOdGrjHe4dohxYS4BSxFXNu04FYOJzBcqMf9WynZ
rZmeTgjmD8NxAfCIQkDrnwP01s3Cjex6CvRJukdwA68Q9iHIl7td5yL0h3lVLcj8h9cPTTzBMC5V
H478meKjvp+tbHmnwBX+KgQmGjllVpF8GY/ZQZWORsSft5zO0F745NzPsL+EyqrSbTI0LLHtl9nN
T4y1oxM4tsW98Ok5fgOedw2ITZCRqhAbgdZhOn4+QqnGKC36+X334ziUVT1M7h7C9HsrxVAHkw+5
dJmjCzxMnofzwrDWVMgbh6mT5vlFbYUlgaJ9j+wW4rtJQHdd2T4sU1jY5yq3Ev1UOJUo2pZLwyb6
UX0G3cMpOHhmk8JybfWR44onji0Lnn30iwTkXXOsJCT0UjC6wJFH00k3FElFGVjp06nkrWaF9PPh
1hHdltS8IGkQ9QAkjXXOXUYYuq2L3qksLVU1m0uKbXl/Lq19OYS//ZZBlVIlWQinAX5DiVINknMF
E08M4OE9lPsUumnlvVNXphQUCGAtdeVlybbJtUyVU/L5detvZuA9h4o0eRkCsGOIWgA3Xxp2CYK9
iHMy2n5hOJVSoFvTo49JdUAMyNqhGuBFbJe0ntICc7skfoAClcZ8uIStAv1beZH8r8T3kkQHlrWw
rToz2JPNizQJ5NsnGvvjOCMUtE0ojB0fx/g3fKsbJMsmWXVNblUrXrM9Fiik20u5Y4vS6G5Wfh/t
wLxtTmZjoAF1dul/fuiEghn/DeUkJQ4CpZ9t2FBZ42JmdeqPjg3z3ewV7nJl/qNE9TzHmVPl88+p
Mt0EjqGt2cWzgGMD0Bcbn177Ojou6fWADZ0guZ+hwEfYWvlszh61sgtDlAxrzXm1Q5Z6TVmtNzss
sNL7+eVdyt4mfvzvfFa4xUj6Ghwh2cTnblzadDJZIBdj4MyBxx195uVgO1D88ttHQshaVHpCAdd8
ofERZMvyznbgUY0Q55pwu2k6ILiyY5AId5a/wUbO0FyIIzZA+Yx60VMOO/F7umtIJUGfuoWGGtHJ
hXFJQBnt64Tuj+l7buT6ynD9ffXghvdnL25Eif8Yv8teEqqG5THuP93moCm35jrKGnXKkwn+YvHH
ksQ5nsZr133GGvphNs2CfMIg5TQpa1+YmpKJGB1IjcT9rV6p275mmLgAeYfaDrA0oTlZsnJqcgay
jSOqA6iZODkIUFw+oIs3Kp2n2aeIyJV1gB+fOnDoDxNtJ3kFp7h0iRLQGmJxSozVr7ueWDflLO84
dOmLCSadpTIJNZ8rrSe7Bo5525MqKbLX+QjUWdSYZIkAqSCNCvBK+s8dGDEcbiTClfDGonAZI3j2
bHPS0EWnAUPCrXcoVwyR6RiwUo5yiVdfck1KvUNeruWlVhsoTHrlaTCFKlJp5bZkeUHxVIdTwyvJ
dOuKxbKhj+0g1FVlnEqvO2Khy/HvW3jplw2tznf2900Bv8NxBlhM53PQx+cCTNECVwq70IdGyfVf
/4QosB5dSPx5t7/YvDhdHEHq8THpJs1z4ml09MOQvuIzJ+YT5P8LIhk2Q6QoZpRnyTxO4+CVPJwR
0Fe6h99/gGB/LlwELoRn56Po+OLp/mCXJubdd0X0wgw8+Yjf5+ExINlsJLdJHuivvMJU37hZUySr
20Wk6kWU2LZrGJjs+v4A96evrI1E/HWHOG7Q54dieCdQe3jhabGgPX4Tp4QWbjdtdlRrxi4/C8DP
5pogINfn06TWJZLdg4ynXuX4Y84hD43OGIDVSaMUJ1FGN+ma46HQLukGG20b0oSTqdyF8Mi34Upn
UMgUVIdOAV0DZKeaNonrZ9UvZGOEZD59SFZJrXiKRALToGG/pUd7F05Y0HucytUigcdrvAGEcAO0
NYVvdUmlY0+vNtjmDe8iXov0Aye2b2+lsj+hQQy3Q50SKV2nMf18woDKE0O9KYsF8mubz5rT8/CT
KBb2Uf5Nt8tnpXVB5em6SLAcf/Tr07AJ/fyDOZJCvD8ITvk1s8erjv7pNSMDGx3zwbSuaijjxSMk
0M4Gs7gkS+Xr+5EupbXnXUUIsE9+45n3kRlFQeYJRQG96lZGUS6YqGnIXRKowo+UxRfGIy/gN5ua
ToUcIwkw7xNfs4x5qMuLU5dPDSOVQ/Z1l5Fh3yZ0lNqIGqf7aFDxtN1L+ltV5lAg9pQWeQuoP/F2
B/8GA+EWwTepSVdN6DziOaAVuBSFW6alWOVuvRVZrtKXTLnUA8clXQHqb52bR3hSY6Jn8rgJ7GXd
FGbUB9cv4wCyDlCop54v7sHHJH1Pb38odz96juW7QOibM2OwK+BPxgA+23Vr77K3LBX3AfGmMQPI
2ZFEaAJ1YgJskbUqs/yDldG9oRic9jk9Da2oytsCkicmh7LSAAqizRliCgXr6IMl1fmuuiMiXQn0
lLk8/fJa0Vks83++wdLi5nwoStxU8NmV0U8yKN/kWkkTObloQY3JtXT0TzcFO8qRDQ3FYCTzgKst
huKNYo2TEUjX0HjvaycIZdm9AuvJY6LcUfyre1TxFcOCJsA0U5Y8fNHqMNv7rsGqM0VPuEeZU9h4
DDJ0MNUij7tYpGPCam4Y87M5VgqCPIQQzeRimrmgabcGqP/IBsjiXkyI5mhe4/g224p4u60rqHQd
8uzoHxkOrTH852D1bwm66oACduJ/JncnYbB/4o9tHivDOjU/rmOAtcU+LY59wiOz0JvhMFYsu0tc
2BgyhKaR/ndQfVsXO+QEXVMoF2u3/cOfA2SWDrzW4WTZbhmC/mzYjHLXViZldjd+QBlSCwNXdK0B
CPRNWVPY6R28x19iZkOjcTX9OaqSDpHKX9/gnbIxpb6mTm0/BlliR8IyN9+xoh7+SS9hL7fXcuEU
czzoUg1ENqyf8cfrDgxpMhtbpnin7cebe4Wr+8+AbeBev71pjR/2RU9bb2wsf6hXnHcDpXNAvm6a
Dk57muIuhUaWlNJa/qiQQWUCg3piLJLLhUeP4TVWfJ+/msb89TK3iKpELNqgYWkdAAV1oXY968Gz
hxXAFwVMoaES6kaSFyv8tKpR6TG3i/O12fqnMAm6O9+fUBXmDkm/SVZsbO+BNFoMC53N67u5Oof7
bIIY39YIMhZZFV8eifHPeYwbgIe7dfmcyUJE7Z6ooP6MdnnEsc5wKhObTdMNQu/8ApFw2JAuhFk1
pi3qs9d+zdOVoEaAXkNKo/lLPt12sQDsE8qbDqrHGwgd/rnRwCSC/ouNFKtrGJWYsDUdFoig8uXq
c+Il5x/2OZ1PdwX45pJvJpRLopnEgPqZgP0531/Xl+OqDPOrDv0FntihYQwsAQIlMNyL7JUlFRKK
axZgFF0s5p1xTQgA4TXO4d3AQbYGXUfIO7U0xlrSl0XLBPZQd4gMlcVAQqLRVERlYTVvNd18CMSS
hJK2HHpuPC7KLqwcxQs/KUqN4ZZllY7A1buLkf5zCJWYvrJQBH0Sz15Fe+SFd2i/ECVREsGfAJiL
h5xuKci2mWNnne55HM3H0CntQ7/xuHb36IwGRHuyfNv1hFZ5EBv5uwEdwbLfLMmkPnBSJaDADjGN
RPSusj1pSnQK4jKriRedIM4Hn4qdGq26OEddlBUA7MO7Exl2VBHDehNJzH5s58GmwrIjPJAZnRls
olCcHB48pB/WlP/co7korXHOw2T4HhRHHbutLV8nQ88/psEWkGjk73fbQ5MdeonpOm/ZbkzBkZJu
6J3F20IPEI+lpQCWBLumord+lDoNNMVggseWj+UARXhJ32aGEoL+1bIdNgoGRmXvtCC812RoVFGJ
VUWzV/uAvC80j2lj90k/KjDbviH7MpS5icfJ09GWHeH+aTvVnj3Yd0VDMd2NKsSFL8fJFEhLXivw
i3/VNNOp2oWvU4jyv5hq7p3lbJYS5yXZoY8BDCvRB9qdXRTHnDcjfyxNZxUwHVShZAl5xclpk7Xp
XJFWpPtXJzVKYNAviV6ir5ZIpFoMetYd4vT49V3MEijnOn5i6kiHI/S16/LAMaykJrnESma/LzjT
TWe6PnPYVs08KPpofcrGLDW3MmBwkVJi+UVTNYZ8Epn+IfHTNMsC7W6Y42wD0N5utoEm9ehfEU0O
xxScYbNuFJZu6dRaUKzxgjzuiO2OxO6vUI8HUFgRsDJpHdnLQoXuKDxD8qvrZI2Sbx85tVSfUH1V
++lXv82+MN9qMDnbTsxMq55oCmR6Tm37NTe7AhjfDYSFdFtFfN9OTX7zfbJgyHr2BC6mmOdjSNwr
1tmK9eL27HkHyxuzvYexh3cTFuCSk5k+7UX4EBG/E/txL96Ck16Efl7j7P46k3IgpIRwypWdbOJ2
GMve3VrLcz4NcqseKBuiZXrensYHkHkItqNJI/ph6HYW3tffZLZOjtRu2RF1mOf6rgzDsUaAfABD
fvOHcWdny5LncaqAI0Njv+pbVYmWeYVBiU/Oq2ImLMjQ7f80cciPJGW3aYkkbR8++tYKwgQCsbuN
W//EWj9NcSdjt6ZeSWwEDJ4rWIrn+YRUb2tNbBbT9C1UZ2my011hBcCwT+Y3qSZBIQBU8WVbSkzX
WaRIgNa1W/PI/0ls2R8DNDVC3GJDQQgirW/mNd1vuGC0fqpzL/dMN99zrAFQlfQfSvWA3y8ZQvNT
wjoNCKBb9coPY2aJ9/pD7eQ/t+vTyLgKliHcNvx6lT8pFXspbh7GP090xIiqs/hxV4QLKxuK7XDz
fLuK7km+UOf4CGi3TAS43FO2x5tMl6zS3fUSQ25BFpEijCxZHi1axs5rLysXbotgFdJ0Q5gDPwJ6
tXGDwYkl8lyyULED2HiBRGs9srb2despOvUWLrjLZ/k/pQarQhS5WgIW+uP41JeLXWjbao103NJp
4QWVZZCkFxmQQfzkPwPG6z7pMiJK52kMZLpc2u+NrqAzA68kMRw4oSg1yggCvtxD1qqhjURyC1kb
Bb2LdOch658ffxwg+sTYcc1qwM0OR4rCt+Z89XLWZMO8pjTgySMU2If7OVZiJAFxn+4k9mYNCVoq
3bKjzM5o6fzw03B4tvzC4tihNa5juLiGnW4UQB0u1JCAp3+ZQsC32TobxJGXVJj3JSumUdg/rIDg
6aR7BzyJyEhhtyMhY9egOodfEAhE/GcXbjjNJ6E+lzmsGlDKhM2aDd6KeOa3q3F8hpeIEPWfBEd3
urB6ecfVzfk2xCzqX/xgtysp3mVDbsZjpznMXUzK6Zxx4c35kiIXSzD0w08/rJjAGffBU0vdiPNB
oA0F8+5IZZ9UUMy9+VIKzSk57iHpvw270n3zhF3m8S6fdBATqmDYF7JJie21otodgyfQQ+8b4SzW
B82d1fJAm64U5GKOdBlzHLuAJrMxb8LOIx6uh3J5vyUbN0OfAalv6r8x3g5SI5g7u8H3kP9asqbp
QCiuNhNhTpOUzS+o0mBfo3Kskmct0xbqTBN6StzXSXbHUZHqb/x6FeWS4hyJDNtCMXCPjAA/bC82
ZrosxI3WXqF7i3FAYprgEIlL8v4P/KBcB9Kov2eoxoCmWGleKYnucJFIgIn/x1ms9+sawrvlSgWH
oNT8Qf7oVS1f1t2l0hkQkGgJ6X5uRC1lC8K8OspyE+U3S3rmzwdKX2PWhD29a/qW44P+wdBUWTaZ
mH5blilR2HFI98zf5nzZzJJgfVbHwwu/zKM4QS8b2LaXGzCyURCda9TarlIjqbN4gDjCg2vYyAtm
h9PEaHBFFpDMO6DML6QZsZiquPdiAPxLkpsFVNsU7BV1OE/XmVcMSOcIbQ4FAG2Hk0brOgzgBIhP
k+ynVD/H7SXX0vDquDVPI4S2Q7ZMmvwNdve5wjaR43+r6iMV1UWzSAthMbEL6lOOU3mK/Qo5TByZ
LNiUS38gbz1aNzF5y/au4lP7u+4RgVZrMLnVw62gBKbgqPkIc93r7VpYxulfMIg0eTzWi5lW7djz
W5sE7rpYFXySjO2tC1pM3nNdtQd47gECjaj5cyl3bT8rFc07YxEI/3RMoq6TKD0rtKP5aC8U3Pp0
FRhEQqkasG34qNDH3Sbfz3HLa/h+um2lpXLLUeaJWb4fKm3i/tWKbb/91CAK7yFGw5DyjSp+wDuy
52HIfUhQkO73vZQdBJcSHzF+XwYRc1sOAQk6jJVBCC47FpnMlO5zjvPz9hJIp6hfxAghNml/fWNC
yrk4euwKF6FPvr1yxuF3cDnZ2WezqgIRGFbayYZcLkRI+cjbhmXe6gSHbEZyZCA68u9+rLSk0SjJ
OsifVzKCNJoCUEoUcbjhz6wRWj1hkL8IdXA/j8ftYKvcxS3IuWTNz8AGYFKxwXYJpn9iPGU0/5w4
oihMwsJOj0CmnrRMWIFoILSG6sW61CQTXYMFueZz5qldhPOlfcqmJAS4RmbaO2i+XDZexHNxcMo4
mM/obDp07rSaeCUxLl4XH8EVLoVgrS+lgB1tFsPqgnmwet9pguPno2ObI7BAUyP1AZLOJhUDPQFQ
A75H843xnHTPwqKGxIaLb8T3JN4DklfePnD9IbXSE21uwQGXg0pacFOTWyNYyHFRq31G1TAerOBC
+5l3Y6D6eBNIY8c9/VU55FPI7aXsSSA6wLPokS+1PVlGJiWTqa7Oc079ZEkZZiVpSP61GUDnUj9Q
w7XllFbivBFfM3YnkbS0NaTIMX9yec1zKMaewGa0pBFGhCCT+ca4U9GA2MIcTfYN9Un5DGjc2/Ab
GnMrXS4ivU7D3kGQZm4CBxfD37aFkOxJj0NO2mhbLfJNIqz+RRYsca5fpCkq+f3Gys2iAlZzUDr+
ay5Fwa4Zauv8BVAk4G+nTgCSX3qqRptmoyf4G5rMT/Kukt47NeYWRIBaczQwMHCvC2TquWT0/kD0
D9zlopK+xOPaT7KWOluGY6m7ahVHmFBPwNbvvIV13qivK0qzEnkDbyxWRU+kZbMmFE7IpzAzY7o6
W2jd8swW/JDdGBYQk3qUgg08pIsgMBfn4QrKvuqvhqht0Siqhb65Kv2FaQTJWQ6ve5ynEZRvUQi9
92ek6I9/pTQ+OqLaZIltMqyS7XKj2pzwTfTIyQllqCGVnp6huv/lrUIYtDp/fhXkQT6XwHF2sXAn
UUcqE+8PbSiICuXYp4fCh+GGCJQtY9lqUXccq/13lijGpm7lle6wW50RHuVnoFHUD+/kDITsC8T5
MOc3CAF/P5smdDmS1Y4fdiCwzQ6KuEJTx0a4sKW+WL69uUr76K/gOYzX7rj6lKvvWYCtoY30Ph7A
KdPA4iF9ME9Pb0feFm//yt81TgRexMu8ORUmCRLMRHWCncytX4Onwql63f4l5dw/rgasCFGYpvfI
0yo4YrG7gPpfwSkrhGXC23PKBfod9cgRr3byfagGZDYoYX57FFGtZxpxhHyxYMSfxFmt6A83daVz
YtAm5bJgOluLfXTb1jlABYa/QVY81lJTbzOQCzlhjoRPu76oTPiXh2InAbnBhS+F9cHVFYlsr6wV
8R2cRHOsBRnL7+o9D7BpTJ2YNXpHUaFXLQdL9r7UxKOi0k0y3CV1MOAX1HgAV3CCRNIE/Kqee7T4
LbQMvNEbeLQuhbp3qfEK8xVmzwxk59ZdC/HXdkYosMjMinUYoePDLAbM4775YuBpH2DMUT7IFA8Q
TwUuONNwnMYcpfFK/wEQohaRHF/MxDYLHwJlAitZ9IvQE1yKoZDAwiE+OxMbwEaSwgF0Z7RSs0oB
44rQWKB+3hlB9Pc8gJE27r4GvbRRCaBJlG0lDN6F3KsyDxrcjziAxReR2JRoFhgKqB0jIW13PbuD
nsFZshGQlW7YvCgYv3B7lhLHPbWNok42fw666n0yQ0F4u1qTa7OdIgAuYyFkq3Nf2wIBHpRNVAMn
Shrt/LYPPJMuM1R4DP135Kjlk94keShvHND5bkXEQ7mWbi7AAaNh5qTZ0HQY7Kch1NC7hbnkQpqC
MzEFP4LnELHxP27ciVrqZHoG4qP9N6tphZHxYMhBjzthRxD6n+QWMvdU9u7yhsuXboo+IfcyHJFd
Vtnds51QFPPeC+n+RiB+6XeMit5pBGxI1IxWpU1CD+5FnMsqVSeFKbmiCGRdwwZMWtLZtdvUY4BU
beQwbGST1PfiFQHbGc7XZXwDGA7D4VFZyqH8uaL9tgfWdaKeRi407BBeH92FyWLJHUuk1QiMc7iX
evPjtpjwCRZe1kUmjr1A9/sEktamio/R95HxpBtjAvykyS7mYGCwzhgkPjs3rMo0CQJ0Fp2HF/9D
EDTF4/do/qiY9aPEhlWVvu/dDzyexzcJYz2u/7760Z08yuViTvGUL6XPjGrBShjxWeif+61TOuF/
V3HoPhQ5m7hDqmRPT0n0iqMZ7+F/IrFU4tVEIFhdg/RICrrjpSgWJpOj8ql2kdh5anbnt7vwrqbL
FzEPYg5nGeOJyyk7uUdFM4xdF/pjDBVc2dGSPfPQ48EPchFvhnbcFmEQevfB1Gnjqu4/EJakt+yC
geNiZz4L5CwIFBBksD5xCtRHSj72KIvm5ztXY7N28lnLvmmyzNgVibXlNbz9V/+Rbmm6cHr2W7Yr
JKXq/NeqnwhWOdeE0+u+CFzH299xeOtsA5OIazEnx5EuQ3LdGc++aA5HSxBBv7GhFrZkwVmmgbvR
9EsfZAyCHk1QeYe1VPW+meILTXVQjYICV1tUE9VFIBQBACQ2hGyJ8EoMY9aAf8Bgvulg+bOhXE9p
FN19TdwA3De+CxFTjOLF73EF7UhiKd/sal6OcTLDo7tvCf3WAYymjRdQfpuu9/5gKGCdI3zoIFo/
PHcvyA0CK98wc6jJnpRBfvHNv3iSKhgHbImQlagwfU2qESiQtDGmuFWsFhAV5m/xsR2HjQ6e9wrk
DYf/4ryI5LmKCZKKnq6cw1J2zug7IHenX/TDemFdYMFoYIsy9TSm2tozZAER4g2vaPA4e1xrKOkP
6RFP8Iw9jIl4+zDO7AgIz7xYyIuCAfIHVrEh5K5umqkphpOn4iHjMz/b97waSPABWKiTVXQkJ4Hd
v8lnkLHbI1Le2qdbZRGH2hiwtsbNRsfIj5ysdqR+lnnM6ZFPzMOWzNDADw5Mcx93ugG2SkD1CpUV
BUMJdaJlxRTbZ7jXjQMepWo2juXxKTtaqHST+H0vref5/9pWi2lnWE9/oNt0HCKtmV3/FX/G4SfU
q3ay3TaFwR12TRqBgn0YBFQhfqF+rvJvD3/JX5irAa8+tiRp/ZY8Np/tJPXonRViNijtCttvlnxI
1IpJs92AP8YL0ho70wLfiNxP/myKMy/ZwN5lE5z6QoVkDe2PqY9pLD47zE0iAgmjr/7H3wWOVTIW
YzSmTajaZFchOQHU3wduIHo1w8dB4LmaVRYCIiB4Dxt0h4qRRAhNE9vEsqZPcmKVSG6lXZMMzc91
yZy1OVv+n23u/D6xkMGCaq70KeC4KV//1kJarM5D2q/8lMvLCUq52R9N+UlRASnRLeT2ZykedTVd
jXnd7xSB7as3drD+zrrvpmccuu7jfYEnnQfJbBYU4/H62VjH4zWC1ZM+IIwR8lDnd9FLYHEq9Hq4
kFJsRdqMQ+BW/otqgA/hpWz9M4mlZBfBLYVXWhcxDBIgUO3VbYi0JaYVP3YN7HuMZIyEDp96HpUG
LSKPcuUQ9Vs13ACrHpQTR2WrNIJW2w3siTfVnM7wvJhfRWc1d5QJcfkQDLh85B4ibPsBdZm2i2yH
n4MDWWC5GWgh2gWy6gPhNTKQrKp5sN9GEYMIBbU/nveD9uDa1ZDOywoj7WQWadrEzQISJGmlLTnr
TF/Sj3pDzlj/gRRMETXZO2yGQVV3ZLPksEqP/jBUA5NhdzS1A3kbDnrNdvyCxQps8M5XZC7EU3Hz
uJNoalmAXNeeZlk0v4CCqnCMfAdSrZOS0MzgEF017MyHjkB7zLONFMJ6RGfZ7Qy8lfBzg1bjfNoL
YqZcewkYDqwQyKA6uNiWmsCPNb1LbMizI+RqntB+685ksF8ADGVp5htGozLc7I9tqxWpB40wX8d6
m1+j/3o+c6uNu+rdFkPgVUT2tTkMyjdq0u69MAGTLeU+0hv3pxB9P4Z3pqRM5tnG585YbQTvWkOo
6Wyv5w2MDhTPCJ+LnZOj5Mf9VSgXdZpWeq1MdF5aLpY8em4aCXRzizc//fkxUdPSd19XxOhH4GEA
I45g9yS5P4FXwJs7OucB2cg1cS2y85pU2GjxUiRCzDE31pwqaL9ZyHAvDO+fr1Ptmfv9EvHxtyDW
6zgkzuMqGjNz62WhGj2miP5whwz7bZXir8kcmCF20SfPDXj/3149YsXG6hN0KwOK/6uTxeDlrstM
QulFx+MGhy/UQZmcnHg7Ws0AxLUmrmbxTtcBFMdfh33KqN663/VIcgKMhqODWrjNbTmP2CWM66mJ
Zc7iF10EVgG3Qpo8PDqyR3NJfbsueA7U2M/Q1CihbYV3KTgC8Z7pZCwfyc4Z8wDNto6IeisgUg2b
4LmZKogXIe8InXHt2tKj8OX92c776Zi1m0d8d2v84ZS7Zh5vxDKZd9fWGcRKmsDTKhhhPd8lmYJr
34iTtvuOwsy2/lAasQ/Np744qriuUKeZaJtO72ivUAOSCYOgiHrp7NP4m5OngpglMXTzETCJB2Ht
f6DiE5nDoYC5lMXzchJ+iGmU7+fcG6nof4kk+G8zklMdKkHa6pgd1hEbxjkhgD+QNDBctdNclPZj
MoDQg9hAE0QNptc+wuoqSoYLuBiurSsa/m9waEUGratwXdFO+jwZOLno8+MgVSrIjG+C1B5rhrJP
EsSJ92md8El+AgGzgCidmGWIROnKJM25sSKN95QebClB8n1e3AaJwRDueE7breqox28gndnp0khs
kxBAunEaWxGMJ3uJ+ja2pzmAmGSe03ax4KxGLEquZOMkRmtIwYsBhdPpm1iTCAXrQpEjvnNoxj8W
QR0u+Runw9BxWmwAdH3RvjGghfEMEH7aGtjnFjuHcEXmjmYhHYuIevKL230gOyQj7CBAbesMwXbs
T/V8cOlCaCqHTAZ1guV2lDIhsgKEhgnTOT7dTLHDiKSKPqoPIPCah5HdyT1g4PPYYuCy4IoUUQtJ
pV+Hrs5C/80rbnsgtFotAA6bimJakX7yOoXP5qNKpm17RFStYBo0e7uFEbl7zvt1qXUCIaqzc90G
jNeAzV0y4dkZ2uQSNRy2o23vFYSVfFODUlEk+lmszg7ZF4ILFOENTas5W8BKB6ffkuNXMt18qb8/
g8FdvjSSqCsG8K0lbLW0/8AkRSOne9IVC4XuwYRmrESdYwUvLQ4pS0HPa1FZXL6Ot2RtbeN1wuh7
83t1h0Ie3S3RRpeaFBWFGElJ7WC9NZVQuGwlPctxZcxZm4NOfl7Uzzbh8UiQnYdNsLgis/u67To1
s7cLPPRfN2N6BPH588Ahi7ObcDUDSRBPNhf/2flWJi43occzl57V+U8XZ2aBbCZJ4uX81voFKefE
o/8siexI4Mr26cidsrE4G8058dgaJshERZF35EQJ6MIlEXy7yN/CK2rNDp06ii/psX0PxNHi1T4e
D/qSH4dzRv1Z0Ey+veZIIgFOBIUhs0rVyEypiYbf4CsHNtYZ/FavmTf6NLW4GqCNCeyPj02f1F0B
cdnMbSamMX+BgpmRutVYRinux6iigcCLwATmj03EogoUiSj/adAjv28e81pbfi5jUwkxBagv0978
mxz56nyaaafhSW+IVQ/VtYbMcRyiBzWHxvHYrUntb7T+EBmzlWp6rFJ7xmOC/5j8QNoizR+EyQe/
WFdeAw9/mpoFfAXL9Xl2Gg9AHy+jvL/afgYjK+5IKwQDky1E3GEISqogKkGsXEyE9W9i73aL3dnt
epne0n2gpNex7zLgKF5t76IaKrlq1TFmTH9WnURdm8fUzBQ2aTlBYE5nSulGWeXOEHJCjr+212zB
2PWWGpzDvbyrGSZeWJIfcVDxQVDTAuctWUY/V7N7kH5FgXczmsuWHg4TazMbXBnmG5Zr5fN1Rw+c
VivxZh4NOXIiC97YZGbLkq+cdDCssbE9wMWGu/iGKsgCDV/WboSpMtvjq763NoRSLV+psb5Z/QbM
E9To0azVfvUOw/+FalBQC6kyLUXBLH2E9MFzkESXtRWC0yDeZYFQ1vTot3yX8wRMJNwGPiQzijep
3JvAFapQzUX3XWYB2JBmPovOIJ3HtVMc1c3Ss9BS+00eB46h0hocjrnrlf9umSmrfCabTGAAm5Mk
x5Uevaw/gNbx6EcW/yOr4cxCkDpTVTgOIPgXOV06/CpkUskBmXjVAtfb8MnFrS7nXILWuzw9R0X+
7EUyZ3cFCc6Hl90ZjsOPaSuPu5Gic03dcXRxVU57W45iji2wSgvsR0OrqDGN0NEUV5WkayxLXrKT
XysilcIwc46vm/Tzx3EzqQH2RugTanipYSSffl9kzdC00X5++DyJAUUb8nBKNWb08dg3KORt4oEJ
wJvbKNku57ianjvRQtBbX3Z4YwGv1N8efJaDiNU42ioiFBwXro1mWSxAkOLok2g/XFhvPJCQ1MJZ
z3dnH6FDLuT5+CvIjQOPVbUDvsyCP1snyt4I0JTNiijRp+8ibsqZLyNvlJomy5Iwo8iURJSgIfwr
+w5q+QbhxzKAbRARGvDUCln+X+yxJBs7uD65ZZ4N3r+NPnRAX+Eh7UGH9qVP/hQYiBqDHvAuCOy4
MoIo841oe/kCOBCscVXSD2iy8OXbJR4/LpK53ML7dbU8Iye/DTOtXvOzmpoTbeg2t1XpHM1ZEaVo
TzVmrrrf8xN+N8jqv+p8TC3bRNDeZRAAGTw5lA5/oB4CwQQyuir7iZP8C7F9m5BftP8aVkqhmz9O
Eksuv5rstz1Dv5KK7LOe7aJyQWwgP7dYxSw2Ym4F6Tz9GWQ3WwuFoM/h6jmR4/W0Qt8GB5L25pMs
w6kPEQ4XH3VK1COJTjuikOOWdrQTX1C1+bAfY/tqOGccIcDjQ0f1XTGa+kkxr5EKjsUlqXJEMZP6
/nsvGXMiWBeyCfjEK3HxMyJmJMG5GDstiXjIYL2REcwSfCsw8LI81KMT6Arr0R9Gro2unAyvho3q
6KfJj+PLKPA15PsCZenrvnDmaNbsVvEMkirmqyo83+zPNFtgO8RdJwJKFC2Sq+q7BcG8UZ0Bj0rP
yesybL5j42dqKKfvLcLKJi1U3USshoMFxaWXtRDKMnEpJo34DvOmdvV91JXsMoFRKQjsPRh62uO3
WEyevXNuoSmHf/oIodmEAYk9sRg5NtqZVxtbKrjmDsq7os51PlXL4Z+5WwSoJH40lUYC6l9EfdjE
73TmyFvVVIG5E2BP1UB+/OL9OeehbJ2aiAInRFhW9ysx5JM8oGbUvh925COm3ZBlLzcAJJToKWwA
E6qiIjXBEYt3tf4DeRgboriNkZqymbkEhbM7KzHqNh9sAouVje6gZ24jYXkQrBaYC1735lhf/QdP
AdwSCCLXd7sUjCrgty+FxDtqnP1yXNIxiIuPRgXg2H9B0my32YbIlcbI1MpFT8MLfFXAcuajxE0B
y+hewO3W0N847g/W4ZX9UnKu3hRGt26mBRHAp+WUqJjHIaPJF8oHpUTnVC0aFaiH5KHAKGvdxWvm
LMGsLZwyreMuD+J4TDXhxKtvH8w/UYWsCZQRYpm/B7XQiPkxzzK7v/dqE3hC5iqk2KqyTm3ErKg0
0WWJPQB61Tu03LNx6EuTxra3Uo7QS3RtjIy1O76C7eEItk/4OMUft/2LQoq6opdj6P7uj8Se/9Yj
ZzXLKCeiYQOdypp1+stWs6tYBXkCgvWt8FnF7iufF4BJuQHwukyYOyQpimo6vlIAChDTbqsmWhMS
dVVJgB/vAu7znPD65T6ExQk9rwKBG3amlw0no3/ajifKTneO8X5y5S+c1t2qHk5KnObvmQaPuWOU
r8m01u6ndpqTcqm73tCsQPsWEcJl/gfPRTy8jIF4zej8rms/Vto3SiOVIEAat8/KMt+qfpfGxaQF
aDyYhFXa6Lbj3/do707wekJ+WgvAKYObK3zJ93zMq++DAu5SsPPkHcdOJPxk04qfGGpy3asKazPQ
KvF2+idHz/sa2mq6CqptmOIymS06/1wR+UmYl1jh/6YbwvLWsgbwc1U1H1c471qkVoYS5C1mk9+Z
fXlCglHeOEThg2I0otZtX7TmIxcVoY9QgMHuKiC0wMRsEERmBS8/D4r5wyLv6DeXX93xCAtZhhY/
G5D/WMOqplmwSpre8vZCltOLYZyq4Mjl/+Ii7uJPX5bD2ohJL0KBBwYVEAv1S2tGi14FPu2j4kbA
/IZLm3z6NEY6i77jfW/oRHwk3UZF3WQ8MLCNbkVrinhc+SEOoQZczlkwpL3bdcTqR8xQLppKJElA
b1UkJwAA52f4cI8LBmvX4UaFYwUU16eof66MvuB0FGtTkHAe/y/cx2hIROF6ifZVQTUis3tC1CcU
fiAA8X2qiHNFqPqmwzUfbGmgZY4wl0MBxIxkbLFcH/vxOT8O2ZLi7g3mpsSEWDk5lQD8WrtXWD3Y
XB2DOewj74WobVBU9DRDJVvYUM4b633F/Z3JN/fFtsB5A8F4Kk6DO7WrgUG0H21IKApnL+TrIofr
TDoSdIUqDbEQZrBJKEhIhau8FKzg83sgEZZfzc+PZz4PwRTAgy3tibZzLj969+Iek5pm0XRaWCba
OpeD3Bxe3s9jqXNY5sQr+KNtvxpjpBFnaW5RQBQU7hXCnaVrL06CFD3PUlhEkLSCus90zGAAdvfd
sYqoTMAxi+b9bG2Z8Hbg8+lqEuKVr5qosckwXNg28DqzdI4rV7s+wTMj24EC4/8hQideRcxtdU1A
BAqyPYStAUhuEw3Ak9VA6vbSXL6209Mxo3Ki8M8wVEuXWU5F7eU0Ji+XlQXZQAvn8ktA5r558qtf
MpnpO6ZhM26fN/1dL4lIFjNxs1p2TSL0trgHuIsxikiiP/tb6AztpqRIBSYVuKbRW+56Z9PMz7Ak
nihueJYfGfY95JCCvSLBrz3iO2ioeypjAnnA02krSy4i/QutAOl+xd511TGy/d5w65EM23UaY3Gx
iiGxcF+X7f/2gM7wSo7L60EZopeFtg9FbrAmJAVbQgCs1onZVrBGVZJTxJQ1hG6eA3FJCzlVXhRg
8zPYOBDPlQzJ1HmaofYXtRenHEXBF0P3nf0ctOLvJGSkDAdVYZ9xdQM2EWSFy5NRdz/EzLKGqxok
UeFPg6Jfb24MLQQLVwQXRKsvYtd94rXJdYNste/7TrhOgUqBhdMqyjQMd+uTAg5cI9GaJH1f6lgB
pruA9YEydEmSDSkDO0J25GIkeiYQVgJZg16JqA2ye0KwyamhE/SSIYSnkSa/1mCAi3unLMA/bZLi
NJlvYFE+Umn6ZROnV1en7sVMhGxjqLmX7xLGcI9LVyH9W7WLI9aeBa1nR3Ixbt/g+Mqx17PnILwU
IcomuZaymxXIpmy8bQh33Oa4Rvo5a1bF8B64XIt/9aA/u/bg5SjNZzoEpDb8KYdFmfM0/33Do+Fx
i7+1SGls1CJy8Z/6acq+Gq1fzeBpHRSTdELwjvnXKnBdyAiAzKs+TlhPNkeaZHvW6rk4AxZ9j9li
hKHHTP4becYqKd/ltnwCG6/HF4zQV/uNKBOlnwo64y8QTyNarQLAtOKr8zPlWOtvS/QGiWJjOXRn
nx74X0h1TCNzdAuo2qT9e4w+Sjc33CzpP7c80/20aGzN4NkaHhmIhT9JwFEnmUxtNxu3TQeuqBuJ
Wf6BTB/vErdVaARbaIOBDgiKWvazIPqwHJCtopz/CTJHssMX5MmT9Ck+AahhHxZWmQaGNv9UZ1o/
EiqgPDLtEFSea0zOoZdaLz9zFv33BCBZgP5kpZRO8U0u9v0/uZAy1I4BKPJ1ft2JnzRH+Ql40D1f
CuIj8yIS1jgWnKO7msi9ECTo3Ki/u8wUYllFUH/S/vkJrjVRAgT0dzSgPh77vTDEgyVM2/s2TmkB
j8SOWw3S0tla0klTVGd1OL2R5gMUd0mYBxFgGRCv8I8t/KV/Cr/7WLoqRiGwlfNTNktq3paoh+d4
ouZKtbQvpz85OyPUl1ztfjOCjUudMFD5TZFBqiO7PHDTWvZC01uQp/OwDiVwJ+9SBGcaK3F0VLnD
BHaDE4pjSgi+S0HRADisiEL0AMlgu4XK5PF34p1dSJ3LU1HG0HqFPh5OMO/dSsflxlDHvF8Xw8qj
wIXeYwfAlUOxfqnwlA8zjZ7vQFmUWNUZsKTaMUcn7loUouV+iasM5QErRb3SC/3kEgjEwmfo0cLu
09zaUGje5GHkqvMBabQTpPFW4paUwnbIDlALwB9u73XE8ioes47wLq4oiMzJ17r4f/YyZRymE4oG
pP5QIsiYCocln8XN8+wyYdLFDd6ovabxbMlRtq8FMZR/PrLtYg+TlMJArCl9E3DXeZoyI0cVsGNP
dfAqTKmYRBnzp7ALZuW+aonfdaetUZN7/OQla2tKjTxRvd3IDyvAQBW8va/H6NWUuT24oAbf25qU
oyuS3gDQukikSj8FkTZrBSQsMADCDOUe8K5Cm314047l7WiAyq8fVe/BKEapHwcU4FDjz3LAdS1f
yjeTwNjdgxUHhaqWXbXIhMdUSvO2nVVhgjpizrho05Sx92jwmz9mMD7oLNgOPwBFKSgUHx5wBgeu
aaHqL1V0iQ6ed5KeRgtig9niFv/JTqH+ep3ErKwsMuPFrQsm7ai0fbD6hGbifx/ibUjIRisTKaPn
2Aef1KLCgvsKnjupQJoIX9Cb6W3pegwrs1Mo0+0ahP7a91IR//+gwsQ9m9KXY+2f5C7ewNEB+lSz
4pc/R+ETjmHDH3ImA2/U5LjcZ2ZCHl4iDsDku8+6wSwH4xGggL1y5I+mffHHOMP4r05H8WSfndM6
PU3HARZ40orRn36/cuQS7gBe2mNRugteq8hno73VWXZ0I9n07SVfEJgoOhoEc/bqXxlAlEkd6j4f
UnhOUl1iFMlfN3UbNdhVCjQmlcpTcRPrFw4Rqa20iPuV1tqhgJf/LqRGgioSvMYno/4Y7SUMD0Pf
RsHXyhC7L7ZVhIMF/Y/hqv07S0tKOyz1fEkCXyuliJYM70CX8zWjOLBLEcop8T7fUwx/+XC9VJ4x
AiFGIcnc9oAcr1OrrYQtJTcO9nM6oh0bSuhmhbpF5+BmtDrcB21wnRLovaULwqvtA1+cVD5S2/sZ
V1WMwqN6mo5LWNscBdYmM+GJVi1n3vLyckOYiaCag6qOQrwS/Am5DnNxC1+PgkyMVGB/tcxjEuVA
LebLEFdyvf/2hbDppkrQfcSX7m5yM+z59wpdGDofWvK+QPzFVhZkHFcwxmxlFOAJbmVXVYUV2xOh
TM5HKMdY2AKfR/ZVXGwB4TpviOsJF9xyisfz31T7pncdITJSpAl9l1ZGdMmj577UloNu+h4w75Lq
GxTVVUfXg3g2JicjFe//DkkbboQzRHFclhVdJqsT5Okve5YOF3IYlHNdwx44jv06eLWcvS9J5xbq
40eZdnmujMghEHUZhGdaDjQaaCwPnlCyetsEUlY++B2MMnmY8WlUNi4Ds+gsXRabGc3wbNKSN8EP
4f+VZe8AyXDtEMwVycRW3Sddd9swG4TA2ymIX8+HWTBZLhgaPBYV1ivmTEdgiNYaVuV63mq1JXNu
YZr75yVF/R8tZUMJlBvrTcCJv4wXErn5VN2gm8N3g7FL0k0Vnt29Q272PEnJhZ//946hbdPAZYBL
xank6kmde+VRsW0WDowPXc8A/tf+Dj3JzpxlhD2kGku4P4HmfF3U67NG898k6vJ02rrMfNExXyHU
mKsv4bxUNe4cwr/uQcJTG1MBbR8kwsNfR82AhphYH8ew711ZIvwQy5R1Ul87xEN0tYu5zzIMY+Df
CNdxdwTrIvFrdYZuKiROKph1obI3uIIMhZtZ+gFCqdvwGN/FEZfhAog1ycsY/Cn4J9PqCuSeZJiw
4M+j73jK6VnVNlPscX75rPWYZdHrOnh/CoeCxtzFraIEDubIQCtUutuY4QSx61rYc1kgn1OLjBaP
87569lssJ3c7E72BDyHX4bmMb1IfPsi30oSWP3Yy9Hg5mxCs7VDmy1gx/lFD7wAGHvCUDRwxzdal
/0DHpE/11Mo+/Wx485pzRY85/dMTvRfeRIwwt6dY+t7nHzBeRBu2lTpWxBCMvS8A+wQM3wfcmbZf
GjJQZND85sjCmISauuz28OV9zgYZupGKWfspWbhfp+8EnCT9pS1an4Pq1vOiHusWJteT/E45uZLW
mnmRGnWJ4MlFUj1+1+ZvWSmWRzW4MU6XF7T9nSB52bA4vjRTwvx8v+vZHijc79IeJCVkLTezfoie
OxOSUzP3/9sogBaF2Hn93dKdJuj+Sie99gYPj+GwU03eZbTbYkrzm92BWiXVCCuxq5MVtmqwC4vs
yxDocUmFe/aKWMxkzLJVbib61h5XeGYQ2LmrVHe+6C1pdqG5JWS+tQFahO4ReyVq8wW0Md/zZk6Q
a5ynLpSYEhvdMjOswWAe1YVKxV6bZcEmJgUaDl4vV4KWS+OoWQBRUVCS+EbjQGNvgwSKtgj0GGhJ
t18G3kIpNQ9/ZnStu2hTJkA9oyq7YtyPiYdmYFuY4uVgGZD6Kx7utL3biI2Q+VirGmxsWMh3Y8w6
AistYkZVw/NoqyPXi/MVGDc9nlOhRkCsBTUd8L21DVdcl/wx1wVzwuDRXThuqi95KG1TrqXHV8Um
f0fquj40PCD3CQVK3hq6PPE6P9ep730cRCW2E0Xk2mha27b2Z9URrv+FQ4nQa32g3GeDc0Z58xLc
99943MGRfal9zXiY0oMk3Sm//8l012EZv9p2vEh3WmT7QTgkF6oOdunyRpNMY0GSb8/9jl0Mpmvn
IwsFdnTu6i6l9sb/iRCRLSyVYXDQVTjc+ctgSHj25nMYFlPUJ40B2My0/dg85gEWVnBO8oaWWLVo
4jofMZaU8/4PqBK6pu2C9XNl2fVi2DQHNIQfca3ZwlJkXE7/yOaLB0Y1mA83HasnhkXRrA0rzNmY
Ma+JBKx/abhhSH1lu6wpDBlZvVXz4Q0FjzSVSlPxmMMJI5u3gHvPxWXtqeG2v0hPjvd+luFb03Tp
55YP0/i6GlYmi2gQPkZWLc6TmpVnIoDo1NXuOviTPreLCp7aeVhRiFsca9QUyUHYEsRZrdPTiX0z
1xfOmuAcZaQRh0IFeLZIgsWFws70gWg29kJM+5ILWWbT45lXTAMUgRmH4TeFCFRcxd84O2wauink
TodajWmtH8bpN+fWRXkV5Np67C2IoinxPi9UnG2mw7DTzPmsB4rshoKVFJKAtoT92WIUGf9ax2D7
+Y4P9RigrfhUnY67CHwYpVPdhk4nyq+Dh3OQTzNZnjATp6y0hT13kEEOYiflc2OKFuXUyYnHwcPk
O0N6BR1gDHBTpz4iZ1hSSroWlfY6rrouIPsng+wDrWJWyxdnfCp8t5gLfL//G8PAV3Rz9FvIr1Xk
dbQeCJ+k7JkwWWjiRduffEMPK5qn4cvZHhckP1Pytha5XHf1NhFnHv5rUXy3469uX92cuquEkQVK
knHv1yeWki0yx02z8+Ly7bFgWwf5J+kAO5xW9w1+tKo2VEYcR8HGplaaNK6SPh32228biNM/FznS
63VrJ217tk6yp1TQVRM4x9huNU5kJ1Zjmnv1AvgdugLSs7CP3BeSUcu4tAQ9zSVJNMC8BtHibEia
Cfzc7+zrC12YsQixGRqtqjJMPGMTRSZMajcFx5qvyLGvjMw9CjDPXzAAnFqS5LriEEh/C9ukX8Nz
MvMvwcpC3nAymIV2rqVFG1EsJxDSVC6vvqMNSWYlY7yPk6tXs/GZFzQ0OsThl+lHV/GFCUkQOQuP
7Rh4z/BnuMjHUNMvuBQ5au6dDyFV9Irnwk2klSdpYVe1sbSXJmU8yhfvYYQLWSNvX/RLuRurFkU+
K8MojBL/U3ajDrI/i/0H41G0F3baCacQMDXjNZetJzm8xzz7xfO4Ct7I6/kNsWCST3Y9cSCTnSWT
xjuI9YLFo7EI6DVIjUyyOcgGeMQr2mtQ1H4MIaWI+5dHDAqJrLqTKxx7vzQtwEOxOB703iE3+Vd8
1PAZYdza+H6UTIR+LwTkcDPbB+XJGvDIxJTtMD1bYbZ13wKXG6JPgow+N3ZKwE0VYQM1GCcC/BNI
+bTtLeENvSRTZNFxxRLgLwacNmAyrvNf5ceAvnUBZTbv1QRnfqn/uq/gTarN16w7YgLCa1wldcM4
8GHf3T2RSoCQ+csjzEo3Dt1mYGob+9mxCZm6ASRcnMDPJShDU1HI7xi06BgsEuovXRHcrupDO3gt
FSxOlkTZY6vYLfYANFFu84wck4OSCah88LSm5mkul/YE1HASXH2BmvnYKr0bCtALf96hyki9S1mg
ejD8JQtnOC1UEGbvBOHiGbBSOKLNiDFXbqVBkOrtBF8F1Ks8YzDDmBLlRKUWIhgqwbu2GInt5F3R
pPi2pN80ynH0cgM7kuDkgxLvItpBR4/AL0EkckjJRqa3AMH1ViAWCniJILGGRKlkedYYy6oAiB0W
ynUZ/+LuBh72bme0QjbjePd3iNnjjDo5Ca8v+zi2zwGiAtUhiy5okAQ9abQcTWHL31LhEw5rsU0q
Lp3SocZLKUqpR3O/pHZOt76utSt7Aj8U7I29iCTHX9ohCXeKUZ3Ya/hNe7DdVY87c/4d1oT+P7fb
qUQA9IaMSIgqo6y9jwnthH83EAz1rylGei5cFg2Gte4mUbRQsihWcvRKfl6utXDKPnwggPNNsdIj
Ncml1FATEbNISM945eE/y5aePqvXJj1jpFcfxZlWDVNXcHusBU9dG3/vPpKn52Wa3V23gXzyFjgZ
1o9XgWyw3mb5DEsaodNTeg+PorFFzXr8yJwf5ywge3ZubiOM8NJDQ/qLEeAEjeVNHZGS5/otlKA3
MF9K9AXO6ICLn4Tz6PSLDyUPG2NbmXQ/PQF2fq//daEKZVCK9diU0gFk8LQwFpbC4pZnsx+qYOyd
ZKUuPsqX4D4VBy9tyFj0MZTNaSjuv6NGLW9oItxctYoWZWnZPkUzXDugm6JuxnQh8f/m57FSnlu5
u5+6MBgwP8odgBctKK2ODWGEMrFMgm08u0CdtR+A9mLY2xqKo9ETswuRirrk56f+KLeAHEaIOlms
36DFKamAPV7I3PMCD3FAlj8iGslwN2ViZccmqvrslnMbsWIc6haBSf8iXh+ORB62djLUNLFhl6BH
WUgOA0BbECVWYF2y0yA2EIUJPtV3/ktGMwowQDNm09zSFnTHruA5o6tpG1W96HmB5NlgZ/mm+Tng
tccr/VqlvYFCxBvSG/qDzbWfAVoG5qBPTW6UF984imCTNOzu4WFwzeEC+ZCZSvt7xob5DQch6ypd
em4tjSXz3YIbgtsiGvvxSOx7e+iUEmAo1SQtKrTRpF53wcyNzpoQ2g9Og3QlULUiQ6WnDO6BMmdI
/jrrpa+Gy1vvg9SxtGPjtlqleLW80evC5jKZNMiG2ISQzKUrlcvovKmFbtRZts18K+PB2JpUodn/
PCOgtxN8Y/bfHn+YD4FYwvY2a8Px3yJRxYcuLkttcHS/pLAIG9p8BcpuSjaO1h/YwLCisuJh7fLN
ujwwa1SZiZInWxWuh6EQa8Ww4zgZm9fBAcnyuEsFqd2hu06CHseKsiuEaaMvBam0xrzSil+XefBX
Jxh+ILNxUx/4mnPrtWQfXd3rNyVyEp5XkwizidEk07zqfGV6EycW1UjCA3VYH470BpEKg8/NzaUP
OtVgqRojDs/BMrSYzBGvSKSqrWH8M+qwEf5NFjiFLy1/iXf7iqaluymngJFODkxmJNENBrfAlGFh
IOgYeJuv9GkdtZHkC2cFc50gOeCsenWGy+HGy5av+pxMR8pj/eYBkymoFWFsX7TTPZklPhjxL8nc
oBvdA4KS61lLqvVRA1CTZErR+nfCwf5TngYpbTx21d52fKJMvW/Du9B7Qg9/ZwlYqmAFosqE/LNF
GJXYn8DEz6u2cv2HOhjDzti+V/oL5SIBABEX8ygm5h4XLmN3lSgAZjOmT4D4yuPLev9Fq/qK+12G
cylzMSUAkSbrkQHO2zFdTmV0EtTV79fanImgmVjSUjj0fsR2YsazXIpk0CG75Q0Y9OMKaio5nKfG
G6A3kF1ZMrrfDuXKMd/fUp92206qwfQQTKpAfH2Mqwyfze0NBYjSnjutGGDAhAttH0Zjj1OBnBwQ
a1l0yH2Syq9NP8rdn2BiS+opW0rA25DZ4uA08iPsAPJfvmgpfCgj42tt6dEFExTDtbKhq2h4J588
xrQtkSr5iw7LsSwI8fEc7rWgoXaS2UOevwCx43cWDwtGs/I/HApgBz5ngDRHA4BsoU60KloC7dPc
smn4UBMXL1Rl1zoZ45fgQNZjCIZ2rWepwQbzELjaDnWECzEePeBV58Uv6NAfXwzuYA3WV4QP6CRW
atEiqjbovDi0iNDgW3FsjXUtOE6mOh+cGNOIE6i2JAsgGXG37+7mm3Y9R5P0FeWKSWbenQoR+GEW
BznkzpDKMX7NYT/YZ3w6/Sw1hUPk6Nd8qEs1sgcSr+6RWAL63BCWCQFsw8zj0WHbeEvnnmxFvXwZ
VTe8+II49SUhFQbX2Mg+hokf3PlnslmBE25/a+irZYJ6HaNo/7PHOheCdjEIcKlblH2PPW8MRa9E
9J47JZLcA6MzszSDmv0nVSsxHx7YqCDBTgdr+Hl7wGkcoGCSq60b48WWo/Kvy0LDmdz+90g7BPBy
mKDvj4NdLUfw8hj1+APQUPvu73gwW0Bx7HOfZ5KI11xczh5Mrs162wuqUgAbJlCci5wQFB5vDCQT
57sJrcFEh1U+PUot0Z/rwLFxrkDovPbBOa2V/mzW8TpYf5i/lrP6mq0FduwaYlFdrx9Po/ZO03fQ
zlPUb+w0W9gvthtOLBcKDjeEPXe/ANR4CFsEOC+YJ0zFsZvb6pwKKPnD3b9U+LuE9oZc9A2pjt4U
dVRiMU3/KDb7aCBbdPzHlRr+3vnN134RmVgzyK/0sDMoyt4RVK+lIMq9C1ETS6fAhbTPbOri/D0h
F0sCL4mbCr+f+XR7OPpDfFVf4PVXZ7mI9pCa7FZLmK8MpPKOO7NtaJfevI8/I2G9i/2s/IMGWbYu
i5h7Pu2Mvm4VMrD1bGkz5WcHKYVpIv1OFlUHE6q6rOLqeM0cgygy6zrUdli42+hYx/F+2YxILyHA
7T27USYDh3j/WqWJ9bezzxjG5kctnFeSfQ/n+UTzjo5wJPE9imqzx5go/mb4LuNLcGjuP1tHZ2oh
sjDtqzi40PZozzk9/uAdmywEs0QgPykM5w3ikZtFmNiKhjsdMKbdPB3J8HCQ8RRqrVw+BSH1vTpU
IPHhikotgq+WlwiMTavA/5DhNez5+zGhRExWLfi0Ntw5frminvQJMfVAZXwf/b+mY8QYqopwo0gB
FG/5ZLfukRmDbn5YBYdgiN3eDzNXg8hQ8LjPuZ/jfxda3vvffmpYw9zDdCfbhtWcopOGMcoFKcr7
NO0brUHKhvLCmdA86Rp3x2QVnh0OcPBBH11m6WQounqzmciHNi/4QYTeTuFcNe/rV7qc3BtXk5T2
Hkh/f+mBdLX9gwiQEoXVy/3CaW3EKDZaGSVNjdWGskYoD5sLld6Cd5fXHa8F4H/PuRVgUet/8HaC
bIZFF12SQ/e9UDbKCGjRhHa2lYwqdxCDij0VgpyptrwqlTQdxOFKfndrmLE3AsH9jZ9uOo+RHj75
OYq/+uknTHzKjqdS5Wa8du5/yfwBhBXSDRIc9Zzt6a22omVtIVGrH0DF9F4cRqnOYYqUhpenBKIu
1YXUX0ztK3uE+uBvi0ihSWVJwKGB+QuFLOitmbb8XMST8Y+OjrCGjerGxUwCTB97nTcvsU91XhPN
qp4GPNjkxmnAKT5nht/2XNGjiLZla5j0wSUGXCSTRoOxFZkxEpX3g48D9tB2HQS/zKSapqZ1dmPx
8IKYMpu78KJF0bHp8JwPc1+MZXGpfOBh+ZEmywBcHw572zaVudBYngXkUpgoyOYnMS79r5OOhAG9
j8YbXnqaT/Sh0KQkVU1UBSJmfCwkXeCtIrt2XA53fESClRObodz1GiVKjYyeu9RzG6Qg9MjoTi2f
34c0k+yVOpqVwuYqO6U8bwxHAM19BWxk9CUcUV+0f8mGTdxcq07wgzNO9DCaIfNoay0gXHCvHk+P
1U6qeV1Hqq1RY4m41kKY5Q+xqtK00Z3HphZKv93cfb4wwATZPmSV6zRkzMCY1dVzRYMBCJjGiCzx
IQJ5ImXfa9fSbEkgNQ1UVG0/AnNQH1DtSDsLbBMfDL+FuXro+qrIZQPkYmWqmL1ayOpAaqfoq7KQ
4qPYHWkjJ6F5FlUcmLXocysF8Q63XBw36hdmGEpqEqWCONnXixvsZsTwNBVI3TvR7R0i7MaY6f+G
SpUac4aSUvrau+NvJ+sn6WsWML/bQS7PntkYbpOU3qIROqDdiXrrO8UL24eJjM6esXaJGmqGhxef
PKS73G5azTVt16d7HNitDDS5LJW4jIJEDJbY1O+M/vTmAotOAlLJ13ePmSGhbTM1TrBeom5dRcwQ
s8coJkdCsc6E5ezQ8Y4Q0lSsRHbIZZ54YLEywQBWNYgt95Lhdnh+PZVYWLHnVhRN2kJtQ+FtRxAs
arDzB82VdtqklP7N4ZDxkkPMU/V6KzEP0GzRqcZMxjVY3KSI1k72/Vj8G8OWIrSEBnU+xPU+2gXW
+WnDPKJ8Y7uv82d1fPEp5z1nb+opuG2qRZTgsIdNuPXuSlr1P4kPYvAhBEldjhU/O9hsG+IX5Yrx
MqFVtxDGuO77SST4eJW2BVnRxQXSNtEEXOxpREC+gF0XHcyrtKqkYZ58QsNX9e2D4PFYI2wJNmx4
UIvMZTp7dnb5z45xSXdsIbpqaE2SdNwXX78B/74RVTKymz4ZEJwPOcIkLoOpcjZJS9KyNakHfxli
P66/hH5XWsZ7kRJ+lE9nyTYeusfLrXDWiDOyy7r7g6tveovzFnBBUZWYewk2x0gBVe54ltpOOXX5
qROW0cPpde2iN5DWTuYqy9c6UkB5m006tQycNE5Md9aksuKkbR/zRfGowI+L9DTKhCk+ePTekT18
+Owc73D/p0H9XsInWUA8/YrIaOlnlZiAwiiTgh7c11pL34a6cUQTfsLEefYkY9uN2KP6xZKja66P
eLolTZAVCosGZeTpMHjvbvLJn1MpxqrzU15R8bRhX+GtGu1Wdo2Mb1mI1ckd1Sr0HtbjGGqUuiHM
SXfRYUluxMpMLP9wznsBy10j8IHu9U2XOtLst8zGMtczeE2ERMYZqVKXMbA8HUHy+Yp2V+eZUrti
OpTxlWvUtr65eD9fcKgaxkvN5giu5HaOn9RqTo3mtbBE6nOGk0TTsYdoXhHLxytTfGqPX3KyXbeR
DM31zo+nbXIHXoLSYT0yOIl3hhqHotT5WLyTl4YdmRLbXjxzwaevSaqJrqLtwrMsJOsPk3tih2aD
js/lEybuzyS2oCuoE+15LdmGujLU80afX9zrtpWYQKeGcHja28lrOO1A9+un3gzKLicceTK0k1mV
QBfKPesHC07gBOUp5K2lcI5L7/S7PS1NTSA2Xq0hThAsRGE1K9Ag2p59VjF32IGBXGOsscuB3nK7
CkJ7rBW70n1iV6Y1f+O1upUCtvEQ5b56JXL5LQYXL+22BUrBU4Nz3/G5CH3AxrO2TmAmwQgl9XrN
+F4H5Cj+PZJdhyTflBdmavOV4tmS9iXSiSZ62l+WrZQLoURpySANiOpRTrEzZtQ5oCyM+ns4HwAZ
+XuFIktE8bFNpI3mNGkTOpUX9eSeQ8rf4+3XlRYdpgzCiGFN0D85n+vgzVC9dguGdHduBS1LGw7P
ooskEeecBbipAkqoWGJL+sTTbTsOEC0VqIACQGsK6h+DJawBQFeR3iZSSZZiQwMuIqsWwl3eQoK3
4A3TNsXH8Cv1XtaLGM9VniZTf9M9CKmQR7v6cqoMnfXsc0IgROPIewUqbamORpbgOikOR7dSbTZc
fEjEdJXqwkpZH0dHmfa1bRV3gc/pAqvN2oXe/opz7azr97XnDEcKMoqyXm3XhXIzvCGxFl0qfmVL
hEdtgiNbezuhKYXOoQkLanp/Fw8wiVlkQ2nKJnmyLNQ9tA3pvyfhHsciYOMVywX7lJHGHviFdIJl
9oXVDBsgnWzFZUTI+i9ofp+8gtdi8THBNpN3pKLfoJpae6DpJdBipvUa78X7unQfHu5zYntlj+95
QHwJ8g56kiy4i9X6NSNrrMzrus3AVHnrrAytpCzi83e3gid3g+kMWzPOZpyWvirFIdkMAliBg+8E
iJijH70EZKCZ8znrTDkncHhG4/Ncpm3JQ8MLWjhIiXgOzcTZ5/RqQ+froy+cVVARQtVK9I1izxlp
Ka5Yae3tz+zLvkZX6mq+BZqq9hZ/qA33RHqdvJkSyXbi287fRMP0e6AiwINr4lgFD1ZfBjJsVokB
xv8VcdYNq2xinsRy3OKbQCQvLMk4wKfsNYDlrcdQ2jnYX3ZPmXrTPEGQ0JGlxYqFcnSDLzGH52jG
lzdMMBCYuft/YRz1XS05bskkrlLmI8y44fTPnFrfoLe18tJnyHNa+28RL9lYYk36zr5cVhPaoJic
xnq7/f8MdwzXCO+96Uvvhd+eFD6X18BAVqMrgix6+SBsS2drZLGpzMkmsGhg4dbvT7BpsmQe0obY
s7kPxFw2Cb2IQBUEm1+xe5VncX20/zpw6ICFCDyLU2NleqfhuWjVk4zlXwmLcsI9CRpaZgFyygSd
KgKz7wmFElyW5HL03MYvOARH+7L6pQfXp6WO+Jlx+hwea2ddxHCdfBzfNLLjic57suspzJpraXg7
tmF+KOOzkr5O52EEjg3YRmrM4pLXzbMLz0H6uG7qWEm1pcs/17sq92vGrvlWvbnDmirJtIaddGiv
oXTU5OtO1/N1CsmlaGuOtGRNlwLLeCVXw0f9jbszjay0HwjmKUYeQ83zNa5abSbGoYjyVpmp+jim
tpbQS1HlPxqPn433ntOkmhhvUtrpwcP64KQid7HelE9Y9niQH7xXHfRrXrq54kzSJUzMakX0PbI4
VGbZ16SDT8RnoX2xNE1ZJ/6nRI9Vn7NnqgTAKqZtEfHwgD2Bc1mlQzf5Vlv7hNQNcVdlC23FriPz
73cuSwwiglXzBm3zxclDPI524jpFgGfwccKlvCXxkz4AqaV7ydJD3/NPm7CjFOk7RmPKE7ziaPW3
Efzwe33lgRJVhBXVs5xKnjS+jJPdK9rEPeCsaTq5yv6DPKC0bL8OesFx7XsJWu6HiJ9A3ZAuEnSe
zrdhINQKRCwMm9kRvwBjgtGe4itIWGGS3zg9lzAWFk06Sj7JjpIkM+rJAP1WyZRSTZP+TVfC/sny
+x+nRl5W2p8nVX+eSvRDzvYxfmA7e2wM3nPfNR1IXw4nU/Mh3FGxVLtnTOH0RPsWNblAASTHozmJ
96Y5z24EHZXqVjYGuziPjp9jkNoXWlDOnan0MGNemjqH8rbtjU81Qgt4GHzNygEMhEX0kM9UAseq
jToO+tnIIseORHjGYhvTf+4nDo93P6IBMXOmNkiAn+dus5nZjGGT0ADU2KNfnIRBzC/EnQrvI3Th
hriBBTg0pIYwmoqI9UVjoNpaacCq60AgnRffiuUJreNVOtqpXu5dwuLGpROXObGG0Txd0Xs9rh0c
haId00wGc9ZUTVb0MczCmGFOqozM6jFgKvSWQYAr4t8KFRW39gcu4Km1f6nfDqMFrUUY5/Por81v
KwERl5SqqRfwyNEpPyytupPGykZnfS15bBTcAvUpX47YoxvD5SwvER1RI2IQ8suVOB4KiB7mYiS/
M5r+0LB6sy+Murv2mR9JfMVLdL/V09cTF6Msq2lj1hfB7whUE9eh+0C6mRLugUs/8WPbIoyWMJ1P
Z7bE7E5lNjE1H3JsMA6dUMq+mKwIfE1Y5UtlGn4lTRdqs1STxZ4Qum0zPB1L/biuzHB04RomVByc
s1OiiEcy+zSQl0ISxi3cfic9pV8w9BLB4+njcgFbDle0RvGgAOQ9vGzB9f0uo3KXzwTq7ghW4zG9
R998H+1pluo96Ar4KA+3fHTV7SO0Ii0AHLnDMDATkS5u9j5hRa97uA9Y+jlIctIcoIMV0EDA8Wwt
p09tIdk3JolIZDQtsqWb4pJXo+OKR0ZKSEQS1XkJYWdb97nB3SftLmDV2MUk9yAUkQqpxIsVvTAT
Sw6x80opdQHpWkp4RNOyBaGJeMbuets/uis7ZQqf7Vo5g/R6ZZu9+/87sGt8FmApjajcgU3Spk80
GGG0lbJoShDQNJJBBO9UZh2+2+huy5T9qaZhnTLBAveEz/cxFXAuCSTmzn0hOACd1kKMvKHuMv0U
oq1CZ7nay/r5TUHXdLm9PTRYulTnF35Lq0l89Hl+MvKsg6NTo8/z76+3zVnkW9R0goLLw+eESgFa
xxMbJVMJZv2vQjLyZVhx4iC/2ZXWGoiZizaQTGuWpefehr7NzBvdSbeEmhXogBaqB9wGUMHlRJfe
eNw5JwrMI9KN8YJPvxoHtQlk+DGPxFVZxAbXhSfeZxck7hEPkik74gn/NJKwARgbpBZ8AdfSkqB7
lm5pmJb/ydQxPGoAYiWe3TLzaAjOu82cSX3fgGUq74s5IowEe5G8xwsCkWnJ0YN8occnI7Aw3Yv3
2jn3dSI8/SSIcRTpbF17IiZ3vy+hjXc5GdkkhqjOaxvEmTF3fnk7jE18ZE3MQTTC/QelFsIhLVwO
32XaTcwswJJ1EsWLco3c1qtqB4qrXIpTpaf3rTsath+7Rp/uWGxU70PdIhTflHtMCbaT44N+OaKB
aAZlwBRFOkfU4xUuO9A6TCcVsv8P0BW+s4iHwKqxU2yrLamyYdperYB6qZafYg3fxKZR1TGisgd1
BG6u9+ZY3F1PuRn8xBfmFTEeulTdKBffR3+JktT9CjzgtiV2lWHulrmPE9YyJOF89aAeUY/5rXqL
sx/o1XxOn03X/ZRsFsrRVDCw2mv3jX+rNvnRS7Jmq3CO7ayTnAihW4fhQ5OA+JFGhy7Wy2S64atY
4P1yzzsfY7rXZvCSjNodM8CTvj8DPEAMa9OAF8tAqv8uEHUPPFbwk0E2wjhaUYulPmroRAuIhRZr
KvAisS6LCjVsHlKCkQxyPEHB7EdZEtiLfnj/5on74lGSoSwAaZ2F3M7t2QGM88ffiWg3v9TtePwB
WRW1oEpVfj4YwAZRTQ2pFl1RRIflO56zKcMJrEEDmsCWCbe3RjLvP0EKp64mU5fFNYm3rNuQXsZQ
SN6dUTiMzB5OkzR/jL/HlT0oL1Dgr/DZe+I82pEoCc+e7Vw1chfwHQQoC6w8meSlfQ8TMOMPlG8T
YXvdSLnkLbliAx8FwIA/OGgu10gFMLwbCnEG0yuHejLkJdQYSbzDTxViGht61raI179NrswY5yTZ
QbwRoPRSeqZ8BneizOdeS1/dtMA14/lfK64B7HYNEu3/oRJrnhpoVc9JoZZkR9xNsg35Q9raqOxM
zWGAMaFWTxx5qYd+tEvcQT7qiPHMkXvoULbXMcj/khsJLwntxFDOKHqdoJHxZpLcrQ/WHy9c7ngb
dgDYgE+zmTb+192FolmQxvLLd/sMdU2Gjr96ogneS6DdTT5ec6larOg2Zc53Mh636qDSnD5OiQaM
UQclRZ27HdIhkAQQPDIkn7DK9/xsmz+wqAMeM/n49kS5ClqBX8sfjupSpoVfP6Qdj/P/f35aQLx0
RYrxDZ0WSJIkXB1x+86gbjvbV4qz2110RcyEjU+6ZYbDzmJKGnA1yifEZmLCFNaVtH/XyalUfxKQ
4V2bkYGVLQrAaoCgX/0jvqdGY8dIcnZsHA/EZOMYfav+OWhbVJhREhiQDsIxgMNZ8SNlufwlluCY
+n/yF/ANtZmmfhVTIW9HPQ800rktJYVWntvgNLuFTkzibcPhqAQg1oHXGlVdZWs7lOfYp75zXZrY
pwAyJEOsv8lo9BpRUUNwGqziWwScsl8IPzaIlXc/nHrrsCUb3jl5yiVxdNS36KJEmBfSpncefjl0
h1DgTRioIsnRKZj1DSzJapMhqMErcXNeGuNoamxhphSCRt4i5d6lxF9c4OHzpNjxABDjuIWEhDFO
ZGN8+VAh/m4IvyBptfgxFbHntoBd2Z6sMkDFOyyxSYgZ5dZJTt/L+T6VXBlE1k8xC2Ew8s061Zgl
nRfaSg4vQFnkyx1ntDRtoMLgRJOxdvUzeguUUp/EHoxSmMrioManP/EVPECXPeKzyJ330h4RTLPg
u4zq5XTygA/lVTy0fl7oW6GpUsuvVbXizXRG7nDVchaDRAtgn/3n7UcQmV68qq0wQ9F8TTcKSgKJ
oYQqVi0nM8jMVNBNqR2Q/slJ8D8MbSTA7D9AX6gitsiwG4ADrA/TUCLdQU3ywpyufEB73kQQYJO1
hSTMM12UtJp9Rf55NSu6FodchMK/LIteUpeVNefDLDZpmWQ1r98W5LuOadDkGQKrhO6j9gor5Z/6
SYbOrIAn4ZeaDoTwszSi5Y0sgxhh0SmnN6lU5Jn4EMxphVQpS4zjT0uriWGXCzxRDC4Qgb4puHuf
u+lCBo5VQWh+NVqF9X/xFBn8w5s9U0X2rxf0GuNBTqbvbHmyAAvMTkA5tFBX/csXywRzlBjez5cj
VR6PCcpONgFKW9PI9zvUK2NOaN3p2+XRi+zQihBcZNuz0oxWvkF+YN8+eOGxPrVMryg+/kQITKDl
2/T7l8fisAmek+kbwy6cEmY1vHvx2PJqtCoZKXlR+cpNC22AsgVo4gyRxJ6xtcP7xd7Nyog25usj
3eWY72+TWdyauxjci8r/sFfMU/iUdDzNORXRreMbKM8tAZjJaYyZmpuuRiTTYOGnC9StggR7A2So
AyRATpI6DXMSE2ecEF5lXXNECeWoOp6FavEPbavh9BD38H+9GgN40Jc+m3UIFss2yr0HLHppmBMm
djmPbg13EzN58CScwvnHN38z8V6K0h3w635HJseVeC7HlpNgChRunjQbaMeCMeODS4a5BMF1u7GX
24nk2GoVnfPAp47sH5z+dU4tUBIhSCJhzXm2pXGnaLF3imr2mVpR9nvzT9viOPa5S/lancYQkgqA
zgURw8DdAOQzkzQWS7exzkM3rgdAT+Z2rXgA3O+ATSNSLwxvcGj7L+JtN1ikitu3eFydpTiUWBo9
kgutldC8QPRxOZy9QSBqFG+Sf1ZHfrgn6x7GeKst+U0+CYIrmhVXnp1MA1KCc0Fz6DyzTHuz0+UP
3zOXYdzZiheHflHi1kehnb0hZSpRI2EcoEazbhpyGgn2ZwWLyr5uoekJLpF2I81V8YMg2+NGC55D
DAZU4miwJifrWZoJZ743Yh0r5/S6OqmRpahEyR1FWL2tOARC8Q/kavJ/U3LiJZwPnqhYP0gnA8x+
VFPvpBtsL8len5HYRRmlEnH9Q9rSRHSQqMY9Dm9IkdqVpfkqP5bonNi0AaL4CHQyKBZH9Lm7Tclo
VUA0iuHclvDDADcV4K5QCt+CLVe0behXNjxQ91cjMLmHWIW4Ba3a8r6vikMFNZ/YGooGE5iR8SkD
VqAoVD3dQQCX/QcjEU/zviEKk5tJDrPW5LmAJhqrJ8N66mG7e0Le4Su/RzwHNnLA2qD5TKE+0QWX
ZZ0zeGdfdiyreSLwtlNyIb4FsxGMVO9rX2IUDEG1W0egh936BxVBuIxAotj6kWye+mJ4ERGDYJmb
UG3u1prF1cVC/rzhaDhx/bUWC1SzmwUTxKW9gLRBQNXox2jRhpwLB2NaMbJh71x7NZjhbepbTgUa
Tkhupe2WP+FD3HXXmRPlbsgJcJuGqmG7LQ1f6mpV53ThqR9PFZgGtU8Z3IauTzwTQYBl+6CgY3tp
aN2nGZYwie0AKC4gkX0GmYUPb2fHDEUVXoQRNaEdJIXfjVWXwGRONW603yy+WqbLHBNXaaPLHNFP
KbI/9XmdGf7X+ot93L5zZ326RALxawNquQO8IPkCvVu82q0r/1tmgyXHWB28LAVo2L8QnyMitDO5
srihBl3GfAcU3jMRt+Qfc8Pnuq61xEp/W7+qjRr1sGk9BtW7vghqDq2d3ZE3ov0/ckRkRpjENO3F
3CQCf6y9vy78ID2dFyh0eQ4GAsWos9fiFfsYat+WLeyI5PKgkXtSLhbEtf9UpUUnkMs+07zrPCoR
66DaiE8M7ufZHmuwpeUMoJOCamf4jAvh4z4R/I8w3DHupUeLP4Mp/vqUElWzi1U7308OLqkAMk4H
CNg6nAKlMramoFIkJ6kxBaaRGzfoCP+ReNA+uGOBoab3WzEtPS/Vrs14dgHKGfByM4pyuLUUEp9b
mskNAVOPa9Cn5JjrSG/2VFsh8TwltBZJofw7/cYi7RGU0bPKo76/B9kD27TeZszdrAEfIO9lcM5D
39ciTzsljVfpBWqdTZ+SFCaOlUdxLw8N7jOFQ9hww8QM6zg8xLC3Jtjqp+wNaackE8UVNYP/WGpo
WphdrNrUqM8f41cmLwCJ8ZpyiNWlqyIDnypUpnSqctKhI8jtUeznVpeo+a1Sm2s9TodPYycOMpDP
xwgFBE7dN1ymBMuLmJpRXhyLVAQ+dFWcyKpE9gchqXZQryXTPWDjlHfWS12N6eVOMPG0REn8A9yj
2H0hVJmX/0QV/MockFqL4rf2DaUg4U1QCZB6o3xzvXpYSO7Au/W3LQlIreIhOvR+VFzMO85ZdPKO
k8rie+wGIBmOrEGPS/DoqfCeZ3Uspd7niIqc1/zki7b+XX0cWnGW8byjL8kwHeeV90mulK7Pdwz/
XZfOs/dp7aDMW6EJwLkw1uv9EErmOl9oNAh8tUqZbc1cR2pAm882wyaReLDgfRCTJ8fgWxaeDuYr
RvmGOB1MyhmlaOZGS3UUhT1V+ZHbHs9Sn38t6Cnw0rlvoJIYmwr7GBzvsDlWLbZ468J4tmp4Uc0k
W3o8EqZqxPTLAdBd5bnZ6hnTIN5fhZRllCcDgLB3GDy1iCVak3q3zYttk60H6tkdNyRmXAJQIsrz
JuOSnpkJkAZUcmDdrhk6TmhW9u7B9xikjiQ4av8I/add21e/fXuDpIU77+U+ApS0YRxSYobWf2b6
6gXluUpfBruO2S7dTYZV8yGw3SpwuGTQcqxKzZvqsNU03qb0mkMdMLJlFdCXy0J2FJ+X9IToZr7R
HSXe886MYbw22DVqL4WHrtEMNb3m9FOxGERn5rByNaPZ6IE+NEnB1asRxpn41c+Zmo3lcL5OMDGF
DvSaKdXBG0irE0BUn6JAUEbKmwXJSf7QaXXM1/Qx/b532A3R4/hBNgdkclbUd1wn3ShYDDX2zOqr
/VQIE2lcrXg957GRh6pRxCDd/FR8/N+7Q17lKu6LJrktZOPRjNS82a5uj2hQEmMcWFQnbqa5S2/y
jKG1mbjqMLVEt5puMQ9IerhwKvnGhZGhYRZ4kuagZ5GVIhrSc+B1s/aE3Bca8krqZATTAfK78K2q
fEoc+LKGby0Pdsu1AxA1y8rDQ+ZcOg1ash5e1GhsfCN2iMp15RkSYNM22/RmWiQtAWUkJpK8lH4O
3K/cc/+2zjaS3p/uWzOPiR5hGhucz/6TE8gUIro02m43u8XuMxlsSE/c/X8WW9kiNO3R1KC1utkp
cUIZJYvR5Fhx9ppJyxHi0IAlV3gk/SIS0VaWdDGQAGBFMZ9Vy+1GoaFg/8Jk+OyB0XaCdkoOhNQM
1xyWiluZfUbmV2gmceoTn856Gv0nayEmVsMHwMeJmyds551NTzxngyWxN6XLHPFsNyk8ep1SpbrZ
aAgxSCph4b+cLQo4XmWh2w4Lvn+VlgbnrbD3Nq5dh5HSCmK8g8GW0eOeufZIG41YfO3hudS3ClPq
KlpIZyw+K6Nd16bE39VVtTMtA1iX221t+kqqlGDcLubri04LuNm2cS8ClZDtMKY0JzHUXi8GTrMJ
oKJk82DAhP370L2Y6WpMEoml8R/tPfSpb1/erJyOC9OPclB4+F+Tq4hB4vnedYdfFEq6eLKcgYAx
DIxfLdeUXvQtgFcDhdOeOEBokBegHvkklAE95qNpQIhRSTJqOTi/b/op7N7YqZnGQo5lIuDKZLhU
OH5C4QEAN+0psnO34RfRREza9D8DPkdKv+FoodBy78VUphmy5Y4b9mLekRROKx6tgZRIJeN5SMWu
pbN64ZYaMJIznlW6YH3p2aA8Ray0ijNQNrSXXXBYpGIfmSLApiPLh92t55/kVGjgZEaeoIjzmpc2
U8tkD6BOgbDMSqGYOsBFihRc3cGjgsGjhKJhDavd4jAqO9NXJnjEatZ9da+Shgw7w6AgeIHgFqL2
SF3r4a3cx3OZD9+ITK4zKwOaJn5wf3Iryg8XvAiBR+UGiA+p+5rICEshfgBnXw/rPZ2zWT3PG/UE
7mmmJbl3FabQdH3vUupK+Ka6EuPUQRSCmOSeGpTX2BtigFuW9F8uonPwX7xOug3eII2OLr8o7WHO
6FjTPUk1I8CwA3w5XtotOGrSSuhJ/GevsyIn60X6FwqKAqJ7kjI8dcW9tuVT0l2Gzyi0e7oLuOqG
hAPaBy60lW7AiIYPFPw5nxp0mMR7oL+rNPLfOMfeivfwoLbDX01w9ntBrm/Q/61g4L8e4d8Ee/UD
23SP/NE0G/tSQHpw2c80W2xflYwYrsSRAD/1Zlwq/+JSCs8OM/qh06uOjgctzJCNk92mlMGwf+9c
BI3FY+pt/bZh8xSi1a3WbYIgN56k4uPaZyR2efnW1wHDKx9SnXtQ5JDcJFvbh8GY8VM4bgTQ8Uh3
saYRrVFTMh7PRCA8qNSHsSYq+XGIH2RvPzMI0UJM3oOIdiuFDNvWOodlPibjrbN77dW9gm7angoc
56TU11iUAd3eNPfzmCytx1Tox0sOu3cS8FjSRtJsS6znOHfVL+DHmHtNhxmLVdYbb4H77y514+Zh
SLYztdmN11kxpqII6ASC/SzyZSK8rcN6oMvF/4YC16HhteLDuWOTUhe66ZejiAlJKCQXOt4m6dH1
0Kuo7uniCNd39D9ijhFRZYqVTAtKNPZ3RSgokmzKb2QNt0fiv+oRk6cZmZ6CPSyo6SYqpso48b0q
yP/Qe7wer2I4QkTKN56jbcXXxxfouDKNEvyvyBDGDDTbHvwUio4cBdKaNEjsOYBvWynHBeD1ta4a
l7g/IBKtklO+1+XWLMtaBDDAx0TwXxcWREZOgo9roAfTYwmmx6KBOPUqxlkU1xj81OOJNrgXoqFn
hfeDwKuzb2eXzZoQKp7nlycRbI98O7miL+xiJUeTHUS/bNvgFTU3yMpyKjZ1JwW1a2qtS1u4Lw/D
ofor5mnIUIBZ/B8lQWZJsADBdZTuiFg7U3lbSS9hKBqtnOlfjxntp1FGaegavZcEeBEUsaNaLtzr
EHBlDcRW/7+xJjwDFnOSODmb0n84eGF6hOdoAnD9nuV8BvUWtGyS66WguK8OuNUqIrKHvbhOI8Ik
GlrfHPSAykGyGCVdphkE+eA1Nv2H/hXapzNWWv09aGqHlJtCAjQ6kHReDzBxGJGh5yHvt8qN2Sf1
OdpQkvR/eBxzauVXTEUYm30+gBRLYHLNvPjqHKlW2xWKBlVkBVvKbJHmOWtAYHDAh9bo1pdFD4H2
PRbFYBOSB9jfNfaf+TehfI4r/9hAFv0QFAJJKR8eIgTl5Pe2QZ10Sj7ltAwMkLzN9r21dOHC+c2s
hTu8bTd2BN1Ji8onBrZCjz3D+qVyTvxoN0JXwzMllJqtdUJeW39kBdVVxojg/yUKTPFUXVNsqK+E
P87y8iHgVxJaB/k2UqMRJ0OZti40rDHmWIj54rv8JP1Up+CUaNMfrKNFRSEkjW1GRiHWAZ6M6HMx
fOYRHY2hAAWYuVYv3ySs54XbSXUGGHgVsiU+t3lX0a5eCUzr4jJMXi4jBNwkNSQaV23mylckqHaZ
21b1tokKPzTA+giy3Qf957IVaeSZ/9KzGz7Gct52PPkwoLPAl/EQD5qSzEx/y1UYwAMagybJgEvb
NJvBZ0LaA7wwqIBEqyI8nJUZS6Xt6tp9DP9yzwU+JwYQBxEVm7pdYLlZmK9kfpERVMGdGWwdHH/0
AZTSJU2K2jQhvg8SXky5og4hhb0z78u2qlJ6WZSxyYQLYPLCBFQP6a3ETS4p8wc1xWmYyMnB8T3p
D5gbgfF28nPpu9o45yvdEnT3dGCZESSAY8h1//oj3OuRsr8UmXdKqLW3ESFoOlu7GZnG70LFf11W
D0heb+RzzBMvUITAezmp3yErMO7lyKR1CinPsY5OOMAmxibhtVSgd5bEAj3ClvorukfmsfXjflnl
VTLLfoKz2PgKK/qkPfJmoVBkZWtj98h4J9WOmvb15l+9zHE7g+hyHVqRSpxMAr+GUWpKqjov6kKK
E4BRNfzsgWovGWRCLjlPS/Rd4OtUrehOHe1uFm4/LUD6gBFF+Wmbdn7P7NHfkWu+AeQRPACUl14b
JiLFlwmvNWhdyd0nWMTdNUou7kN6piFlfkaVA2rA5Y1X7K/kZwVNGe3ySzX/1ehwQe+MrhaG+aqM
vYFm05eujJOU1uQMN4ZX69bilE2yYAha3+wEEZyh9wAJUSoi+B1di9DEnJFZdVmg2U5E433ZDFtU
XZWw5gTxo+EHKYhd/8To+Zh0ovLp+YvOxeXLTPYW3csPc2yFPfhnmHiH3x8gk/7wc2cGcZJneqKl
9U3TFeDf8uKtpn/trO7l3yfVUk4vPDIa0XdWAQzC8XdINT11udZcIXICICehvJBxbxyPidR6hUYs
2XFaIiU41mE+rpeiW4CF7ADxU7XOq//pPgW3Ino+YkAQFhaWZAz9uxGYgKkhGjehC/k6oa50bZUt
Ran2vY20mBj+tQ4ZYh/Vb8s/PBWzhCVrbqWNuWTj23GbDjHlpDQLRhGCic2DJgahy0lwTQUOVVKJ
WqzN8T+WfmoxCeersBPzpC75HGoFGjwvvamP3vQaTD8/eRyjNLwW4LEQPocmDrXVfoxZFws80wRA
Cdzc6rh5HEiA5sbmf7kyY4e2G+bYA1MdjOK4qfK4ohrd01qoXacYqUvrxOIVyNQWQ6Nq5pmT5psh
p9SQwupBIGYp01unlEE8/cAtI2zDF9Y1pKGKNLbmtaaNI33yBhC2Kc+jeHlVVcdiXNMNKzCHPM1r
irvGg9RexuqwwkYSALAbPwyAnGiZdWpkXFa4UVTQnv9uV34Ah+Gbkc+5g2J3mAvCJCLEBsy0VKUf
WDA2sZMgZDwRnZGmwqtriw5V7Ihr30kBdr/Mfo9NSWhJeAX+0nKhnZGU6uJ7uAxCAIJLupQdvrs6
UMSHdbCDWtuhInA03drcAyCKTVcHt3J9xjncJL07kach4D5UqbNxZvW3h//Tntt7hEadZ+ruhcYV
J6GZ4wMBPyWxF1y5ugZdg2XRI/UweFM3qonjiNAtUgTA63qtbAto5iG1/R2T7Cw5kASvmEGDb6/E
u3CHLeLm3KfmBidDFjUXfJ61DxgSpB1QqvEnZSHk9barNXG3fWxy+QeTKRAyy9zR/JLUhEbC25HF
7MycKDuFmAmzMm7BFFfavMgrSFhBwvJt+//Yeqs///AjuuxtB5xGTBn/KgCs0E+yzotPloj3q771
wgy/1qmsjLUrYiMSaj1v4TF7tMR1mMfxJv1JajyeIGuE15XaMDDgSEmtzFxBDlgtr/Z6E3Qn7D/Z
qxjXiSVkq6BYKuWuV1+qLIXGGcCQfO1ZovzEiV+DGVCKAQ2MKgrV4BANOOt7sMg2Yny2WA5R56jA
8sb3AzxTE6sqtsu5Rz40jqnG4LnJX4IC6ZJz/fpDhz4DCHZGK/qyMtDSRIydkKNG4Z4ib1gu/rvm
P/h+HraCQ4Y9j/tEqzYKSs3tEJtqsppI8PRrpJAZf6p8vkN1tJQSixV/51xnSSKhA/4Uqx+J8PBX
mmunMIxPp5IzF6822PN+/sjwT/t8Sj2rNSyKtNjK2qIzlqCHhoOk/ez2PeXlvELyOLSSdoXbBfUe
LrQCu4FLTfXVli3TFZTKvF6zYsWfg+vqcjqAWgxaGP7PtgwbJjTIBv+vFwCoJPVfPkj4x+aj6U62
Y9tLWQnbEHCQ/XH/RI5iPzP2Iu0yyBnQS5EMJEohUjHj9dDNYShJMJ1yc1Dbrb+qHA+6uv2/a5yS
n8m0THDaxbXHjB4cTkHBhj3SNPWWoBvrY+Frfm0HiPHGUa/k1XchlS8L/nhr+qEevWNv9ci8N4+d
R/JlmFUKHPMpOYlJTb6qKgAkXI0+cWmBMDXVz6k+2VNzVTGiwXiaQ/ztOLbwO0Mn0KIzKjD02Wcb
AaT6X/RZwivhX9Wf5wNvOREzVerHNlJo17vAri78OrJr2ZYfewkcrL+gEwlfRYl3GFcaoc9cdOLd
PSRjmPGa9oEziIEKI+zGqzLOnG3SmjdbGGhO1IZWloy+dCkfeSv1mvc7fecsL6Ftl9at40gEjCBe
7zANq9VUHHrqAvX6en/2YVe1qTEZUW1cOGuEeu4DfvuH31M/xOWb6GPe0vRLODYiJnWBWz+EdY0A
gwGZYyGdXvqyK1J1RZTUP//oGHbm9kawzVNr6+ifnQNqEYXdhhsMhL9Olx9d+aEKg77RAAaClZAw
w2GOqQo6Kepu3vp/CLPKadv28b8Vc3eKwDKX2DsRuuk5YPbld/y0H/yeQbkQyZcFL8td/ioVfIH2
0W7wE1kf8Si0og3T1RE9AYh6O7P0kyy8b0GLjlyXpAD1sw9PaTun7P0qiQzHiSgyOwf8TalmLnOK
S8MggL5bTvoyITXlqx8Y9M33gdI78OrTGG6u4+scDNwgZ/4kKnKb0IYcQBtujknwEM4Y2Euyq4MJ
mbzyLbBX+jgUSHE7KSVt9iLIdg/39Eu0Ij/r4m4Gct3n6Vqnqmn1QG7+OaZXCHxT5npWmoBuQ/1A
W6ewt6J6Aeo2x7MD7KvK+SX+VD7MlVffmGGTLl1DF6Qz4uBIgWoRQB7QtZzxHxyxkYp1y1go3LV4
Nvk29CO+oi2oTAs92pay7FfcNviNaWurjbkZJcUrFfpFu6o40hf5zXk72szxKA5FqhGy49c5bAe4
xAdga+t+mUQkoKhClefrEiiImAYPicnHtV7nIvsREBmTWBOT/jUtV/8mCk/fRcel+sZb8jHJFphs
7Vwmytl4ykC54vcVjOlXGApHjgVkyXYscOPvrqM20BWQjJgoLCFhUEayqeybbMNLDXi3exZX1bJO
B4I6eG/B6r1kcOC8XyQhldX2Y/CBcGEtnv1+xjG2kZAYiM21UB5PwWW3GZuHLHvhPRrexm1PXRQB
SaSaCEgpiPfs+FJmsrHUWCVDLtSOCotF/xf9a+ZH14o+OZ04bgtzkWtE2mkegHBwP13m1j2fmqeZ
QJt5xG1KbBBq/j8/eapVehFkrwXXJhbcfJURrHioLOFw7bwq8pDxIkYWEWKOkHiDHAIHHN/MYNsT
HYWF+MSb8EYKXXoeKxi/ZCovN3onUhGBRzeApkVJCv6a5Jj/L3qsPi0+advzc1O1xVZ0CQxIijVc
M9kHQgywbcB4a7NY8J5D0/cOeKMLQQDmkJtITB5RSOwonny4WBL4Aeme4Ke0EnENp6V3SIkK7ATM
slrFGHKCDFcJ+yIB2bpTCH4e47Ohp+HqfqgJNNXIF82l4uVcM2NRkzLGeHOg8lJvpEqLPgs0hG/g
B1gvMHgTR2xUZM67MjbZNFuUTY8Jzy5TWNT8AVzU3o3LR1+H1cuKuz83n+A2u4PvXjqoVg0wSAeb
znthG1FPgu+tr1TIbTbllt6qeWqNa9ZUa8tQwkVuqHkgv3uqREpj0Vqq5Gw2dUXVHJyN2ZBoOJ34
QApZDCC3PXwZNONGb15XlqUpaLCk6xYDffpESnguczPpAaVo3+7Hlt8xdbuwhbb4xEXyj7aJohgw
DFVdArgZE0BOpDfJFollqzVpxLyLcFgIQnQfnF3rtq0tlie3cmiHpEFWYj/XDoAwixcsFHocUrgx
CMSbp343eqsfKrjtpoln5ynamoafrqba0dvsS7hKGraX36ESDqvgm41BSY2+pfkG1ZTl3h/t7xP3
VyeAQgtb8wjjE63Mb5aYIiDJCko4KBZvC0jWdel3rWTy6uXlWlJN7uS2IromEuJn5VgA+rJY7aI1
NHii41Frc6ygmdCf0addM/hP+Rco5WaBxeHGqEyAhiYCIAoeI51qtuWbp/sVhHxg1zpig8N7xNVT
+apAXobkBHXmXiLw/WougzvPAgEkwY3O4TH8YUkcoHfprVHPzq5Z+M27KbCKWSh4bY1E7AEeRAnO
FctUZbItYyCuKykB9vDEtpiGAfLpo+xesJo/Kyfh9fFUSswvbdb2S5X9uDPHIy0wwtnTg4H9ZU/1
SRT5qk772qZJA4Sa0WfXSbPg7vwMetUE6cIsDM8Rq0yNO4N4JDRWNgemew0Y1Uj6nyoMOfi8SxDY
NY+byMffo4Usangt7qIS68IQ86Pf3ujKXz+3iRur96xQGybWBuixRvwqW/rBDKA3Hciw31f9VrS2
l6mqQ+4u7Ce/BMMV2Dob0lQjvEh0IcySc7HOcU8iV2IZSfLDQGzcMEiWMe3a/PM3NvD6MlGS9UTU
pYNH/qtxAuRv3k7WdPSJANUFGbBp8vG1lKRrjJydZIU3U36yMAleSYzpWTKUVzt/HsjDOAvAqyeF
o3gWakTEUfnqx5jrHMruglRhL65A88EayjrNBvCb0MVtI7ak7U1WOMvb8ne7suhiKMSeIscTxRab
h0QRWSbM4dnRqnrpyS/ud/FBp90fKy99rYoWftiYlRnoEZSLDnVV1I/LOcAmfr+4St/3pEpWzWFz
NQTdqdUKHct/YRvi7i+HdzcE4JlKXh+VzJe2IV42HcGrQ4zlPmGdaCNVr+3Qh/fdLVOMp5bG9NR2
CUd1IeF2YDwr6Y2PxYMXkctDDJvfFSHP6DH1OKk0hjWHR9FBTZgsY8TtGbR3sI0bte1IkxzlWlNn
Lom+aaTN19WhUNhP9Iv6w6/YejlYOKeGiL9KscwhMzO4sOFBiaLfhfFW7n1OiQ5Wxx48+tCEpedU
wQzmp9dhUDlW1QPfZuh6V6s3XLp7e3N3vRagoJeOEmvCiJQIrhKgkcAL+/ZNFSuDauIGy3liCeAH
si+RVucR/tIwnTMekyfytgNGgFuopFSj/kpVbxQIykTxABd0KU5Pol72vKvZK9n9fkE+APiiNYiz
3NnDV3NdWB6gtHQ+mAtwqvKoF497FbZzgncnm9LFV3u3JXWmWzsyf+ZKodqYZVyIuFOjeVYGFoD6
1PbFtA0acI9w6XDEN0CS8ubXUhTXn77dlvCR6oPgXwMFjz8JKS/fVS0v9pfA/U5TCM1IhRWbp8nL
coekoha51xJgd9lhUeLOX2mn8oyXz3xG/KbWCnCCr/f70G1jtMT0WIVKx4LABAqmAZYqucbxDoNr
7YdPkXHHKbnaLnOpBdp02NeJMIUyUjQz8TbNroj4kZfiSOv+derwfDq7cMqbjaiE+n6YK3A/8IZN
5ZvvmJbiElcjneb07kDWmRRYYk+2GQ5o+kgywC0ns2W36cz0guzSNzgwEWibSC4GYkzm8zHdYVoG
v3U9vD2BzRNjcylHjmmrxj1piMtN3LuGO6CHB4Rc66eUZRNF1XJ417fllq3+y3LEffsEvR+Iaf1W
KYDMMJFcgqBmLBasj6SzQJ2+u9oKeqwJqhGired7ZuI7ioj9SVeiVIAfNwhmIGj8Q+/XY1DGCUoN
dkBtQ7V0fy4k60d5WtxG1RagiTWV7CnBi4Nt58usRtoRupUd52SuO9xmvESLYzPABWLAaseWAFIo
Gum+DGdouoyE4nwH45yvm8UAmOPgWbBeL3bqnEjNQmvOztwM+GdSj4umlZWSePY+zJXOi64EJ1ol
grlEetwmFq3i5cjZFYg6/Y5fNLR9M4Df0LwdXhmkqCKe7mGGuf7L2W6YJr3EY6JX0tGFJezaNCqs
SU6bxMguNaes0bp8Re2G4aKWE9JKajLe9SMfmsrcybRvJ6+llssP8g4BTW/Gv8tlDIk7UWPq8fK2
UKqr4SJP+4ciRTay5dOnfobU/K1YP4LrV0qscLfdaGG+PPreCESXQ7eUgYiQxZsizGca0SZOYvO3
dbWijUhoJCMllH9XW672hMlLlFaSy+1T2+SN/HQBtRFPBTlcClQVl6mSPUzXZ7EoD+08f4apmfjr
GSyWSGIpo/jmZ8r9HWrhLfc+Zm6WEN64EIZr2mcJfMj21oJ4aBrefQRreC8vxdZfu9GSnk+LMGhd
DfEtnjea5ygrFhe4JR+vxnxdq2WV0oaGzIGanywIfXH1An8pD5tJHLps5fD92pugUGeYHlUoqvyx
Q4yyM+o1i1tl8yizFcsCiV1qLtCgtJHZDo4d6b0sRln8K/M/UuQFLJpNQ0FzXX5OKHfq5tYC1UC/
jUGoaRX6d9wDEs7AKgqbxhZzVR5ujL0RQaT9gUEl2e8p4OR1CMTWbg02ES8QoTYaB1UQA9tXfBgD
i7uDVdIXIFIDUfhc/QTZXEG63C2qyUec/s4nHUDMDgV+5o96VJP4wqQhPEc9AGvWlaQxKEPiscH5
46N1hv2QXcfFDR+AH9aXY2HwqdrhSoLpSh2TmjAa0J/DWXOxOOnGFKWsm/La7I7K3z4DLje3wNEo
/oqf3YPNzBJgDEqmlbDy7zzEqXERQj7Iep5jfuXxmvZgY7z9FHaPpgsAAmLB3Te+uHTvHLpoacI5
MEOtdkj6f0BGaLv+YkFiXX47akl61NZCCQ/epFME9qm7KQTJosO/ciSA6IFdNYBYYjkH+H1W4zZc
gU37EDr1R6Nz+qa834vdZCOWTOplkjgiRHVDo5/3ff3yIfBpiNz7+6HIf5kB0Zx57Z4z38GKgMdN
MFFbBkUz4TZRQ6DIYTosLdQ9SV0MrIcyld8MEG9hg6etPw2Y0QdslKoualK/1FYgCOkXXVKNzYfw
dFzZ6sm7zdRFKTbhxHQpk6FWWtE9NqDYupAMN9pQ7pVAhbP79EONA32E9cgHol1U9MbWTkh15Q24
dTngdRkzTewo7/+bfaXPUnBa9+b41qCnzIGz6wbSqgD9D9TVBRDDQHgMropDTIwgRgb58PfhWork
TSt2TsyPN8qE0+71TeyzLgJzdHjQEMgR2fjhq+EUT2wG8DVoOZYsDi79WbI4UvJVPiCmJPoMn4xV
GJEEd7acopYZqOKi/Vabr36aYjyjoC7+d/v+IwnG7ZYZq34GvhRvTA3pPlDJI+/m0rx1UhoriRSG
b4G5ddXkYQm1wqws2tSNOm6D+SKYLwyHp/StPsBKmFnuLBzGaIvhYZpsjDRxDUKY8WYBoVTJrYLY
USwrA/ePABQuYno6Pra2jNrZijAv8ZpIPBu+uNNnFV2ETiA++ocTvNFiTcC58+H6HB7gEKU7Jd0Q
MAhzkUtzlFVEHgu0Sf7IMvGG4FvJQG2y7Tp5gWCZ9T7cP+lip4pPHSgSmMPIlUk8LEN6XvENAd4k
yfdVIAca7+2S/+mIiOACql82hC+vPZCMQUDrb+1eUWn4XWUTyi5tye4GfMKhWIzJ7dyVM2bd+2+j
3UfXXPC/FfqrH4QK85jsBXb0Sl/Vj3ADLDPYXJXZ7XNNOC4CYYL7eBmIrC2lW6hFQdCoMU5rIrAo
G4Om3Ng6s1tiIFzsZM1+DxtKGYxIjCxrm8gcjoJed/3rbjN2wWBV/OoMQxcupCyzFetr1KFKJ/zT
NDyrGLv+c+UZIS5I5AecpADxmUR+DvdvXSfVuhVBwTu5vAaXe4y458dCczM18zZF405gLJX5DTrU
jG0O30t6N09wZwCc/jRhaq6s37gNqUnmwiNt1oVD8M11LbMdDQsVXd5l3eoOngUHKSnEOtY95IxG
H6N3ln3H0G9DQM3ZTz4w7rX3WN+QgkpxozegFMOpeM0g+1iqmNpI5hCE98tLFAhUSy+VzWCiLEqX
N2MviIlGLETv2dkalMVo+qxzlztFsS/eSAUjDoOMlaG1lid3BChtssBpdh3KcfWwXstlTvPguS2R
Dle887oPKAxKpwbbFscn8N0yCSC9wCmeTTCZLiMFPPsgi/HDAr+QMLeyWmQBkcKJXSP8X82T+igY
gFiJMKcC3Ct+3nt+isUPCB7TUCO3wzE0Gg9LT9m4zIxXui1XUnr4p3FDfpkEkMy8bSu+dF0FS70S
ZI3nsYz64XEMMVvmzFxFcVT4C8yOFa0s0GdS8hHESxTpq0OuMXeg7k4jo7/UOC7Lhtqt0JASIgin
6YAFKSxHqN//Dbz2L4pnsrdM2qhylC56YGYA2s1BnbUb6vTewVqBi75lO5atxmjVN8sp+h5XRPmW
VY38QpFnzuj63dV4iQvOrkuFSm0QCF09PUMy8FN7awsDUW1kmriZudelnUlCwaRzDuoGTdPPxl1W
qz8ZEHC/yzE/Xqyp/8DSuICIKZr4ww39dFWPHs1ulmNp1Rz+fZo4FkjgkajzZbv/Zr5xJ8czHSny
P6XjY4r/eX9Em59mdGGWF4Ud1fETGNFd6goVQXOC4SW6vIPyj9nC2p62jmSpiclC5URP6WaiJ7Vc
yyUHin+s4nCZlaPcd2t4V1kNVDFGixhQaiuH+H+tiRIsjnfIKTjzGqTwRX3sxgmtioGuihKHALRU
bR7r0FUW/8Fdyd1RqObyS71tfWZpwqqEHSScx2TRq7PGFh3N2R3X8stW88RVByiDTKyDkmidtT11
5dqZh/Z+F4R4tLnMIvZTnEidcSXOEzXGoXAsJIK0WfaxD4XLh0fqoDtezo5LZyzuiKdZnIye5teA
wZl+4qBVZaIHC+Dma6eP/gyQSfFBbx8/1xHO/DVIe+AdXf4h2v1CMXMN5x/9YKMm4hPUwKEptmzo
DHhM079Q0V07IuwlxIGOLGOy0s4ysXpfn9igHQlpc3kI9YgynyyKWl8rOWVGiKV1O6qlvSI5o19U
yYUZ1MTkydf3WeO6RSWiS4pfRUMJKSMuqpZqlCEZpyH8cQ7iETCvy+Uy5G2dzB+zkWnJLTpPHaP4
L9l9iDYPl+b2aArh2nAk7PBA2houvkeWnehscjbxlvyaXN8zC+FCVq1tlj/NwzUkpNf6FjqXFJot
BOaRILiO8tmmoHXjRrPATu0E2S7HsgjYdaUJnM/4MD9g5+4ePGM/OYt31SGyNF28fMa07jDyUjTZ
80LXxbgjfXvikWfXCb5h6UzxaUQbE2auEszJcR9RFhO/LYVQegy5nzht9M5BgTNwZOva7pgZc55J
BpsP0gBev8K4Sfx8s3gvT9b7uav7hhLR/nlf+BO1fL3n063X/ObenzY8PmDXK6qUPkEjvlmSfbLu
xWfFpO2U+vE0V4sNAm5LUjo++uqp7ry2FoD7O/n5/GirVklrrX/8SGuHL+yu5D3TlnPgyfjD0mAR
TlXQkdkoV9yXre/nYjRwCelQbX8tSxxJ2ApURDzgJgsW4D8awjNq+lO/Mnyvxb211aAzTTh6bE55
XdQdZnZ6sRe/Sk8haetO1uqstMPncnxUgLD7++D0vMYfg4L/pYew+iXH0R624/WMy6OXyvN33U+e
du9FFcp3L3QWMnNs9h0vPOmek16/93Wb+Ic4QlYlOB/Fqk9C1Wy45YJxz/mXPUB2NSdhnOX8iw1X
2qBr+tHxpP1fEQuJigrwyEaznStoi1EPwM/dAUZSFitGAqiMqpL5Lmufk5zMzYk6vSopFrshIlEy
zSfovbpHOVUoTJIdL4noNvCJI+riUnMEiXidlfszOBCuCrukeDXlCERoMpNidOtcM5Rl9r8VySjm
+1p5Bv69SK6Yp3ILPhBU4J2LC4uhiXwr2xLMb3P2IFj3cxXOHT+hMl1C4LDV5dH+3IN8UrCYOdA5
SFqxwO4HXtJquYXyg+dQ3yWJFNhA1TlHxzUTEqk5upMU0I2j28ZEnUHvcC7Pv0o87Mmro39mRATe
exUONOEIwiDkJ6Xs31pOb/JzfuinOX2xsPCSfC4InwSGUx0GG22q87t6P6/7/QclrpZ5ZrxXiQOY
3IZm9hMIWcjKwJFQ5JoFPLN94yK2EkcnizwRsZHKhkhlckQUOlU01m2aM6swO/mKKbtV1vDChp+C
mSrof/Lt4Qtm1SXIqg1DkwiP9oq8Rl3iFySTK2ai5bW5/FH4RAfIomTmVtgMcqyZOfuMMknuIEe/
7JutcZkb5wf/YVfY+Kohe/MR6Ld2fzHKRYOGsS7yVuiKB6eYUMdaS1TMxZ6vtvnB3J9iHM7bYFP0
heHNTjXIerGiYJSztNeVniHKygRZgfOd/Ee1g3j7kI9Zk6bnVjzXVnniNeWkeyoM9Sf6MV3G1JMk
DE66iZxI8Zj+YJftx8hFyPP2CCt65+fkjK0bRXkFDq5j1/0ul6t2FtJJivYNY6qtCxxKCsCOTvJn
eq9PH6jlpxv1QAlRFCpLTJt5dr9lcCFagb/ZvCqZFj9eJxhi9G2AwtVYSZR8BdcUjONgE74khnnx
HlFPGw7kPrP7WAXIAtv50A58zCe36NH63nYI3mc4GcVrSEUjl3bE2SNs2CP0ONAsqXxKROL3FDtV
8xA+XCu9rIRtPionhtbdNfpkmrwEr13BxFOrlvhytwLT1IzoU9B9v3v8ukhs01NtiFszCC++rUjV
WaOvDj3nOTXI/46VnXezWNAB4mCeNeZTP1vpwoc/ACBCU5Merz/HugeBd1IZFsIpwuNw8+6azFdX
fd4uJ3V3vx/jNlp444WArK0c6mRkoGetu0B9k5dQ7Q+/0dRFFSPkdwSsqlADmZEi6bXqaxtsvBVw
7beBVzC6QV055rPyDs+L4coItqPNPbx5oDYOa2GbhE01QrJtiHusz6Hi8ogcYnxDm6NKmEai3Q5E
FXalS5RRgwniC12zAgg2o/ZK5PWoYEnp9/J4rcSe6f7mHNTOEwilvbYdqZPlgoKNj1lkOm57KYgw
JHAIFYeYF6ZHwVbkM38iHVkhaDCPDn2Y91ID2eRusyMVlIqgGJ7XXzxipdl2qwnE84UlKMSPapZD
fTf4EzLqYkO7o/fyb5yxi3JJgDqSE3MllgdZT1vaOGKbPyJj8db4YRddlSgcuq8tlzmmxoMxIM7J
wawnoCVWdA2ozX8z1Cbia7ZR25HQ9v1R6Id1q56RZHd3xTDjbvl+EChILbrGfXKBI6h20yaW+NsX
W9qTa7TmfGfP2RwyKWkINZGg+a8YzGW2XS+f+HC9QHaK0vustEKM1gJ2UobmQ5YiCykhYgEO3yTw
5ALfzFveVlQvk9OoUGdg22H+bC5IHraj27FQT64E2PM4bxB+KFablsfxbqhnD8havlesG1dDfZkJ
ATSIPrjikVrxsbvQOVyF11P9c3l5inavfhxUauO+OTVOjgu7ibIswYhVcuDUTWbtwDFp3QsnfjOz
XlRSS6SJpOszPrWZRO96UgmtH4ZvYLZPrHBPOC224YTb1aM21uBz0I63rPYVVU3Tq2FYt2EyGU+n
M+WkI5ygU5sRKDi66PFMrxDkqR0MUC048mxTTHfvnxcVsskpuycoJa64gPBDPB9aLIBpCEmiqxGi
Ds9SsdzDs0Zk9KwnKe0k6iIAW4PA9Z/KrDHYyMCWJw4Fipc/fxVrR86jPDxHqqQFvUCY64xKdzuG
YZPYyf6x0SbjC4ZHeavqLiWCkK4MLqGwJmsM7XkWxJwqbpU+b1X9atZSO0anFjI4+NTt9QRBmiAT
OBm0tBCTqmNo+KDAHCa6z+rDaY7bU0zTLAoVgGtYm0eBBMMlpnBsFIUpQzJ6hPtUu5BZ6HRrgxf3
0h3ymYXot7hEms6IIDfM3Bl3veoTyUNX7jb7E8DpNJTEWWf3hqnj57/HGStwg1aQOHy2IsVn/zyp
SpM4zAE7cX0to3zJL5f/Uoj1qKqrPdchYnq9Ee8JOdJGcJC5bwXMZG8RW6TrWj+8xjanni7nJPy8
v/xOJAqu0s3PKJEvqdXIow2HIDGlxhxHWgtpcyT8baNNEp1fFy2HDqLIJTKqId2OoZsXrBVjkn65
dZKCbnEKdTdhRE54UhxdGHkr/OtN4oWSl6CuFYo0QA7DfmwoUjLzqCBElrGgDw8Geo5h7jfIUk/e
28zMrZ6Q/QMrXbIJ0V/ESB9zkrVfWUlGlTZqYCQpLxR74zBOv8uXHvLrO3DW38FSKNuruDpYL8mT
jJO0OghBXr2zwGQhFmRurTKMav7pU8UJ3vBnI/ZKPnoru9SFVkuARsTTALzOIVmgJDS7LAq0RWq9
MmcGZtJePEGTyYmDyH8fCtfRKv4N2vCc9832CSR/4A7xllKgHNXKu9r5ePX6Obx4dUcgJ+78a0sh
r7XMcEgEfnj7gfFefp9MNH0/htjH4H7RPHjO8dQ4jWUg6Xbq4aZoAmvo+S96bl7YmALqQV3XlIzd
CtuGjvRYlG0tFNs/o/FyjpTL+uavPD+Kw2rECcgni7oYR3BMk87xCWpEJN80ZHiUdjYqDD4Zq2E0
deJgEuS/AoWEKyHcuBX4v8XHBs+sSFTeeblqIkI/f/9HWZ5g7NwDcJQ2bLt+b2c03Ca8DK+0bi3m
75tvp3DMzHxgHXbSmQWWgYMu+4VOW/s73V8Kdb56dKG8muLVrAXv5/frvn8C/dP79AichWrY3ULL
jOC5/Hc1dtFp65pia6Ws+3BZJN0zXnSgRsK/a+qQCQWDXeQxYhE687wJpPKCQ02FQbOaUidp4bvs
fcnmYgQfq3J7LC8sk9W7jU0xmFSp8E7trM7JyjSLChE3yXIDZFb1LSurfE0TXxMxteVsUprZ4VBK
ZBofY2/C0Jr0P16cEV2xknvWEemTHmAJr9gI6lNkihy9u6adj7vs+P5dAqc5X0nDscLITENyPpC1
QNET+f4w4gZK+yrP5igBnw1XMIsT3mP2MBKclaxbmXa6t/axiL1m/GSlWsLICrWcG0cKOxK2Dn90
Vlf/9i7F/QBrT8genWsO90EyV9CNXr16/mfnMVbIAq5aGSc/oGXJSCIlSGJuYocAG7/fr5NqDnyZ
MLDJKmcODZuPICZKxC6QtHzRT6r3Hu2+cncKgcybRr6F+UL14VMO4V0z9fvL18ewcy3LMaRbmb9N
66zXEP59Ztv5Y5zI6I2r4Kh00jL1Cyuse6er4nvCruVRrZCgAVWxmDNZyGfnBGZCec2gc1qefK4g
BUhlm5Y9Y2fTHXm1zxNOzKeV9UbK+/LyA8eEfWEsKnCYFQndrP9+Bq6pfIqEzT4dUiobuvK6vyQr
sPRT60bQznABoYPDlXjGXZBRYaoJdexINAbH3NgsM12bb4brEY+QPBAoDs9Z/DdWfAf/sd5eTXAH
mvCS9s0NgjG+vZDOzXfolELLYl4WwFnNEQgZ11MSUItmU9WMcm5O0KLr/qE05IV1VmBh3i2SAIGh
tYpZpQk6sjXLKqrcmM0xDuALkT1VnRkatESGkt+VP2xKX+e9GrLmlG41mDxXytaw62RNDa4Sv2LY
rvFjEUYqp+TTNY+XAvYstrRWJlcxaFG9Kbqa6QDUwL+b8dIhb3JAEtjun/zk9NEs9Htc31AW4QdG
tvY8sy7KnW6SJuRuFZBf0+46TpLsfBT3yci0lPfI0zLduyLVkKUvmsm5cbjx+M2eLxudv4iOeBhO
pXdUlR/9ExZ04rvTHo5S+fk9RMdEW+JQIaS4LxG5q29+W9ZBl3uQTidQu0mlSevCefaQyo3SNVCm
QBLWWAPItbEHKRmvaWcRh2ttEO3UEEilUjNkWrj4tLVOZ9MlNbWSObNVxnPQRaE6iZElM/LFbn9o
G4XvywsZorYuvlvN41+Ss/UlHD15MADRwBeKWlXuQMftOHHXIfx5fkAPrVGxJfABLKECs9xdDrux
s7sp/IQOD5jOC+dA3HUlqmHayjIY3FKiFqaYJboIq7vhDWOgs4AwQnWgoRyCf5M2pH3w4PJadoRA
krpZgZ8xsLG0Z30I5jTXzrzMoqlsMVw4C1DvqvCDoKqiI4WvwUJ/iW22/wmMNSo4G8zl42ttUDOd
mVgxTWKAeIMZ9+PRhJuY6VOSi8vE0T9SZxZkrVDgW1B48MVgqEqpjvCeZkShcghHAJgp1hCo5GHV
d8rDj992GMorPy+nJD/XPbcL1yMGwoCZGIljpY/N0JUT8vy+jiQhGeGoj9vWupBoqPph2lmYiTxx
J/4SyNGUWIX2O0aOT5QdPTiEX1cZV4YRNcxMl5FID1PmJ3Rsy9+V0XYaQg6T//w3+VNxqK9i5ptC
JeFgkYv9cV4IykhfmNB4A8mOn1Cp2+evF63gCFWnqNOqFQN/fdvom6lBg3uyt0jrhp0ootCMuhZ7
BQzILGNWcDU6JKdhNrnUF11htRdCFOfjnQqM338Z5j/9j8WeVBg455B+3bDTy9VUNqUhbK993sAv
V/7C+M6kU3effG7Vl73ysqVt6pxIJlGw+ovoDEGA6HX2ZwaghmIcLyKeBAb+bmn9AfEYpw56b1Kz
BhfNAbdLNBYpcrZ6Hvztheg7qR0/7sTxVWo9ATOFWQM1kWsqXpAjcsWBFdDzdFVzGZEpJk4+O0Pe
hu+qtiIvAUupRm2RdIDMLtxogO/taZY4Csas3g0GY0Um5tHkB3T83B0lxkSX1rD3vQayHHb9JV6X
P/5SIsLk6xYh2E4Ske1keOYIpUkQFeEpony36Ww04UgQX3vJALyWRjIAft6q8kb+couMugVALJcP
JmUKWIqxsYpOnjXNs1muU1GfwNoTIp9f7PyJ/9H9kCjlCAOu4YmsmGiF55OxQ83zqafx484jXlOH
0JHhYRyE8s3yUfJpR1T7hnLhR1dAxLR33acx8dVjURSxDOqgh8byl5qp++90WU6ScW0veldGBmEB
ToFbBoqj5HsIbbakge300391udhvX6hQ4wboTZRqQggGMZqpcwcJKNoeLWxbjwnxtHgT6Eh2+kel
nBSI+TXW3111tlB5RVmrN0og5F045roLmwk3HFERyOKITrQAtB7h885PFCPoyyoEN7VF0cLLCjfW
+PTnxP4KVLBAQ+G48N22vklSZmdG519SjQcm+lZV/2DGHyMvtu5WCKLKO0hW/m+7/XNpiISA7kBM
e36ouNnjwmpV1cFyNUnRW3PeCsJhl6e8Kv8ohcKCXj7Oy0RJXDtOqSvxI9JmKsAtZSwNLXvH/y1L
G+BWbC8vZBkhNV3kaGJ4kV1RipYvcq9wjVcDTWjBL0NtegidHjeZHcXSDSXvB69KXxin1uq0gmGm
qzdZ77FOLPrD1U7hnciwofgvy98Rh8l2BJ9PCCTL5j9JOXW+WH19u31giFNz6GqsUNUktxNPdJkg
pwwgZQ1DFkyxlXASIL51lINHSalY3xuVNxxQII4JJPvr+bGWm5xgdsGL/Sn37SkA7qw1iKp3BTdh
SQ0XSC5mEsJU0mK2NjTxpPGJG4q8dMc/GcCo064zlLNsoaSFGq4BDFeIK45H1BOVp/aUPSp4176N
rHcSNTy8macr0wut3F9a9oLCWIjmEvNLDv/WN4mwuXqWMO6IbsLONTjPH5zfe9HE8U9o8FP3reb9
46uJUMC7mzjRNv/PVfPmFSY5VlSS6R+zswrS+Wib+D0Y8PfnPCoOcNu8niXzX+ivCSywpMPlOZ+m
hqmYn1UCGroBNydvT8tmo8gxiZJFURpv8AzgcnyQYtVD3suaDe/n1v7E1Ju5ZSysF+sjFGK1r4ne
zubf6oOH9sx5eNWHhyi/pvDbtZ4JRfGK3Epi4241+Q6BVj53jYGm5XeAWOoMbPExvE1zD+qv3keX
ACvCSD/fIRiht7YwYHth4sAq1Y0Ju4v/IsptXNYQEonlNUtNREsW+x2075amtkFtx3XhYtwkXOmo
XYNdDUNaU/pfj03vv6I/HEp2XlOdKgAcDudHDt8zgKVuO/qxA8KZZEkeA81kphjFI7qLDA9J5XjJ
fHaOH6ObC3rDFUpmPG1gddu8Ja+XxF53u+ikq9rHf6ZFTUP4wa/+2DOa+Y4ls6axlKyXC2W0r0Fi
IGvX8rczyvdgCJP+kPPm9U/FUl7FPM6HdTxa9MyrPJgyPq0rQ7MxdlD0MJMfIjHKlMTd5iYUlHBd
XGpwof5XkVRs6jUnMU4Hgalgw/aQkUllQvCu30yhtQyTOa9uxs48YraRlKPP+pdTZIGGat0ubrFO
SD+SGa4t4WW+sijU1fu2N6mAW4NnCAOK8vWxqFNQcvK6wnx7HOkyZJIbxcjVgcMaOsTO1C7a5FuM
EJHj4Z3YBQQ8vRrJeDJFF6k3c/ambm1yOiFJR4SGHQgOLUHv2RH7Z+Lt9/x382Gr457g0fkJvzHX
G+alxiNx1IzNnyCtck4wjKF6WlcFFXgFeHCgLbL0W3mwgHLYGBQnEAtZ0cZ7w53Z+G634lsg7C5I
oK0197g4hLSA7zkbgC8jKzRtlHxUs9TXgDFr5RwQHrYLGpWx833bNMkvO9JagtFDnRLUAg9DZ/xr
6iuQUvk3+dfaoAtjAP22fbh8vonOB4ChBpZQvK5YWkbC7zVDTJGgiCFkkS0nUA66y4b/9n4TGiDf
Okfv+Ianncm6YgwpsQk9nUmNzYYokDyYerBrHN6fS9vvC/mfzxeTCCEdT6wQgcoRH0MfAvCizFAb
1q2A3+MU6WVFee60aKvNN2KLc5HCrUtMZhyfsELaD3zCc4eewTYKKmoAs2gYHBMOmz8xj2lrohnJ
KYogZG+vNCGUD89U/ooi2BcTBkQWBnQ6vPl7wsBEi+H9XKys4o2Mqjez8nGD8UdB+QMNLDuX2/ts
TobEqCerwM9uFPo6eixgVfSa/vFpop12NzR48Kwp06y34o2cdZoyZCTv4eYLqxnQ2KBVJueSjTU4
FC6PW24SiAvZAz2+NbLljKg6w448xHnORIPJoOJubfjTxz1K0loyLnN/WoO3WzfOV009h3i6zdKO
vEQtZZbN7vka0dcv0F71+zQOdPERKaT+pBQ9Dzm6G6EqbmHdIjHC3BBISQwoo3mA5xOT4pWg287h
UsMwSn1Lq0BzRat/QA3447YOONBDUbHiAo0RH5QAFO9qD3wicIOmu7WkG3jiQdlSZYZwhEQzIdVW
waNakprAdByxISnyYNgdgdHyIiU19Ug3/pH1jXOQT7/GnEojiAediIx3hqdK6HClvEBLfod0d+uN
w0q2hQeoyzthMp2E4UlIRvjF+qjX6o8CGTOwC0Q5zN0AOg4GNPdFd+boa6xs9zQ5kPUA2u06cT1W
/JyfP23Moz8YbhAj+R7AmOveLqT4zi66+pCur145MYw41J99OXb5tppvi36aLpKzneI4xwoiDWzS
ItckznkPlIAGgco3wRZCGjNs74qxkZ4Tx6kn0I+08/RWSqf9Y89L6K1KPb/dqJhCFct9BOlCI2Ap
/Tot2TqplsSHFmVQ2pesr+5VcMq4Aj0FEGYWzQHwerOYu5kXNz6vDbIPYwldeOPQg9E1xxSEUszh
TEx2vlMs9pVDnx/qRerq+rGX2nErIZ32CZ5PVM/m0wqgS3VV6DQXhOe0z34thO60POoqRaqRgj+d
hjVBTAFB9bxrJhnyli5UufzoJyCaodol0sInkHTbNPoPS7isDVrXnkeD34pUuP0wAtLuXvu5yVg1
PDMdjclz5YBnK2NTvPyuVYWCseBwT3688zU8gIPAfoQI2Y5Za/n6HN4PKw04Ox7QDdDPgJATdAGc
JPVp7MZLVy0R7aZephDlcwfQwYkocewk6gVuA8p5mhvCaoO3frfMXUqjJPRi4IkIftZcnl62s0+h
PDDTbUfRvC5s2YzOV67Iftfr3dTAMiVh868eyFQW5+WeEebn8IVy46XGyWcfXOT618NkssIrgmM8
eO9bxJd2pZMZFNKkYRr3nxFufITGdIuulKC6zvktRS2MxiE9HRNhpoGUeAN9qlg3UElpootnu/um
S0xOvDwsE9vr6MoqdRiNqiW6+Cv3Cwdq36jWk+Pu+NDLPiz3ekz8uJ/DDhMHp4L0a0x5c/96zGPH
opSVbLRIJ9SB3biRykU+Wz3LPa9QmWnAWu4b+JTnANISQUkaJtCMGYzGH7J/7Ew0ibCsOCwW8qOv
zjkWZ8qjzSHo0+MmCytyP2DP4zhiYuTvwQnrc3ZI2d+fs2DpFZW3ohmuyXqrfNUWnyuvWDrnjlfM
7c2JrLgpFz/mD81eiFFFsE8OeWYtdagSjR2oWn03xxtA89wcjVUvrdFd0Jw6pQE5gCLNYbD+6abZ
ggp6vjQpqsrS1Qm3vD//MiCGOuyahubiR3rlJxN+HBvceiH4jgoDWiK9mf0K69FevWCtXSyVGdJO
zqMNQ+pv64r3PWY/ieXeewMyTuJIynykXtuG/wfklS/oTOY95rHDPkls806fWTRxqWDzDC9SqLlP
++Now7pxwYQDULDKlkxpNNfiDBayv40NIK9S6zHyBC61By2mh+m5RGVJh3PWWRxrRShgjcvd/tx1
Pv1yIpHKOEpAWG8tOrWziU4ufeH3vUby2e487OA5UucVAUO2Mf4zFABfPcxF5WVSl3ok/0H16IQc
68rD/3xa/xWxXWnsRX5EOKzpfzh0T3DA8q9xeb06WFUkHaTcp18x7BBaFaPufqcxft8ysnCXz5Ak
KIdxCvh891lssuuj65MTeQgCXoCpgy7eHgXz5nAXvKB8s0Kj+2xluv0MrSKGM8ughmzoA1Nw6R27
Lp+7n5hVPRnWmPEBoNLLZKWzcmYcU3w0xLtDI0p96frHfPJe5UMsyaYTDokSw2piRocFQ6Llyq/V
05jKYR5dk8lpjd8MD6vA+WmbJmKl+6hp09IpjNnBaTM4YXLzc8kNzimXQcIDTpV39RADtZGpb/aI
T56JtqPhlZZXF4+/nIxnrd9/67DkDzlsk9RWFhugruopQKqc9JXb11G3BsVpZsTqUZdqluhCOWnY
HIhqFnAtIFN1YWVDHAKlUF3IbWWZitejBE5jH43Dcsi+TuQoUhv5KcbtPITjVD5QTz8xUGLWGiUo
vCvytEkGh1RdzIhKpmd/Tbyo45SREOqsuAV5UDATKMhalCOjgmJcw9c+H9I2opoc9hlmhBh4HWA3
C4AKSxMRT0/whiDujbiIAtEQmZ8M3ovPgK0am6NIvXmQjRWaE/Pki40/cAfFVy+2odj21aZsE6k5
qoWeL/HvY9JGBHwsFCUhSnNtFGFOmjskFE35TUALgPUHA7vqDr49LHOEZKlSoRlrL0nju1B9FiaE
cYbR60GN+LNZu3uDkdj/LoMmLst1+b/Jc9+BxP6jiNbdnomHuI9+y4OsA4voPQo7e9kaoQydRHDv
sMsLie0K6gGSrwI5V4oNQRN1NOeuBegLghgomIdEWFB4s1t0ur7BLFvX4qLjEsASq3f2YY4QvhCl
TzvYn7NPZCcRHnLzRhubp6T+yux4UqOo6n1MTUPmypib0DAduXrx3L9YmJkmb4CeoamTqztMUHG9
n5FrwDPewEUeDf+77UWN5UxSaUN6Lhz1mraXuV1M4lDp4+3sBY/rai1sIFDaNZ+Wx12097+5rtKK
1r2dE5kSewN5vTGvdeVNQkM/W2Fq+HRLBBUhPcawx3uIuzSTg5YrKvNz2n6Xw1kd0p3ax8QvXLTq
LEayzdB4GyMCEH5HUFuDAvkSwkDBetWPsz5nsgX5NC85Mwg1ffp6e+NcWKpDWRvfid+HB4erZ2NA
TutePTZm/9BQjRlsYwgh5NafB7HHFwVAu6PrmtbU+Kb/xnvWVx/VZwmwdFTMBIhbdP935ZKZpgmD
cRY7XyXZf5r7oQ9I14vqN7AN8bbBOusXVCM7N4hNQ+GiXl52ZgjMS945hK5fkzyN5sNYD4mdnd9h
YSWAPAQKe6V7LuEGqfFcOuB4ZucdjQJxz1J2OVOIWChATFtQThrbL2v5JAVtl1WEZZG9b44Zfbbs
+LkDzReKnGde++CoHZxALaRXGB9wiWTnt3Lgw/gkH+1RGI4K01c7h18AH2z34ovHTyf92+RB4jWg
9Sn2pPwcfXtM+YOjb7d1Hgdz8IiSLJcUI00YYHxnamI0ysCnfJsHijJZF98w3q4e0EmF7+hdUj63
W30HFfnr+66zO5cmWMLdwJlu+/VB4m+AosppDLh7yxbv00rc3h+mnvAHroy1DRYI5o9BRcs8+MSd
85e6xhekB2C3YDBkZ3Uh2nJF1VSl856BWIy2Wj3NBC6X9qZscr3g4FH0THw7c03nd3zwLnsHlq0j
x3XPFsO3BzmkOB713njWnKLA/cKIn4yqVgNFwkuxjL/aLR3hWuYbDv8GKB097sAZuCcIj04lJLe8
i6zpiyEatlkZy1RBmirqv0xJtrFQgVkImpGS2BXgn1N7zfsYWRLqEaMgV5x7qqhUXu3Qxa3HJUb4
JUbKRrxpUdsfr04QI2umUQqZUKT/ef4gh2VuyLlLLwIUYAbtkadR5DGvPrD1rNI3cIZl1HqxNhMA
PYi+rq60Tlo0aWeOITx5sNA1p5hlD4oOrR3I8BcvyABd7oJsHYWeJyAWtu0THDf7FUz3Ek3wcfBX
5RzfQ1Eli/5jwt7EOb1o/EMvdfI7yE0dOjmKlH/yT8e8tXw8sU3fuROcGm89/AHI/m+Mf/brV3p1
mhmbUaU60fc1j1HrLE/++9vaxhVePANQNsl5AFBxQ/c6gH0BtwAkCxVffd2qOvVKI62hb8OP8BzA
l8QRQUn066DuB0oJlgTHgoMmbKaxbKlNtQO3EFjr8sUxiOgz2vxcuVhiTyueXUDTpS0W9F991x/B
8uCPbRY+4quCyDZtoxA4Cgc2xTNYmsE/vIqhR3rtsf5mxHVOF1ZwpfbAAK7U/xjvcTW53bqu4yTt
QsMqlyJBstuZY+lSqYmBjEglUsblrI/XNo0S/cPRmTzyYAL80w8wx3/XMobbmXwMRtJ8uPAQYezq
NGnjQqEjSKiZUtJdRoS0bwVJLyGiZozH8WL1yGnTOUBNrzcakna8v3DW47rQw0s+3RbrrrRVWa1a
+VGYdBr9cYm/HKV30SxOh7b4anN93nFMd8JP5FW4zBPedxj9g/kk+YDIipr4wCOfKG/cvFqdvxLS
ZTDHnqMFCWbjAn2Z2L+a+4Pw3f+oNkNpy/J6+sYMkOt1gJaeGAo4hnSEXA+IXCP2+KQ49lOmkFF2
4hk+4RjeKDH7/MWgeDgN9EWbcgag7eNxcDQDNZF9Rg8K58vukYUTZWCgDErDhVTqGXM0lsuLSrMP
66Nf2gfER8t+lMdVTi5uY5gLheJpbJPDYX/BswTJQqRHXTAX0rhwKrmQMwK7yuPy/WfSnFx+pJgm
QYYAVSNJXiNhoTxDnrpiqhBdbA9pbHn/wLdwNgG8mDAHGYxQ5TKW4I0D8Qm6C0M66md2NVVkPJAN
QfFK6gVp/behQLDjsdqfwBvD1E4sJQdflSyi9GgEIYUnwZJOWzuCiL7r5uG23PMRy7PcYve4Ccew
FrmTejpohTUFKYuvYuJMya1moAQBisb323P+oXhbDl4tgUrZW8yMzTCdiZVNYLfCK2DAvTM7/gfe
JgHJCoyGVgO7RNNeZwADDOh9M3ltv18eDT0kcS5k8k0LYUuxd4PZmMJFe4MCS5dAjf8sEZkvv4QL
NIHMNg+tB5oEdAdR40EAK2ez5k2nCQlDquF9UN3SFCfSwyUWVF1yDzPPFJqcOHZvReRjMgTrVF21
rJFIm9YKHumPfglMdn8pEwe1AMdxraFRWw/Nu3C2ai9NTC96zE+UAf1VY6IteukRR0gtKL3TS9Yz
LMkHR+HOePZq2eRpfmYMyIuCAS8M39eAOe1i5X7gXkkJKVJ41ePbBYJejeXnBhzkZ05efjtePkpf
h+X18ZJz5A+k7MqhxqIBD7IrLyURCYPbOB6JVudooJ+pDYwHNJiooEwHhVV+4+j5icxXIG2Luicf
cmea4wK2Ioi6IDfwMhoVKmquy/GuRQF9DHP8Mt9L8CeEFHPmF8XCNUEnfP8C/+Q5ePPZMtD+mwMr
mWBwaPaYqTtYWstr8mfTTAifiDxhdLqamBRPNeVHNL8dJPqAqKAR8yHIC/GrD5BUkYlLuhVYeX1H
zwH5cPWK+QRtmwQjlrH2+qKU4fUpNvKwWkR2voQvYmGNWQamhZN2rnRqpWcXGQfec2ykIdaVPVaf
nlcBFG8Cv2caBdQguOnaW+9ez/6oFhntmO2+oC+yG1D77ujxU9YltZDoLzgLW2FNeU3qefKkhp1U
1EPLil5KZBM6OQwfg92Sf8HaNugfpoR5tMMNsIjRyfe9BNuPNGJrG3q0OYBr46Nt3TEsJbE4VVWx
PnCZO+6NiUqNFXDeJglvP8QQwLhg/Gc21KV2vs1i9E4OVRNTxNqi6dUZp+MQ1u4UqiSHEfjzoGTZ
jCn/G6No9eTgfHsWX2i1wD6J3kJDRdp9P+hMzQDVQ1XBGd/gmYRv2tZ+2lLLsDca/PCmLpIcG6Nj
fM8pdysqKuMweWXngofgrjg+pWFDj6/AtUk+UXlC5D3k0VKrr+LWniJ2LW5f/CQJoyXEbvQzjSdl
70pw8xJgWOK9Qd0ADTFuvfi5DLUWn9b1VaEaibP4ri43Ns2IIT1baZ0Pvbdj/0NM9K4CZqt2Kq09
PCLzhoF8bkQWH9TXBE/No0SxX83wSdENW5rrGoy9XDGT+JYbJ7n6kGJywhRFVMPa/CW4GgUQR1fC
2BoGN3/sIgW9zKNEyJUsTIY59cXCdFDBdVYvOg5B0sA83H7tXGwHYZ68L46oFK1RP5+GK3SkTr9J
yCp8yCHLklSfIG4z8FdfyHOVeHXnf8bzLBoRZpQd8et7BdrC6RMa/FNbJX35TvqvtfqZMIYyJt04
1ibHKHUKf6JAnjJyF8x7lhqtdYP1bQ3Yotk3KJ22cauWfAxFKqklqhQc5Of+SjNQrDLnCVvJdEL7
DdCUTAlh2InfwhoCVF04o0fE52r3EAV2olCrqTckaogs1DNi4R//MYkXKSeHZd+u5A1V33dhLE1S
NTjIYv1xychKf52ukFqElOJEKKlf2wSzlT5AneZk/SHdLvY/POgQyKsNeNp12dh6lblQKqmfmfJo
tLBqZBNIpMOCJpXmrY8e0Sjkk9TP9UAuT/tgfRigBdF4BJqOmbwMGVvi71IZzBkEHMjQAnXI25qW
7BVfhav9aO7yQTgi8d5BFDnx3dteQe+BRisF+GjUeN2HK1JBNUYERhnt6WElpiGGFy4UlrohirMF
GH4NtuT556icgjjWnkj0wz5cBBq5x4RIes0AgbO/LJmshkY1nH8Bwe1nkSs7LKbpeNv2gjjrd3oM
ZqHRzsFywtBbGwiNvTWmvQrUOFipRIWYgzg8slE2zXACQTGM4BdLXeTCglNTFDkzUMJqZb4UHoIi
kECX77oI+nojkayTffC4bccMO6xp+5dzLQQVkvK/goL9bnKZzxSye7s5iobqmBimlakliOw6W1Du
n8+6dvfXo694sY/M4IrIZV9yzl/9LZdj9TrDo9/S+qgnYy3YdZCmNfp/32xSfztjp25ZZpw5ibbH
5S/6wqW+SY3zs/YHuJbvnTMjzzX47SlcehO+Jc/NWidZ7OFha6Zg7LDENQ7fBxSPxi+dMmddmbKd
vCpZ75brvVzvLsOo7OKcsrHziCnb8s6YrA3UfZbcrh07cBtH7GNlWg2T2rUnvjYgZN3WhNJ5fo2p
u42kD5IOTiTNODxfJkRJ1xZ5wyfHd/V92yOvDC51Jo2hw3SGESHejVjW9ronUeYwfrdkwiBVkxIi
7L3w103teHI6GY1b3vGxFViGVsei5Ff10J+muR0rzbli7UdmE3yauekN/Nd3D4X0tOGExa4q3XoP
EBcIOV0xyFZpMJulYu9wFw0PN9pR4ZMV3RyGOloihYXuNo7rJG8WTLS3NRAbbjh/0onRgj+jhIOC
T7gFYoFvSV/FRM0SjwDrdyqq3F99gzDf95AhrU6fp5AGNoHlCEEwOKk32YqjzaeJfrg66KfAcah/
gdpAD8HpGEZaCXUietzLTLnx4g21CXMFg89/R49x4zViUOlDabZ99mnaP+bw6JDUL6uS/E4Jyi8s
osp4LlkQDHcq8t5KSq+jcyh8HkPVgmjDDNAoEfL5IeoB80ZVQdMSuXvtJnJiZU5WZXsAiZ5TqCXn
9uigUPk2QlmOrHuHsAM2oyD8YW3RhuIqP/fIk3k1EXksSUlg0HA0BjqTnoBfHr59XtDxzy8DMygt
jdhkCoxqRZ8Kv1AEpqfUIHNGek/o0DD4Yg6TKjGRHoapGv5UvQpaQ8tZ61XqZNfF60qAM7avjiUS
FPOxIE08W3MJaSFNoRjUZssrzBWu9DlVn6PEoPijAsXk42+HmFdWhRm6xkuM7TC8vcYaeXAnDRCC
oU6+dUDSmnnB0hixS6/NliALQsU6XEWNFV766RxMnpyW44bfiH81Ue5tE90eB3OtPDxd0pPFKg+v
jc3VGwNIm1W9ii/ilGJN0znxVMy0A9m64ewS/iCUozB1cC6IvYBFNHgazuwHBIK77sLZIU+wxN9M
HL/yJRSHQr/UeZsT5OZXY0g6jMZwJvjb+8vPx/2AZP/WMddhH4PF2QpkzqDJWkhrEgDUTk0hhPCn
2FkWPalGUD3g/mtbFsPBR7b8/Ze3ZO/s8V82TLnBoJ04yNYHWEReyoWHDkwc5eMtIfa5Ic5rzYxZ
63DB04xfccxrJCS8pEPqvjGngjzE2q/V3Bs9CI698w/d5I7FDEDNr4UM7Jh4I4QBovmVZA0xyNjS
LIWb3HE0nCHgODN4r/96z2ZyYmeSAlGqm0rgiaUkdlzaVEv5cUXrrC+IsLARWV4ZoC6AwWpJgzEj
kLT48ShOIm60AodQwZpLd3KMcEsLi6LsXhGm3tkkXhO2KSH4x4t4jSacfY8YCHfoeCthPyExJiYO
qdHXM0ivyzwxmyUuPaF3LoVzyfrIsoBPhO5+X8Nd3X0JfME1fLSSj2J41y71DpS8A5qHY/jhqlR3
g95fQsqSutTH21siCHw3C0AeR/dPm5FabCkbVsRJuwa1TOb0QpgwnSMmiD9ZREg1ogPhXpyfb5NS
wtKCIZvOvA57pstcQPhEn8YbI/dytk3CWSJGUwq3HzOmW2WkJccFerJN16RJQYhq2odKvVTpNUAE
w8vdxeGMgEQdaOTRle0vE/RdbjB7zt4PF12RN5p4MTZvFEujTcYXrD93/MGfoIcZzCpTdZ7p7K/P
Vsue/JdfO56QI5jO0GB6lniHUjdqnc92BirVMaOUXwYtpmcOis+xMX6EY0wiXE6NKzk59m6bcqN/
d6LH9w255+5/0fhvv9RhQrmgoX7kIjCFC4pZz3HABA1a7OnkKwYFG2J0FIlIfmpk2M5yf/OlpB3v
0aefBGG23WvIgkybCja+4Bf3BTzNvVmHeSmhDbPVJb/ocfKayAu2d6dzxOGSWcsGAs2Z7NgcWK0U
z/kC9GPiwBznYmTtPNFJBfe0Esg2yFV9N6HRLHQjYw+YsvUL9NvmkwgYiTV4EwZEzPgcAGIpXfZC
1rniL6u1/HWK97+mnJmRd7gNCK28pTqhIumP076Pof0Rmc/ndlaAOLqj8Yi0EEjYXnCglMhYSUhm
blXwc+hfP/8tyBZrSM9anbOrSZnqM/WdWCGzytT58rSu5JTuMwzjHb5ygZkL/Qhzp2vqE3YBGP3y
COW8PPw8kLab1BX7onzAieIx+MIF00YEDPf38S7saZ15NNAfICADiRnwn4hhwriQoySmkOghD8uN
sFdbnwocbxZhjFOR2T34nLrCl/cMznbl6fxut6ZJRlP33ijOadODhcbNuPmdRglXFaUL6OY6KI6t
C1PXD9nOPI4vQ77sQ2JrI4BWK1GBbd/Elj8BOyJLYflyePNY8woqQcnk62l7pqFPb0m4I1yqEl8I
hwAPsF2nWrsWjPLdFtG8eThyAGRVngK1gkcwVfzXSHVKPoDfx8gQMXtg1USOapwWkbTAUnKib7JT
K72pIaNkewFGHFhU8ht4Z0e4xKSI2MbvPn5/KfgjaUrJGdmCSeWrx7/ikm3O4FsT82CdHPA8hIxJ
+zJbC0fi1sJ5DYgl+nnUi3SniYIxkmaM+OY+RweNe7/fhaRo00CkFs86+IDQzsnFUMsHbRHAz8Iz
z8gyroSpUYqCVo4di1Uo7GG6HNbVGDDxr8UbDyLGtXDbpEUegz7625UDE9AUMzAzvWydXwGDjgzx
mq7M6Yj+EnLGeSVioGqTWGzOBE7pOhf8P2r0+J5lFwh24A+QiJa29on/8H7LRdYxFWG2sEEgyTfL
swAvEnuezZWZlvUFd32rUZnVkV9vR9hHcGf/HzP4viHWYnJ28mljQaMMsuSd/EqGddgHznpoV6e8
wclgnNb2a/uQAVoZhydT1HzxCVDZiUFWGiGLNZK9846eiP0Wacfkrpt9O7S2/ah9E8QN7xEWIakh
pa31MkWX/EdyDQjChIiMi9FzliUH7RwewzMeu2UY8cmb7X8GWYQN+V3cDgvvoOA/hsXtIpr8g+2j
xJBb9iPo02mdEOPkON9CFq0dbVaWk7KB6jVPcp4ZU5vrK4EJbPfoMpMWq4idjfh/9xmeihGZln9N
K1QvQyVicI+vQHyiNIgZP1gKL43EuhcoUFnFZgFl3BJlyX/XjDJ80ti+jDjrvjRA4SAlx+YVzk4s
eZu5ajeJSdFSSPYv2YnsnFVHk+OcPE9PEcYQp8IVWG5HI+5J/EYo+VphvWCKRlZt1hkpgfxvFzgl
uP/6+LgLLkatpVrxfo8iHH/Ppyot/F8r4iIFtbkfz1iUR4pqc7e5TQOvfoy2JPVdllU+UHC3ICw1
EOJJR9V/kCnn9rpa1H7dmZh+szj4qBnVwW3e09L1J38mk3/Jew1BbDdB3a5ABto+hG4LV4e4La9n
Ybd7PuLUYR3VxW8gn592Nu7kOA5xW20OZ3ksa3ocD5Pg808stpP2Cnz8uBvYL4ruCFOgqcT8Mikp
4QGPlpfIRbXzq3twFe0bUVsSTxrI1oOlfD6cWtGjxqnqpqLxNDtJ1ktu1BoWkV9WfmB4nI8IJEm6
5074heYRacFos1l8NAE+gP4gV+EKLH368QhPnOrUyYJhw7hHiY/gTsf9RU+QpFDMq70bmEnFBsTs
dkZcRV0GhjoYArZ7uUQIpKweUmW5bceZiOjLKbU4UbXGd7w+yE7CauQ8VEbMPvmk1ANBVUqqakYm
dy8mphdgU8HBWNF8XEGmsCKamhLuPGes+bOJWC//c5jwMiE40FjPQ4XiMfEWwQhY8tvhZO5jJDPI
/oadjcTAPZpB819MJjmHDznHx80Z6iiABDRx+4ZQz0hiwn7Y0yeh2do8KLA5zbzzOAv1kBiC3gGY
R02mMGEu2AToX86ACTI03DclLOpbAau5Lgb/Jr2VS2pHW1taYxMp3Ax7YSZeuqsT/v/WhjHCR6q2
24U9ehIDaAadQTAen2Er/hMcKat57tLJu1t4eEwfPD2KQSM2b9WN/BNlijW5F34Bu1gbXeO9obDr
YwFAN8wJSPNM6L3TvhgNRXUeYFfCUeliwsA9+UbLTXy3n+XS8uu0T5Oa+mwWRBJ87T0DgDbwXF3V
KEnh+FrcAmyv8wJdT6uvyUtX0RTvvsp5iXpMkisDccF/YV3xE2sK5Sdh8qg5CY7pSCjH1hehOtGa
ByF+7rJqHtmCQBTNIHQ2oMxLKBKieYFpBknEvhW5KWx3pmu5kgwKz/2btdUPNpyDSVlMlHZEMT6/
lPPiSI1uGG8//wsWeICNCEDe9lbFd2TXuxU+KgdS2ibLtZbyxA2x847TqLve2UAAnLj1FY7Fq7pU
psA+/8VJkkAU6KupUzBBpAaEY8SyXRX8P2oJY22+t/HWUyuXsTK/3V06Cpke4iyPVUEYVeOmBvBJ
mbRPpwGr4kULfN4hvSM6NG4DoKtN25TxuKnjMfwzL49wEDXHvi/qMQtZNr+6aLyJB7tHU7pnwv/b
RBk0oWiAQud3fB/6t6I4dMFZB/kt2SE9eUD6a6PLqYfnAfG7nlmTnHlkVq5Io6OR+y8PA4tnNU73
TksnRLKZoKlKAoCfiXiRHC0txupw0D//JvuakMcOT2u5/+0RMM8g3vUO4DKEDxrmgS4HQ7QxHf1r
ysJAyESHBqLMdVSxxUCISyzjNXPFAWGGa9CwH0ZktNJYpAIcf7r5fz2CqEs9yefjJvHiZVnuNmHR
qP3K7AQ49ilXGIde9BNbIGqYDocUIfzTIzw4n3mviGdCcN4vgwX/5EQrw3yrRAf156IU5/EKDVnT
0x8iRihQSSagwIeq2el8LIqFoIPLMpvseGUWHcdRclJpkT+tEPKmvmpkI/au8Q+s/xt8pb2l63+6
EZ0IsnbEEeU7iBIw98YFRdlrRXQIDGfos6CstIszgCFfVqQmWr+NZXeeUYJBkCT2L1IYufmwEFwo
pWRMMtktdZ3rbb8tmNe3wxx1Ue22Vdh38Fan+6Ff4sMsmn/6/GLK3YF58nXGG9yLLLU1chPafN3g
LEfYg5cS1LngYOSkAfjK6bZojng+fYgrVVGiuNvaCbV7reDJ4Twnr5MZgpd0Qf9meU0wXWf9yi2O
zAOuDOmpRDnta2bZBNCpe2noEyd7mD7bf6NLTXw0KHjG3OJx7TILG1Lmg0QKI3o/TAIyskMwaLig
VGZFp3DIJ3cvkFCSgSPJh2jzQLDYVH6svWZSvVA9cnOONFt3cezt/6jT+BJyu4OdToEuhIUhkc82
a7TQbrYCV0O5FH9RQRgLIioKeqY06vlnK/xYYGHLF/E2rcrd/nWL83K3bhDUBiY2PwTOKezzFHX2
VLgg+OKTDZp9ac5dYtz4iOIDuqmnHIJK2nybUNqTCS9iK4EvBrpsCLlaPGolKDz3hMqr6qH9ll21
NYoDqZAlRol/V1AMQd3h8C7gu05PI/I81ob1qZqkJW7Nm4Vagw8RjgW7Ui9x1UXBUeKsuv4JYEub
vmoB6z7oy1H3ztRyOhSs68OMkhnCBRrZrqZlkK0p3LkjRO1IboJzb3zXuNKJn80/xuzKm2bNvPuD
eExTdIeiuRzXypdZbLoCOhKIc/yV/KXKqx6+bw6XXRN83bPOFlffLMlsVLjQxPzww/HQ2OS96c68
6Ude6GaKAqCKzx70m3mkpYVwkio6Z4l2WGfSasFAbDQzSx2RpiDwpxiqS4pfhUi43p8/0GWbJKwK
wkBjVVPOfmF0lsQ9TPky4UulmaFr4AZp4rTJ9nsINNqFbfHcSNJkfXvnbm6/N/jZGxOgJZ/99jAW
cH8jlTo8/+elR5CFaAza7VKaf1N6Ux3LKKIx0Jd3czgJpzh27kes0PXZpY7QiJoQHHKt/ORw+l5X
f1elJDNBYSel6Pe/4XxugwotCSWs9fFvb+H9YLHIhY49M5luL4AP3exN23GXOuuwMzaBFkaPf6b8
5XaGrlSe3scQFvoMr/idwwWBJeR5TvCBvDnj5/txeHce87TKvLUst7xbPKjaBbyBTJyF5xotR74T
ZRMneI1lXegFbGQXpfdR9AZk1+2X28rDUlxDEmxOXneKbfljV+xfmTyG9SErDoKP9luPkwA7as4D
TkDb0vBSytPit4Kf11u/5bmtwVdkB6hspV8kjD1TEJdXEXBcfolOvriq1qo616aUo0e399GO8sad
zE3bq2FQUk9XOPMH6Zflu0l/Iq9S4TmQ0ewMqlHyfU1iYU5YIE3oaXkNPFeh8iFi0vcSWYtSJJIy
KvG6bApEZXunQYmNx4fXv/AFk8l0lrZXnuTc7HqdcUk7hgXaGXRUQ0zxKPX5sUsHQAJVUK7ttn+s
4qpqLAEzqVnrDLLWxH0Y33HWtPQDUnm7G9QpKIQSvT1pfbc+BxThk2FGRzAGIiVjoJmDbGDebYXJ
X1HLHOdkGjz69pIarp2+85HcyVMkkDxNUpHc6cbm45MZxTPBzSdRK4EWpKVEDhZecVko49hl88d/
eEgLyT76OrONGRfAzAjgB93O3sg2JL2wkRkjNSA2SbKXOfYGzJq0vcyqTuTXcqA16HeVpSo7fhPt
AAE2AkY846i8WBq+rDgi4izBjyc2NQz5Qox4sKCVObpLf+JnBrTkPl/X403ttEhTzkwDOwXC1xSX
cLXwXOAkqfpu5dTlxyTYigCISE2/qqVolQqeFWbFQ3405FjNem0NHtRRpaVrnok2wbTVr2U9lpSZ
9tTlBPXbKnJljedC8yK+mqeTHtP5O7LzFZ/FMwJbNNefXQ1/ec3X3JIsioFY2mfLzklgVbIjD2Lz
s7N4vJMOaWMrrEnYpA9KtAILfU2PMRHTm/72I0sKvd7pSFiy2op9B/LC/Vpz46tAaYzun2ncL+Sc
Ft8QbzFs7bbQER34rYDtqK168N7mSd0wVzX8/Xuk/1RWwOA9mBwge7KQK2ZeVeagXzc6Yz1r8MRA
TfD84/fkZziafIQiiJWYYaYrdTbgVCMr+YPITKHto78A6I7ietzUqdHKWtleV2v0eMgcwrvFCJPd
/hc+HnXSMs5nMJvQL0yeZU/56iK6iN10H+kXvtu3l9olZHVIqv/+1hJPf5yfTh7ynCVQXx25eCib
bW/FWP3Lm3r66H2mXnpTeRkh0YzM3WSXxu0Z3W15TOYKDCcVBJzGQF/90WbaNHXmE3446Ns3u+Dq
gWkILFDioevyna9J6UZW4HJE6jvQ2JY5asZvh2zUOElMyN/GsjKCr5n/NhcTpBsNguHk+HAwgidE
PWfoivXB8bf1HVZdsEgrr3OvmQXEryC1kXl3WmODKkrbNVUhTmEM7aGoGx/3JfK4IpVtZamIuyOQ
lChm4LvGZE6HbdRPU0iWoz71ugswNnR7PQJa2yowuZsykumnLizPppIYL/rT6XVmixOcStwjfgq3
auOLuIk+zMWo5da0YDukJ3kYOdy1+3sCmEyGoywt1URdLvIfJjYmzf1hjHMZjgAC1DRlt9pcyW1g
rIH6ULHXPbiQouDQkIpNhfBtYx5kQWi8bXM0txvtY+ILkavJgzji5Chiacct9JyoSL1EL9BM3vj1
TsXLw/w+SbdaSZgDVfEO95I2PvWLS/+UE2841hhZJ25Ys1i/wbTeA0gHxQiXVsyZAVW3aoN+tTTx
vNA04lH5xHVuu4DuQaf8e7XNeliG+WljhyrOPFa7YJz1h7XRZNrecwX829e9dYfkNgVdb5dXzZoW
sx6FbqyEe6qLIlzEYsoGLgQnMWhXyNgefGEG17vEPJCuDTy9Gc/bdGGcoNyFzKZvNkUoTH9SK1dI
0+oXyPc18zkIIYyQ709J6SEAA5EVPpeMOa8Iih3Sa4bzf5nigbXCV4rBq2GDvudb2Pn/RW5a9lrs
ez+CA3agzNkXdonBf0HWNg7zOIsRSfdnfzda/VKC87URJA9KhtJK/kJwIMB5qKV+iGpR25D5fPnt
HNnhzg0Q15CGbathE5jYh7N5+uorlEBetcn1rAYy1CVGpVpm4nl9HxP4oHlznvQF+p+sqWZOetLh
gA0vO7gB2talvwv1uK5H381/9aI+an82QnDDtZ7Q7s/YZKMeNu40GqiYwq/QLnUbHDVBm2AXw+D2
yE3ksOHvz0zb341cmKoTEvPwokegR03ATd+YfBlCkfU/R9thi4Y7EYyA37aRwo/tq+5h2I/ey0W7
703G+NOOifY4bp7U8kofJ8m+Xk+WjJ+iD+r23anJmEQVNxxMrJzyqBoez61qf327ySxf1RZd58rv
2bJNgcgHtyHdE7ZGyJPdpVB6zPmQQNRdeXYHpp9IX3+BAO61sTDWlU4fk/iuj0JukdkV5gqQrVl7
CPIh28DIix8LEyEg38nLWm3f0ijmAesdwcj9mEQcCUzenv9StlG5IVfzmKELFFikkaCkNVAc7CGm
GnIO3+ZDB2RlvKYQ1NAb4VQ9lR416dCFHhIkyiumsMp3Y80M2s3m1RKvHazuYPufwKVmD7zeZXtC
WXEMoxB/WfDYsCaG8Zuhmi+eeoc1B4pfkUlGyXxbrXSNg6rz1HE653dWwIkVH+rpl0GLp2c7nsZc
I8BXc11BU1ukyX1LfkQSUjV/jyZsHjYAVF5YLeHYR7DE9uRyCzfHbRFf/rEk1cOThEcV8Xoehsq6
1EEb+CGk6zxqM2dyWj8Xjf29GymGb4sWqXiZh5y3MeRBdAmUp2nWyWPgn5uYEocqsJqMYzSgyXeR
plACm6qJG+BmDiqZuOBrhm0cl/EBLTt+Lc9AZo6HiwiFM8WocGo3APUGqcHQchbJtXf+Jmvxo6k7
RzKEJu6GYT4z4tVgnjTH+JndHktYcjVHWXq+aXqtfwYwX35NI+ZuHsHQgtPOA376ZiRsZXOrFSn8
afql6mgqqoczxhjZLTAKZjDkXRPjH6r1WPebw/SgRkN1bKlKklbaxk0JHFehKInAxVlv5iQudoA/
J7aMedkkqp65KavFrj83cNAINXCGo24gGTZh2X0qVwL1i7C7td6mB9iOFmyV9/31NQA8T5k95tOK
2UMLlfL1MBZJqIRYMRoQi/X7zihACQBGCZOJ59l03hRbVeNgYPKnUEojq8cvr3kLXNU+ofo6kTuI
JO5fAUSWeM80cTBFNm1GqAMAx8nQGYUQr6qq7zBhA+4o8HbUfV9WyRhckpapW5yQAykihdwnE80s
ry6RtiyCKqRoLEH4GWEoRiQnHn49fR8GOsMGVAFHcL9lydeo+yqc5Jnw44CXXoBRKRSgQWMIUP//
PL9pPW2Qhyf5d5D/xzfsHad4KZiQUIORieT3r/CovmaJwfhJN3mWuZJ7N9EMh/ERAQY7e/zHLrWU
Y9bpTaVLXmf3c/DnSpwYofJMDNMhicQNQ/iSAAe0BI/jpD4Yo0SjoKJhrpcC4hOocsmn5DefjdrP
D+67c1Gm6gyboyANW8gxGyvtXh2rmg56uEl31oe1/NVAyv7YD4JujpTTee3nFgM1JROKstp1+Gly
JfBEZVaMQQDje2jq4Gr+E7xFUFcfgvRBtTMaCSdhwFxWdBzAyYTxhwyLuzI+QAiSejJJIBRQ//be
5bThGwyv2TxW8jX2BNtMVeFKqVfc9UrMbNWjufxH7f90LKzsneD5x5FGQH2xPvLd06s8d3pxCYpe
LzI7ohWocxpMyd+3/yzTfO7DQfcUDVRC1DBnhULWFiT+3sln7vsBYexlPB3RKPotd/6ic/UugU96
db9AQDtdGxKtRIsHsOWCRLDwdhCueiYMv/2yd+mAWrQ4XJ3urT4znid+J7cI91TIBbzuaUU0x0JI
9FTmaFvxmPx99Py76GOxpEgKXbf3EnijH3H5OFsC3eJHe1JHMGoA4XBnNAlpkMx3A1MCdxzg2vgI
euc8lxx+Ws22A3d5tg4Is7oxUAaKk0h9YAKmw/lf2QVBpLCKI9bMXh47jzCE4h9AC5fO1YcskL45
ffv0HGUEgZgrLZ7bE1t+nrIxFuptCU3IFg2h3M9JrhJr/BXzKPDo2A2RVDRHqWNx/TW/sCgRVJSV
R8s1A7HkJjREJIsSc8660nc9fOytH67Zwhnso4ZAS4APdnhieTydSClUieO0408JT2Jb4rJ+d7Xu
G65EF76ywV1A0aEh5AdBVqP6TsEhT1WekyO6bz9q+gI/irfG7SH5eCVdlzgvtJ9NsgbVUsM6yij0
/YprFCIfxbyq4KedfOhDORYI7a1g7jlBIQkx3Ggr1T88Q6zGYXDOfLV/1MudhtVYOFPHIRFB1sGD
sGOkWDrv3B7+wAj1vAfe8kJu/VkbtBh0OnteJfpqff6jJeDAVBvu3/bWSC3hbMA89rOA/1gBV0/H
NbAlDiBkpgowgpxseQkSsxBftsc1WJhjV7KUQCaat3ym5nf/iM1B9qn2WXZfRFqGo6qJonSSI5su
whAVTyGvHriHDu9PZWw485Wwme270MMC6vxGyEve6JptmzxdjXwus+McRGpjd9mrsHt1zA8QaR+N
5XjA7Mh+x7wDKLNpAtqqCgBdjwXoLS3tHWm8rqS/3dC03UYK62zVO5NZGD+4jJzhuWGB00NoszFS
B5aj6l7G+U72kZ9jVy2b+ig0fVgpmHcYxUm66H2ub85QPmAcJp4bdaj3WFV5rM8P/sF/szmSBeBI
zaU5SbMgPha7u/79DMivuY5uZrHCnx/0qscomjARyaNFxPP+CM3Y4dPex5K3XYQomUE4PIu4x28+
0XpSK6LLRgc9h9Bg2/21mSmnxeI9grq3bs3B1fVChSsEjhfleQC0Jojim4k+d81VtMe6yMYLkzeQ
cFXD0tp+N7rEdGYuHxI+3GTFk4zvazSs0bJeGUGZxmrK51nq+9FpfiT8E9TCNSqTjWQxjgByswwU
SA3m9FHoTo1qwGKpWOsVBlK5gpjxeoW+de7T6Pgww4k046VD5So7gC+83Xeax/+9XHNp5osw3fRJ
vdBwZiWJc0NrN1PKcUhVkmMBaKg/YGiv6oQgDUDpnJUkJJP2KE9GniL9uigJMu0vRqFKF1D6rXSk
zkImd5XzoxLa2YxzOqLlOE8rzE59E1Jx7Xhtc9mK6xtpL61x8X44Im74K0tVBZl/hkyBGY24l0PP
hzgozopJXG9CZU5rt2lHA4y1u9E0gcvJHv7qhgH9M/5FtTUkUvg1F5Wvdczik2kj7yRUh9ECWqsL
nkquCYBqtro1uTCNdib6W7O7MOdwAYq1d+K6pLt/Aj2ruE8HTjdNZCeP29ufqJhFj4HEfEZzFOHQ
AF5K2lPLTZoeRdoAV9G8tO1icI+pUYwn8MzR9jRdheXEVkQINx4rNMnbmQ72wiawjQd3HAitkhVF
eyGxbNUObSWUisVNjZD9XkLKwcY0pWvXcMe3V+MYV6BxA0ixQsn2lPrO/8UEZVGPu+pBYuLRn2qz
Cerg5LjVq0aMvPGxFKS6f1EyzVzEeZagU4Mz6Q5KWtxF2fTBkVOtUkiJy6VQ2uRsj4XiBSiKzZZN
K9oLndfMzTrsnP2NleJE/iS/QufJDvxWLKYhlmr+ruFO6COfUU7cnN5vDhbxsnWmi6R6wO1vr8SY
ccT8eCGs3eg0acRf10k+0pp8GVQkKvqr0SFipMeym945qaqD0UlqUEFXIX6WuGxMaxANxmz/eNrD
KBadjTTMxvfYc09g3LM42mdzoB+Qmza852t8PAi9pjvoCvZyumbGB8wpE+r2IMnAZl6jc2CITLlW
wgO7s3nlohhnmpEzg0Q2qCspaxlA72K3UgiMJQ5D9zYpnZUCR42rs4N4amIaOihTT3XorGHaEu0M
QFObHx6BIv8lRGSVlC9oANuygn897IgrYEPSzvUABr4LdX4wzzrsu37Ofyw9pHgsT0QT6mLoq4nZ
DAYmgGtjCllHVBhyciclyI/wIqAdfbGLirAClq6UE9iGcyYVxxhyVxEODVREwpiGPmlTme+LkGqC
OQbfJ/QC+sFCHT09vev9pgWHC31nS3BCqSwiUk5Y3c/znkdGvYk8Px39QjR6bIPU+2QY2BtfC9rB
AyqNFF/Nhpd/0aYD8Q9Dk0ITfm99xuYLsop4iwYlsHyBe5QI10uVEwn8h63FUCtIYxAA2PN1tb9q
8DEoRd5u5dmG8oAzSmlGokYnetuhgd0LQgqqUxGHznXodiJXMBr45b9ZqYf2bzU8YH2Mdyc/Tbqj
0bfl7pvoGMKdwfmGS2Ku6nOMVQ0YXemCqV1U10R2LLMi8PkmVko6qucQ6IQAJ+tUknerOkU6zVfB
pw4+IIhbnuImD0XuIG/Qmz0IyemvqB4qqP2/+eQ8Fh8ay4ZxZZuV3+Uk3icJVNlphqad/rsVTl6s
aV2hM/lQ7OBO0dW2X3m5UisTdqw3MH+WlguT2B2ykeBvYoEZYyLT6pti5gFflW4WfdIDRFQQqX+5
dDUKjeN6lNn3vTVka1EhzeY8qMGM33iTQtLBLTgUwLUEZANgXpB536ICjpZ1eOfiieSJsRdloXDB
nDEj0BTo2hz9U2aVfypHqgv+hUTMYibSkz1pALj26LQVswr4QWTLcRYcSKFLZ4p2i43Tkyjoa4q8
IFo2tWZKkpYEVP3qGviH0iKr0L5advHcEfzA1W8IHDY010nhiDR4s93HCS40m0tSuKIOVRkjcTYB
Ifzpzt8u+OUWIF2xJ3MKNRJ0pDbKx7bUDik5jcVhM709Bmd0tSg8v1gz03vCSdxx/NhAqmUkCLTY
W1jLGOHxjOZrJ8U0gk+3BfK53NtlJ2CsGzcdlFH9J/vbaW8FWwUP7F4/pGSaZfu8xQgavLdVCF8u
1uXjvsfQsugAlNVSrgmO0Ked4wgNjDgQgNJ0TUXzvfCjZEJZ6+lB7yQWOvJgSMV77k1CY7IOomTj
iIu5YCPTfrFuOZOW+P4MslShDZtOPBYcLGHQtZizhi43lqILNnfQly0aLpI2fSrEQAk+lCBXK0ib
vddDMh5TNhLbddQp5/7jCJerOFItv6qwdaqAi7uAcT3mwC07Lo9lWUWvb/U35MZNYk/lRhmX4qx0
CIy2uhfS9YwUSGkX9ah2/LtDHsKOpI4zw/fMhYhFn9IlDHMmf7aJzpgfTg/tvhpHhlaRx/wsJU+p
4YXLlxjsMDygFTTh8j/ey5wrEKVNsFNqf/VntT5mF7qqw9aZdJuF/DiUmlWbdhJt5tNFQUA8WrIl
UWqbuVjIyIR0XIHc5T17LIDla2WEv4frdhX4P7MOl6IXUh/jzUWjCbWHLv+nZvEd1TYr2hZGgUut
6ZuagHjdT1xLbaoSikHHkiLf/142WIB8W+hDNPc0/levqFZdSE3LyOgRE0Nj7TtnCLB/XWqrCnup
muC6q1cogZE+L8VwojTs3HUcjN4pqPauHkVLsrCYjQg+kI5jVCxU1WIudMATRt/6but2NVR5XBJm
0ONe8oXk8CKmnwhKdHZQtNMrVbZMPZZjRXYrVWEfBVQDYqhGqd8ov9YsC2bXsjj7nblda1YFwJqi
FGSY8xlJTVhJgwYt4jWYF3bRIm1xDMMignKwxmrAVpu2z4RJ3Ln8NhC9xSEMSRrHIih/x31rXWzF
LhGueh4Q5el0F8lOZ0+z//b5NnGMFj7iFHDmul5dIhlqdBZ9p1a5dGNxm/LNZccIMkJFZnXvK/Iq
tntpzrnGYTJlYg3BGuH7OUC2qr8hddVXsg9DYuqr3JA6d5CS8GzZzzFt1FIoFFjowp2badgGTfHH
e4k122Ee6fgeyVZGQnZABL6+PaFhsE8JRbKFaJ0xX3D+gQP6EWBk7EOxJMBy3iV+Np5I1xGsuNm6
tEHPZQ3MUyHL0atdgHwjHRfxsm3IucV+V47X5hEJ35OwQx3eqJMbzMWhuqDZ9Ic5/7mC2ciR1nYN
dP/fgQ3fxI3vAu75w+FBzLPe/j5VZtpZHECFTILYXLBRLZOilF+JGZYk8qMdZqv6bi9J6kW0aDww
B/5Si9gnrQTl5EeZTqEJq//4/rtYObxDiZIDL822CTdRopN5HSxE/UtrS+4S9eZbHKfBPkd70XKg
7kCHMbUrMOU1XnuBQx2Y/n7v+NMDGdaD41qVwOdPankCrJrZZ4HkDq8v7YO2+oPdaZPBjKyWJ66x
7eCSgZFVFPM+bFfElAG4/FvAIksP2FVCYJDaEk8N5UrrG+IEJMYR/zqf+nowjWHrTNbgF04/b1zj
LIV49NBu4bOH/o3PVOQtBhYA7+f+t+Qf+pqI/N8dJQI11O97BXOVxrsjP19+k4F4Pu5n9nd4QtW/
OTxB+5iAFOYUXW1ApggbgjPOzaQXz3ufj4iggnuP7BKYJJGblJuLUxwKb/lAMnvb3ZMcWnL7TjUa
3O/19TudG+4knUVEIBnuES5DirlLT8zkWJukGQLF+8OvNL6XTAiIH55TVhUGiX1VHQT8RWvN3ADN
1Tz09727FdVd7tgOBE29GjchfvqQGF8ZoZHwKUqHHSIU4ir3X0wJg8XLPCzVTLeB9Hyww+wnaLJc
SNi8FuUwP/4irz131SYiwxXnv6UMGtEDKpe0zxQvkGU9QMcV3kBa/2akVWiqQn+0yuQz93iyZGwh
neEYMF7duB0AqpzguxrrWXO9M89KaN59veyCrieWHCkAq2u56EzmQPWXH37Hr8qq4k9Vur7HRp+j
NZONQLKMFmEfOwPza2mnhTze3oh3eswoxgwjdvv702VCVD8zSi7Ws2cPMJXsHcLVEa5JGfO2+HHL
ajC/oVA55x/fn1NioGjcjghbwcNTsgXm0Ry7u9+p+/gA53EmKqSh8xYyAjEsroAMof1DV0Oa1g9+
xKQu+Meaay3uyC2v9zMDQIeMbCuJzaFYyrHQE0GPWQudVmYvXEG/N+Cquzf+q8AbP4EnXRBfAlZH
G+cOiDeVNESYwxJhpqNoZmMWOu6O+i5rX75AnoXJR80NlEN0ios74GvE1dJWR6F9l1o1wdj3NIPV
67c77mDr/nyRwC2t6m6xcyp8jg/fb6EtOJtId7X+MtavhH/yiFMQdaGrKELlj1Rds9hvv+q+nwZF
hkIJ2jKv+Uq9A+0Oi7zJD6LG+dWVR1uBrdjB39RouO9o3mNgaD1LNUze0eYmn5gl+gT8UaNJIXhI
2NQHxafDA19pv27vek7UtoP5I6+GqIoZ4Oy5CFA8ha2Z8kaKA3uuGxwlAb+jaCYLT4gNRwmREJZZ
T4aECSaL9PsOiq8vDKsOrc0+LyPITfuXC8UpzApxIVsdXCuuhzkbns3j1izjH3XnbIVthLTizhji
fUWawcrMoxVsDRP4/HxX7mPQzN57PouS4fhRGyMKiN26E28WqjwSnDC12zTwPTqV/MvShPDxiwxD
mICEFFirdQ+KDrbXyXXYXI2g06XGr1d2Gs6O7B3+ayQuCszAz3KDWQIBbaIfdETpBiz68Bc7kyhJ
65pusn0QDp9zOSR3W/B7LQkOePAZW9q+1X4NQSwjhdJX5v5sJNiHg+DSrmlulG+YqLkJd3mK5Tsb
T4BQKc04u8VtUfmE9vXEyYLfBpJE99DlX7fz6UXib1/4XnO+ZnsGlh4YLZQJXWOIanFFpbL9oBcM
d6ZEE+huiwoKeeklz9dxRPjB2uSeNc7Ub3XsuH3686OQkJvEmbVNFHuWWYcFtcqCQB3gp0goLk20
Ive6ucyQFniK+5P/mIIoR3zR1y9NVB368s1EIGtgnvC7RhxwnYD2XLOvbrB9931oz1H4t+hjVsQa
26S7Lko7DXSs6bjFTYkkIyX5ZFxxYG5gB2IlqDdjViR8lbLhna+xgWG+NAcEjivnTq5OOZKgIb0G
pBBqbXguz3gAoIPoJ8+kIDxOJwNMfKMrVP3w1cxJ1XFuAVI3DrFj5wPk35HCdjjKVbPdqiiZXiLK
s0IiE6UC8dNNI5VYDaGMDfcZsMw9Lz3P/ObA9jfdPbcwb/0WGx7MrjuKhK2EYpE8ukIcvQO/cVvH
zL0gDk8+TVrNCVL7F04JqYmuA65f1uMXMUf5DZYxatceq6u9u//y67cYX5Yk2IcoEzKTf1f68rli
+JZApk4gKpjX7XoO5LH8VL07MR9EpjsRdUN5YVdeRAbcG5+HEMZCXFFYE3AUtwGrlzJ/VWacfp2g
ZvDBC3CJo04qfzmfM12v2/DzyQjh/D4HELdYj5VLxK/SnB5mGEDX5LVIuLgsOt8Gz1J3EmF9ubCb
JdZNMksWAb98uSJbafozmYQwhDoAhQcR8GIp48Qgjfs4RVvzzf3JTN86xz2ur9xF0pVUAfD81Goz
cxs/66/915BUhJixHm8rkPf9gpd2SGL0UddG1DtvcTRDCqAuI22thfiIaar0EYj6kYIfa0rk1+Ii
vw7013tAZPBarCnih9gUB1qTJhQUg6VNnLBbkkNPYXG5Din2y0oM5W5ppbIgph0LeUVYoazL74I6
57Ig3cakoVREcaQj/5iaROVsw25Ndm+YKC83k95V3WaAG/G1gypuLmjQ+4IL0uVzywweD5JHLLyF
FluEgfblQpmBGOG7oChzAz8A3xy6K6niPfjFSmruho1+/DA0qfTrNDO2RF6yhVNrFlB37n9vqIqv
A50kJtE6Y+rnJwQCwJ3O1fGayupV4x1rX5kJyz6VvYrmdUgGDAvH9tJp4ukA4Pmvdj0GJUgAzo5C
qTUnRmdYoEJQnPBMvUYLIBtT+r48qJtKpFFvJjHfN00AvbTfFIuTjVCm5BvWI8db1TvX+tfGizNs
gm2r8UWS1zrjNdM12e3g5c8sI6ilu/M0QGKJAaOovHVq/RsJksx72mQTi8oFdYm2up32kkPW/ndn
SmVISkR0KQamBrMvsqNHT40Z+2QXY4L+Vwvf1mGtPRXcvtxe4OYPy+9J2P1V3nTIsRS3V4yWkRz2
zIlxYhhEh1D+2UbTt6hvC0W7qm4l64LoTNwmWEoebP3oTcjdGDogA6HU+K6C6fwix8tDZu/PlIgs
cbxuo2jCW01kzI4Vz4WH8HtLS5KARSttVWiByL1O1mfgnOkx21IGn0e9r//YrBkpSBNrlfa8E5qO
0kYFtA1cGsVi5F4beWmhXRQHMkPoB/IvI+9W78MPYI84hwOn6bH2tJk832tPNE03ZzL5xVN7hYbx
Vxss64lOW6G4Hm0WvQb/HJzW13w6g44g/XnN2a6aiVr8guK3S8ZmlXyq1PyWwZGJsvQsCkGff55Y
kGP7FnCkUwbnHRSvCkfwrQZQNR6+I/NZf9Q9IHrjudntucMNxPphbyxHcbP8AcxplUzKj7tHD06Q
FjzC0MI99uDfg6ySqZZbC+Gh2K14Zn3+Y7APffSwVXgPf9tdoA8rgzxbwHo+uwX8sAmcoAGdXVaj
qU+TvUQ3u31tz744CIw3SFolzef4x7RKjFMpcJONpmUZ20Oshg3l5GT+0pFJl8PhoR+vyX2jwS99
mSGoGJG7Ye99TOAPR92kRImEHnLzGZFKspW97Zubflmrsl1x6yY2HPbPAnxSTj1EJz+HxLJH92uA
ZsODJ3hRx7yNfYfg1YZomhruqwLghetaG7HmSbDXvN7Y8wd04CJL/H9cObcxizkvSptPKw9f0QW1
DtyQmXgGyYKOJgN+ekYGU+/i4AQHLnDG71EDiryLJki7zcrYZo/Q5QD20iDHvVs8f/dUbs83tPZV
dyITXPe/ikprZ7vP7oSDwcLGYE7gGBJIOtqSCT2A1b0Mf2Zfi46KVfkMlVgmM40il8NLLv+QVEGH
NKh74macmr0E9kKq7WV9pvodrBF8qB62ims4+OTMAxABDFK99wCuaNRF48ukc53YJlfZrKGNoO44
VkQ0AXcKbyhAIhDc6YBCxMsceFRL7t8ebKFTPkhMvho9n/uVfvVfiOapr04ufzf4lzOZRT54ucH6
Tbz4sIpwBApGxSBZ8ggc+9b0HH78w5Ey+GfsRhPBv2fpmitXcN2Mv8yX0zSnlIlsqignCZczRCoA
UrUBQqyLyMqMJsWezwjZytVFXWLAy8DS/xo0fUIsEl+JOVnXwhgYDDVgtStHrejw62m/3D7gygo2
3b1CyqoQwl3UjA3nO9SRvJn+8upZwdC8yBQ4oJAl9g/jvwWD4K1Z4H+XnAGmPdeIa+kq76s2/WeB
Vbh5y0WTNU5L1VNmzEDfD5+GNrIvcLv1VL5DCMNvdxA7+1k4B/q5N1Y1nPbaXU3JgfTjijq1lDps
XE/a6WATRBSe+Yn1wk41fXn4txEHOaW0KhqJavkjdVUQ45u7/Fq6R98CgX70P9pWoNWMIyb3qM+3
NjrOm7dL6fmdessWH+EYdJioIhBvH0QE/uto60h8+q5u8M7yq5Y4ttGU7DkTyZdUh3n8jBvBFDhI
mLbjlMG8Nw1eJHgHjNNuMWRkJzDaFofOxVxEo60k9XdeLgeujkUs5I4rsf/t/RBVd6YYL7fqCNi1
A8Vs3PAZHDI6JBci4yWudUx540jYD1sIuDuDhk5h3V3D6HIVyHNUYQ/iEpWjVWBLHg/ME2LuqEq+
CSCOfqCjRiEI1fJ5iyQgmsM81gtvSriNf3zRr2ZNQm0qeREqS4x9mj1U5p2XJf97Y/FfhC8eLhAy
+pOANmtFwc1ZW1fJMmL9kaeTddj9rTorbXNUngMnLSS0OQ5ofnqkGpgAUnYZ1aLvoUtmIKvxqeFE
+2VXQcMDKgb4lNSChlq5IPC1BKjpZhhvLocdAo5iTwep358g3i06VFnDuOAX3D4X4yWOzUrR9Dyh
W9HdDdT87mUXAgw+wplcU/6zhyLxf92TaxQhggAvt2v40ItD8OvgQyFNCwruaKWFEmgARtGD2zh/
0th2qI55DR78JPa+qX27eoLuQrH+hEoUmmuJ2VhfRY/HVhICFm5Xo3CW7JAL4Rg8ID6Y3BTe5FxK
toYiDIfJkskFVjaJzs9q468uEnURTCcG3YnihxJrsc4Fc6pVRMbuBsrGz/7ywLWmihacxiwmnFSP
AfrKCocV7PyBVSgLFlezc9wRaOgQ3to7Vw/M4iL2l7bzEF8A0mgCy8j918bexLYlZ1TjdreS5qGD
5vAM3nfisUhQZMftnVl1wezw3CS/MtceMVZpd+yipqMTgCzg/pfSQYYmkYMEB2fIwjUcjyWu7xvM
MhESNbc4+huxLEu3bIZjZUmAQMm52bVB0LNZjJnMcryauTA4WxOqngbeXzuRuvUA8679FyR3zaOH
l1Oj3KPqzeZkRPJjCGxVrm4J5wvRG9Mmghy6XYljwJRCkmDMMHhCuZKDPbh97kdHJHOjHi93gvED
+aIsvkABZiB0ITvHiC6tjiH3u4SPFvc1F6NGNArAiuMRwtEjn8im9SSJnnW8ynPASD2AfAaa9Ww1
u0bAoz0vqOgsBfF1ZkI1PQpny+EZxtePvDNHjvBSCJJD+82+Opa4VPMAE9BDsJNqZMCQ64ZNd4h4
ymDMyrcdURvAYqYYJx4jbuPBDoCevItt98KuSub6NGj1kPRM3qNxJAB7MaDYCOC2a8sDjtMQCGKS
53OzMA/jtn0PuP2HFGevy7l8kL3rmnj23NOcL9VA+ibcmV+gtji7u+r9L7qaVQjfPvCFRAg8RKNt
bzppvcbCB2CJxvf3Pix6EcHl42tL76BT1gzw+45167klYwyvtsYZsWmtI2O8N1VAv9uvqS8PRa9B
06uL3QAQaAREFP3i4KmOhpqJE6XhcwCPdFD8klYfnrKilHoJMFNS7jOpg90fytmVahy1JKfg3D41
BHkw1owQSRRcx3xSrduh4pHXG6YrcLnRPwdBa0iHsTQ9UY2oQyDNKmhY/+ZCgMMDCkgR5vLvywxT
KMWmFxV+Qc8oiGXoAiKU5mxnBFlbSJu17UhMLlKwFcjlZekdgrHAlPfIVtTMvV72hMaGqkISXC6z
tKSxzPlEBzAs/gaBikSh2ySIS0F0boCBC+gXpp3s0YcCslvrHpm5txmxmWKafFNCnDZeW23NP5hG
JM0qao1EEmnH+XIe+Oyvy0wVB06Mc6JKVYMnEvrYQ0NR9w0Bj8rEXyQa9kZNJHddjhKodjgDXmG+
mXAUqogDJnZaQ9GPKj75C4Iglb49rJ/H2lMOAFN0zX9EtMSkiarctkMR/NMBQqXgnjbZHi7vaXdc
x2l9+u4IbeEeoe6wLgAM9UjFBhSErXQIflXBEf3AJqrz48o3z3CgpTHto+EU266DbIuGN+VprGjH
muwrnDJMtNTC1/FS2MllwwgyFj1116F+35RoF83GzvZDoEutKwE+1mGNRl4Hx11so43NCctgN9TP
nQc0WDd+67/+5ZXJjX+7ajYl1LMojpLzawPvKiRGNWqZ1hssRj/zHExLJNYRdCEYGyQlNr9joCUr
DfhVtKR9AMHhjLEj0wnI/ugm/JxyIPkKmxef3I4HUXAFB8hGQf3z4gsm5K/DFFvBEsGUw1HF2ty5
J4focMbaMSIqncae/fz+tm55GsDG4OVLqZqZjNGBJ9JskmcsiOXMYMiOWjHq1ni1G25s+64pBuk/
94N2IG5I3O1b0a273EzoUh0m4JLKjhIg0pV03nAU7tLg0t/gb4YFgw77xPHCx0ji8pJFKVccKIN3
xfHl6P2s3yjmgTNPIeHK7uTBYj0vMbypIAndoq4Nkf+/VRsEkrC/O5ieV5kQIbho6U9e/2mKpKl9
ZDU9JbM7JY2gaSpO/l6AfMQiRrboq8fGfhC1knZc2JuH+S4+WKfOm/+ATAZ+i1C7umDpefGYThZ6
obR1LntAtjPepmH3y+ckCPo9YRMG1F/AglBBGyoejmK4DTntwjdOi3sx5GC/XAApaEp/9K/+yNsQ
lJ9II7z1Fx7jzR7bfXAPJhtpZlBrtXplo1Zq0xmRgSp6Z9RfX1WJU9VdhvduWzRdGz5G8pH0XYJy
ead5GZ+94FOdqlLaeAiwv1Ou0SjrmBbGxKthR+AmDKW8rvndqdRGIoSg8OJ2/nGx2uCS3ea1WP0V
+hSDDPG7jDZYFVpNB59JSSLaDxuv3EVBefCE29NkpxesQs714GY4VEInVL64QkGrent5gB/xm2Et
uYoeUoZxyvnxSs/ZTQHhrosmL7ijM08cR6FqhQhVAXkxFblnA0dJPYnjAaJLP2ks+5zWosBaxtQ9
pYuTvqlmy/kb76+X3Q6NY2LBTEaxrZFkRy9dTElVT+TKTpYiRSMtBb+t3gaDRiPmw+fWel2hEhab
NC5d0EnoC/5UoawUTbw1g1G5hS5CZ498g9/e/k6aois0JIKOnTsfLzQD+SoWCf+neY8Pe5Ag5ygo
/cOXmkfc9hu5wSs6y0AVQTJGtqsjM5PeWrHKBlpZ0nl/oN61o1ghY9h00gNjKRFHQ6ZuygiAuFMk
uXH9GalkgusgDzj2QB2GedqNQtUicKmH6OwgL+H2QbwaIdtRh5awDiEFYHNqAvoowv6hPtp5SobG
j4U0/qLt/h5pAjpF5RcuKoHukIM+fBpI1/ZpFUtSVOdCkpVWCwRZHYuID70JBte5oqqBqLLcxq2b
coXOXrTzqG/bUJXbQ67MkP7N3wVc8Sr4QWovehdQhz/ZhXWzi9okUzkQgXFixFiIoAP5WvcEUZkS
FVRU4+PsPAZtnP93M56h1IVLXQ/ah6OUN/zyFORCo7kw4EMNDNdlqjiecmElW7FRTNJFSQYDpJ1R
+wAzSKc78ffxNsxH1yutMUR2nYjh2ZrSisFdSPAatCT6B5IOlPQvAGVrHKP1zZol9XjM5a6+gMYW
/YV085MkWQs+5siRP/pBAbz6njUpe5rfodtoj5Ay0TT1YA7dhFyNrmLJe2aQsiWBbTYhRWCO5od/
N01kQtLJml68lMX+128MTfw8USotk4pSTWPL/diBg+RogBQJs7fuJwN+3dXQ5MGOUC/5gEp+UfC3
pokfjNNzARN5g5YOqWTWDgw+uC702qq7fZLn8ZZP1eheN7plU4wczyGhj7aec1EJiOpNzbqb9eY1
ks7n2CKpePCyS5lTfSKRFY9EbzMM+80fG0hVwf3TrBzHBjjL2UmL4ioyXlGRbVyB7GydSyNzKaV0
ocW9irBM5Wa4EigONh1fHnexaQ3YpDjLK+KKri75SdeX9mLhb3+QVgDVZYH7ciyln36fkjmFSeEF
tvJ9DTqHVajKzA3rJYA2VPmWTgzUDmE9waJcFDa5917DPaFdbs8MLt5A28S4jWpa8b5r+RF5UEkB
eYwc0nhUa0UJvysQJL4ltkAnoh5j+XTenofB4Tc03oyaeVvXzVkYsmxuXMDseNlgXQXLulIPxAoB
8y3eM1OWvAk+iBhelaWLsoezQGLZwjodojwJUj5M5DueNZfeuNIgB4/D63A4CGEWjxe0V5bYN41X
p5wmBPhBaJrsnbcbaLPyaISN/suKw4jPEA7Gv/GoskruwpPCQ/Zs4LUGjlzdAkZGQFXk16ASqkOm
Q26b/3q9uaroqSfMmFVitygkqgDzhDIXxrEWwNS4AscQgOmXxcEBLUK1reeihCwj+Ey8TVC89xIi
OaBBrzmV8I2au5kmILDn8IOSwbYvUtiEvHphyeLYFUs063b15kjIMNFAa1TrmslzRNW+ADi9Ws5W
+wBg8dqoM6YlgirVj6Lk9rGhGLwL7qogaSpvRdV7qUGfxp4UZFaB54APFFN7XUM15zAfIF78+wAM
UMfSO3+8cFPK6u0Sm9JHBfLv5nCuwQ7vxhL1f7dk0SqMl3VqO5qQXdidN68U/r3bf8bKReUZeR8o
RaRAmeizryHJbbL+8AYhT6lwaJlYv+j/yOZ5cxdtyuNvxun735nk+NMJhE/L7Y0vhtT0cXP1ANLZ
OB0Q37xV2zkyj52i6oN+l5suZ/0m+bYoFZrk/caGvjoZcTT2k0CoKF2zG9lCxpRp/0jzAzUGVfXA
oNV56o5k8rW0u4xtGv6DJyM01R5RJLhOdA/TI1AA57M4JxcT/rHPm+Yk5qVuR8bglzgvSMP4ejde
/Gf80vRzSWNOJjC18aUqG1Cxyn2bAXMZ1T5Tbl4qEB67hbJdnYHBRdo19E/mlNey0OXArTE5IkD9
PModv+sdNKlTx0EPYT0kA22SyxizTCS1m+pdN1DKyBX5Qrte5FbPVnvCHxoPw81mODHfx7r9CleD
hcqx0zkVpbyDBNol9t8ZGfq4b6prX9UHhqKJd0Jn75vUdT8aHu8uNlSdRr6Ph62fg8owt3fzYPo7
e5qskIAk1Kki3d4LtbAxHRCyejLuj8JZWqy9+SWaxxHO28Wo6zTr9apAkPxM3Ucib9oZfYDeSXBX
6tBuXGnRAxMS5LzQlLbzTRytUntNELpDwjzUIWC4TWHCYdPlP9kdhn2tXh9KHgvtbNz9LI8iFKof
5mlZjXriaHOYPKdM/IeBGQeVvx4x7zb3y26sbL6xrOVwRV24CZbCzHp/T0MkaEgmPLranfPoAL9q
YIVy2UECg80pLaX+wAOyYp5RNhcPSEoauCsskHwB124+z24z0WTPfGUvZd3vkaWXiSoFbkBJXR/s
kHMfrcVNnjgvVuP6a5E1FyWAAusWNe+aFV7VnX7HicpEYp+we0K8Z/DltcPaPUuiBEm3+W7nyZpk
52Yxk0197qhLTZx/nPv4mzbfEH6qgnyz6CN5rtDabvr6RIiRT/QRnj4st+YTP5L8t+H3CciF985i
eTeXZL3R1TEHZJxmORgEYVXICDkCvk8AlaoGjRp5Y+04iEyFSX+DZsgqfKRImLfpIy+o9xBUkJBR
ddEfYUJvbrnFS67XcMV1rA8wPTNMQy79h/XmB2sz5FgsYStgY1af7crtVG8ukIseHaB6+mzKVseE
XkW87AhrCionm94PMzcsWSH+NntjLF83v94K+Ohb+W9J7mW1B5t9TiD+3MoD4Jrgve45SgQ90uT6
e7N98C4UIAxxogm7jIHcDbivVVNuOuX90+9zULU48rAHh/7qOVb0GsTY4CF82g/J6x6j7JX39AF6
+eziYekqphTRnompgNfbY8wZm7qyZjqwcjgsRCtZWNACf0wdfdwgpfy3ktwHm/b6ayOtIXcQMIoS
N5NXdEXvItaYjSIvKUaD6o9ShNyL0Rm2unV5KN+D7fmLV37fNmVho+idc9UuakdxVpcuZXkhd7DU
FRxGHIjtojM9BjWMjrYBIG89j1JRJ1TPwUt5lK2mY/E6NheVSz0nTybcMlBUaBup/SiEKDKXkKWr
9jzkF5RPDbkpaHifgJ1D01Sb5XvhmLa22CfELXjYZsB8CIuoUvAML7piJEwU4xHILuMZ/w/k0gyX
6yOJkPY4SoPlmMS6Sap87sN1byt9EoqAY3bQXXD7zeCINAFLTksFSIOnNbuKxdwEMYrRNiamPpoi
oDrW9FjJUbJCnTsKGENNRfq6ujlPR3p8N7xl+enoe+V0wTCSaHO1F8TmAg6ASaE3OStUNptim08P
xKzWygsn9XkhzGWfNF1s7pWrrBBQfK0bot/5v0afI+hU18tCVBUmbgxSBKEBo+4jgsST+FY2V+lu
ifYXYvTGWN+Vh48ofKnvXgjMxYLQQukJONcoe+R7ezlNSQlKO+Aj+JAW1oA2X/T3+th/lPHU44Mu
bW5t9myOjmfnoF0HcUvR44LqK+0BbPvye3sQBJPaZ5q18DzO1LDBh9akrDol1ZWySCSDIwEn1JW/
spW3am7NFzOziNGRjAGQCFEK5RW/L/kOPmah+IXg6jjukKpJrf31CPpU3C9cs3BNihqNcYCsyV15
4cvSlJ96mO+4v4p71HVd9M6b6aKCEPa3VU6I8KsCVM8dlzxOiJu8VFJzCb6GzpPd18KtVC08Hwd+
z6FuyyC/Y0RfySHnGk7N0Tmb6/lBON5sod7KPVSLM2vBTQdZyFy9PVDistvQEI8PGHA06IFwTutD
sqeQxIPiGntugLY4Y22Z8+r8vaEd2qgFe78cZCF1uT3Rd8n2ot9OsW/WST6kYERK9s0MtwI1RORW
EFRXmlrJcW5VrDKOLAOm9p+rsMJuVl2a3mFtQKigIjv2P4+jyeia4ZxzRypuDTra8p7mcbuaBQqo
5mF8UUL0u/rCjF2J4+G1k7s13i1arveZ7a5YZz5m841Uvw0e3Jgr/u2jwIoT/U20JjYXporPgTNn
wlBKbehZibkDPp6YAjzsH4GLC6RM+UZqYQ1q8yxScUBlODF5czN94Zv1i5y37VbjFLGf/ANED70U
+fsyTuDpmMgTJTE4xZBDwx9TZjrsikosCRT26ICatwtaw68XtzMDyEg654wgcNunyvHosIJAvrEJ
ayDBeHdYRPSkGNMgtQVkP7tbgBZlx4P8e81+AKR1ST9ZaAWycc1kYmCu4Xl/QV/qrXvYPcpxNdNT
W53w5ayDip8382kw9ynf4s5A1m/ToDj2oXc7Nz0vKnK9lbpq4HXwYZqgVzafTJQzpaJfzf9awcVi
VhRaTr3T9jgqVbq8dwfas3YGAZ6ErfQ3lxYbPhJX0arfk8DOHnrpVFHTut5BKJsClx19VAJGJNA5
i2dVL81gAN8WnODoy1lSfGhg4POaQo/YjGDdK3uvlEfAHNpVjZnsmoJasUXaNxOvJNwfoFTdSBFA
iGmO5qDBmZrofXl83EO0HweRUVVKjmlQZdlob9/GtCtaSVQg4xXT3RGVbRxSV2rewE1iKdYu02vG
vQ0xtfrKw4HDUihVUk2T7iZw7WERedkSrBa4O9xqMbLuWbkST0KH2sD1IC2wTLiTsosgiaQNOXZA
lJvgU3KQo7m9mCtMroo2X5vjmPXmeHcJnIz8pqSEOZ0vNG/0LNKBkpv57jKyq/6F4E42BKq5phjb
QnWEQb8bf9YhRIGHycmflwoZqFu0iENVgDpbZDmnR0AGfzpKVlGDOgBPooaoMW/9wUA/pBg5y2lD
IlrR+Mtz7tEtd4J4j5+BZcpszD8J3qHlzectOq5stF1l5VYsJHzizssGXyRNqfCCbBXKmTV0cgdC
KlhywYpo1eTxxgZ8VzF3i/84o1hVYvwdGSjskbQEnenDY+8EM1P+jdVR/OsSs3JbZlx3kegs3sFf
qAX/WXi1hHxa2tXe9MFCQgbCWekdhE8myHP8pcq3s0AT0MRecGphYq+lKW+C6SNTQRss+E2NfA/A
ycOoojCNv8P/J39O4KW3zTuOcau99/Xw9R4k+qPWlw2C6QgUbiYiYe9U4c0D4Z/p4lx8HBX2lDnH
TTfvqYbIU3rV8mWrWMf6rsnLLfhtBHwPyyp3JUY5aNRY9L1q3yKMEgkgQ1V8YArTYLdBLyRC2h1g
LHj8+qETdWoEJEVDe8uJKqoOZNJ58pvTBfA43p9yMG2cGDiM5sC+u2jGJc9a/p4gpe+80j1AKHP0
IBQxpkmtgs3tcHTQijaJ7O9ApFkdL5hwamJDOIQnLT59i4rtotiL7W018qByMnvSM8esm6/HHvxY
jolVzWMvzns+6z+wkXBp1sRBGfsHja4/hiQd9v4I3lBv2bytCIOAu7DuzMXJltMxNCbVvTy6WooB
rFhuEv7rit3xd01HSz+EP1OmYMTqMjAyfDHsshdCx9TcZxEowRrevykwTEt6YHz+KfNJRaPxanvs
wuqj/0rJqUlZA9hEdl4yzPsjKykQZL/esOpgUH70l1KyC3O/6dofy3zIqHoclS3CVipSeOA3BHPe
0p3MNHwyoRyRPVbOu8+rj7ZKoGHom5GdNWPyojAFIUtvOfeMWbnj+P9eP7h+tE/PlMLdMmX2NAsu
AygJF/mV6yBDQ+ptJu0Toiq3awQOQFkoM86EA82Gr1Pcn+//xHGiYlUGLYm8HsKi22zkTCc2Hm5E
Yqwgpxlr+q2FFQIB7Y8/eBkhndSPXmz/EuKNFwcapv/QgMwwwuQBe067TLmQg18Gp5Yz4arruoOP
hFNoJ9gLk5FQGckCr/qrET+CJ7GewEmVYebus96+1PujPM+uvICrpZ9fEeqSrWoak+VEmhrIXwtJ
egM1NESpGKVeDTvWr8O/E3zqS2XsoPRSdbkMi0P0vxggLxXjtrC8Ck89U0riyiXGCkkuOXn1mpMe
+QKnLLGgz/FF4Ohfx9JcpiyZPVFqg5LNLEUtrm+dSMz0kNPz2q7h+dyighqa39d2PP90ozc0oTlr
q/lurSia7Rid80bACHUKiQ96hgeawnJ2o8NemyqCc2sCYKsbc1mgkFtvEGgmZWxD1z1+AHjzTRac
+Jcq0+MlYB20lZmTfz510llLBbmVu8Ud9MdiASE0bz5vdbV+4nRPSpbwn93hb7R44e4oTiDUGdYL
a3e2855vKFJgfsPtevXUezLVCzVxHK4LjfPeyVxc04YtIZIoh2qNNuqzWEMAFCvETB2lSkLcuA8z
8sNbP0ldgduPL1wQOTV3PYAB6V5lb6iSJKvrpcyUg5r29q8rjbG0stuAOCq6OIG3OD63qZa9OJ3u
oxcUKrBBR+ccz9833XblT/NlAbyN0dvXbTOEh4ACv+HtOnRhQLlvdTpvapZ3I0MSAm8xcV+wHrYz
1hHP3qE0XFbiwG4KcHj/Y4BxfKCPJJ7SAwLuvbwfi4VzMLIsnJRFaFIavEWBZXt3TsfcQVda7cYB
wmrUOM0F9MSEp1gyatNsESQr9qKeAbAlEiS2Fl5hpMsXD9vkv3ppUsWd4JtV6JIU2aTHqlHTz5S8
1SwomgQS6M8cyhKU6b6mkxt3oCMMbHuCtHqHka0870VANkKcHvxLON6h1D8IVR9Jai6suP4g3ZD/
tdICNKRyqXQVRrh0I/A8RMkqbiu+y6amttzkyEd2cm/1+09/C+yHtlPWOp+D6za8F6w+ELQfRjGK
Xx6gHoVxf7tyITee35VA3Ct5e5S3oNfFstF7uVxBWO9Xpkq/+Jrz71YPtBpxdHHO9AhRCp/Eq7/Y
EpKWVdQOpNJfVLb38Z3SsVCPfSVbBEI2hKAMoa/wq5kjNd4eRh2xOYe+QTz8lTHTu5AwE1yYKIFR
2EAv4Acru23SeOAIGMdM4LOhBGAjIQpS5nlKtd9UmbCbB709Rz74ITa/cu4ABMTZtWfMg+936K/r
3V2oqDcCl9BdLQEAWYqc0O9WqByRyEYDieNWtI70KajHJxCQ4AFMDN9FWJHHobIpZsUTBGvo5QVy
LsAsgFe0b2tM49YXklNI1K8EFDzMFBQU5Fg2fo+Sti9TkVLDJFMeEAd1pE0HY147bgfTD/y8M1B2
25VKqdCjTuPwGgMmUGUGAPvoOIjeloBmp6+Oddo5DNd/c/EjYM85/KGvUFauviK8bQhMCn0AIgTq
ADaqG5jUGWMt9hDH0Lm9D3ZYXSRJyeDmouvokWnQuGkiCRPaqmnOZsrhHjeDHAmvvFIFT7bdHwrP
AXaVL5hFUz1UPjm/7AstQNMQtY5O5GpPaTmQrs6ZS9yn1c4mVhSSOD1BnU6dbhq77mOyo0FGPhXr
nt3nWOcQHa6B9z6bFoTWcDPoWpXh68mRhfGChAOBzZlNQMyKTSZoRs4WTPuU6+pvfTlYhNdJuZif
xfhUIRn3hqG8cFOlmOnkiLN53XbSIC+cjmK1nLHtBEGDpG750GOyVFbQGch9SypJuDgdeLMU/mTt
wMnCgFv6f1Ocz0qQTFfQ7EctX2G8SQ9pKs5huFwKWMadVf36Xdg7UyYksiz1seuEBHkZYuB2MP2+
6QziUthj2/ZAUWc8wyNdmd/8BovMDQph/Uz0jDpY5QxLX5qEqmwZYtLfulO93htV8IDJvy6DwfTr
5hMyp2EBx/5+UB21oowKaiTA5rsTVH/MBUhlKVbaln3g47Aa3tnz6kU9Gz4FUmpzpdEMWxPE1jaf
AfMl+DnSqHR/wzfvYxB1C8wvU8dTxvnnawBxS9V/9wceK6i4ywjGCns25NV73ExnMzfO79Wyrie/
+IOGolrv55c4IQeESNoCv2Mq+mH2xrjaNxykVCb8HvHeUez4+Z7JK5XJFkfTWLG9udfz8powrVA0
SdL2jlJI71C7vRS+qvRAMTAznRR3r3Bk3FbHX92qiYTRHwOMg+LxfqTUMTWCCveyOZuKJvFONwlF
Jmq5LoGjR2INa6E53if9DFJHwXSIZLpkoLvw+DQ5NkgIbggVepy5NbQwa74/oRYwu/AbrlQLpQWl
dfwKOnb2emC1vB409PmEE1VyjbQhMdcEOcgyw72Up3EfaPTAhloa7r5Ci0INrlNrqJYVEFLXHTpc
f3/LISlPsTmXVEMlCO9nCNVWlf/QABEJ7bOwv6WtMXg8UHbUtXmwqIZaRK8B+/dGYu+Kn0/H5d+5
qYIlNsScWoHfCtxl1HimGN2qLSpAn2R3DD0lvgECRG8FN/9jGhSyuxE+viFGpFR7BSc81TP1HuYJ
vslUKXS7iiy7e0LsCEOgYg2DPMlE3Lw3xGSCq0r41gHqP8esuO/CNlt+Y6QR5c3bd/pWy1zdiJHc
pWjcwYLfDXdQqq2dpgq8c2Td8W1svSAqQK5W1zHodAbZr0QHTMkhxGq7z3WJ+6oc3NBX1j/DpNFf
89QFIfVDYqct4gzPp/QZAj0cvCUaeMEKHpXFYEwe5qpCfBJ/Nwi3gIgn/T1cOYdFuNsZzqE1b+0l
as2quhbx4iVQW/Jjm0GIqbWE8VdQNznpzN3i5qbF28R0855aw4qSQZ7GveZrQn3YrnvzzgcDWUQm
McOGD98GL3GWPFRjL5Rbwv2N3ToXX3Zl5WHFS+9Q/fHoWgwDdyguuqfjjxtuV9u3NYnNiBR11jvh
W8w1P3wGOrDOPaOhNz2596iGutnM7VAaY1mmywzeFHq++tQmitpiZfXVcv4itn5ms1n1yxeab8d4
1Fkw532cAW2e8gi2besdmT7q4e01xaZMh0iCBHpOhwvRq/5fmfgPKFTxN6Nu9oeI33rlkYXdxX+Q
d2SYs/GKhaAfgdm7ysbL80L+KZcGDxzMg/Vd2rAQZ9jqTzmksDO/XPoK+t2eUZqeze2frrBeyQqn
GuWwLORZphqOk1hROW24AhsaePPxhC4/A/UgeCsgmWuKY7yjzWGjfdQgBclQNgIdVMMoHEPllyJ8
8BSnxEmz+84DupjoEXxAFoz7LLvEzukauQerFRhcJT7tYRFXiM/AkEhjkxUGE9GzFFXmh2yxBC7e
etHBwh8/AaZYk4bo/2qFOhnrkZw3zC3QTSnCCJFeSDlL02eDQOQjnhfEp9i7FSrq6F9EKEXXyZsk
60gfRZXuO3s+kXOAcUu4jKs9uPAxdObXJdaFdBUHF6V9VPqtzMeMu2Wk89omCa923/Ett5cD80T7
Peq4aOIIbPLsBgWljKsVnQDHqMYv/5jyl4DTVi080t0Ibp3OGOOTlRlnJxOkjXPxIuofATE26qV8
PzykkwFuErzebFQ2fTdjm+3UZIC+LB2XiOl5bq53CH56IJsnFxDUcxlaF1EBeEeWcJU99NepJC+Z
clkrOQbzUU572LZFxSlib5kXccNHCh1MCv1dkd8qU4Ib8hfiFZvRGcgYAHD6c/mJNfL7me7HsiTp
5n3lnZmbk31R0WxpXxnjLzriA1AJLb7AwLFbxt1B7Wm77h5qnCLdF8+W/cFq6uuqpo33Sot9/2C7
198BYDe5iX/wWPCH+QAqkWEqjaGIoq6SG4UqrxmaUXbFQiLu3rFkhaniuV3WNUkNcyizTWwLYwJN
FRStd6lVcbvCIN6GobhCMfObRD+/KIUub6K6npOdRC9vKC7AurYS9dCIxj4yQHGZqx6YTMlJ5RzS
UUlQuWzBxtBLySZi19kWiAwyks5V7T31YvMDmKyXIMN13LhxsW/Ka+PGjNpwKq5QYt80Ywuu3ORB
H/LMXQfTRLYhm0OAOgnik26LFtNQl/sxYasPPa7ZprYROCVtoampsM3OMn3ehpQ2ZfL1MCy/FeXD
Ps8W+DM7dQPCFL0hZ38/JP47AHf01J95+5V70WCNHrrvCU1ygLdHuN1Cna7oswqo5wBypBif0GAD
y7AftEVzuLeIL5EeaqxOr9EO1z/GWSV/gtzVmsRoMDT7rgsUWZe/L2Xqefilq9I/JdV0Q0V6Ou4D
+hA5WB6QRIpmPTaq0wPgmHJpIrgnXIjLaKuVh0wzyWGCD/mBuc9jbwMYXNquJHqhK1OghOLvsb4B
bpz4f4CKZfhuqu5b152ltMsdDuyI91hxyKtoUVzOMntzmb4gPmlJ361/xKCR6lD0I8rasJKtp46E
zkZotgyMjux4t4pstRq0Wn+XHgTmSJ30r3P2qPAjz10hlQv47Di8WpwYZ+BOMm8lYaPs7qXYZFKs
kdBjzEYoBhWp9eOk9HyfRviiLt3gRo+VFtRmP3pxZ2krw5CA4FCytHYy7/b1p6SFHce4nVIj3nj5
kMPAl92JC07jcmPsQVMKYGAdvRUwbspE6hFIxm8pZF0cU9O4zq8QuZbHqcrc+tWXGKpJBXceb8SP
MSBZpUuV5XYSvgS4gjlY+v4OZZ0NQGCoU6XfejSZGxhzYh8MAR4Pi2fNrpRhIBySFRLKbanSrooj
6kNgoikp62E7uRtn41bxnmQfSN3ayjxoeiMlw4lRHtfhukccA12yJBNzmorGhDyaf/7xJvdR5Tpj
mfz1meNJqyLNDrMdzwCnvFJyOQNU4S9HUtk1tackAosZ3SkgB/wCkqnmzn+IxtpMq+LsAz6KDImm
1wJIly76zWh63Z67Sm3L6MOLEskEnwdowEyZFwkSLemYn4HOXZCbW2GRZuT9ThVErtlbt6SJmRRc
neB3FhoYAt0aiiGhndDrfwPBBZUSV87/GwAHXX5R0NH+XdVWJGWqrWv3sjcH2rS0LE3CWlxlb0UV
gqMCgAvaqEgfmPqlw9JsAxANeOZ8DxP2qri5z+BMHUBTlm4ZqudGYN8c4OzZb6iUFV3p63nggw2k
NMSvX12dACq+nUdVU4Jo+7QvNdaY3MEQXqurEZJLZq6OidVq/dQO+ujWqqcMZ//4t8NFSX+8tJbj
HXXuqPxONkRbXv0ez3jKDfAb4n9mXN+oSOhCjOwK2qAHCyK03/hb45ut5kFKvqzE5Nw3wQ9NRudh
5mmvJUPTxsxsAcGLWL0jUNBwDQv92hBJxpPTaeTJsSxe0ZUqfCukvfAh8nN6bQk7kvzNPH9KvY+j
tAL1koJhbmfH5vCsuMiw8Ftn67sH+auI8F5WmYIf6rNUMBwGcG9WWAdZAaTg3Z17WGDeGbIMJkGO
xJF88RpwUOFC/T+z2EghzOBkNLBMqNR6uOaMoDk7wGpvCagJj8l0aVTUHZ6VC+Fu3KEXx1krkRmT
gPyh5+3H4VPTksA75EHeTtQ503xgW3uteyt/IhEzls+9Ms5sgkDM9Jm54818dOCfbhv82HCdmAvX
fChixxW0RF0R9n9zfHcnraKVrzfWAaEJYc63rGLfpon5KVKzCIw0rrl7oi4sabKNzr/rgvunD1kW
cnlRIhahZCnZNMClJO7QZHdbiSC5GwW6ndEQiPMjnrNgOZwX3tRTzm9YFAhF2iGVIZbYYhc8bIzD
z+NmkSiyHUKNCbyRX6HjvRTpQOBw6cw8gFgMFP0DKgoGoJAp7gwBceyJeFMqjco+1Cmf66G6jllo
kVGC0hPHD1rUwiEqv8HomuGpTNAhUfYMD4pEkKg8iSyOtQjXGeibg6fR4Ii8n5xtGx2UvZTRRxxj
FvtJDvHPTBZyv5v5DVu/EO5Us1gZZgD+BLxWrvpVzL12koFe1YKkPA+BgGP62V/UPgcvRIj1S9eu
8ivyD5rMWHIASnq674lLuz6c7k+s0vszPuozVVxQTYhJeiPt0bg5VjZlc4UF3Jl/oNP9ESwPD5wU
WGVtNhBkeRWSDbfItdozB8Tn+RhZ+RPUk7C8HdH9E5LBuVE22itbtS05JTmkg+D6EtDOwmd+swjB
GeZDTN5s8/eY+41dyy8e5KPRjkAbpsskVAYVovdLR5YQvDseFhwdTMbxZs2k0cYkQMBJiaCa0Eb4
voVNYZkPq7M2f+xdBiDv3QIBY4OOCB9/wD/hVRn/WKWHjtCBUrQtHxmXJcvqHPNcWlJ+IyyHLcuQ
Kx0XLhgTPKe8H2HcVtXa3+sZoOfz4GhZ70XSnzzy4GP7aPwKDrinx6JykcfwJwO3V+3nxq9JGlBD
UBwUJcEG+llVvXmdSShIXRfxXW5LkpYi0pJHrrLtpzFWDN3JRYPJ/89FW6xS+mKYkqiuGeJNpbjD
Y8CYGReYugVSxz4NQPVWyb4R0l1G0P18x67LwKZr3ycVkWRUsVrmZX5+mpG/K/R3mE9iEiTnz6fQ
hlO3XY+rLxShe7wNo+IQlB1scGZV13ixOipMcDrYaVQfHEdxdHLZsmPoUS/h9z8CGUB/3PmhcMxM
XFwEKpEjaoF/Zi+ZdhSeePTHZ+YV/JxW6lWjkBhil+oqMFicRMKXUq6tkr9KAZCJsYmfhSqnVdNc
bdEXWPnYyUXHCwiRQL5VE4kN9vRse+eqn+icJCUyhQQM3IsrTcSjquzYslrnUVYpxEYp7WLXySg5
zRWRnTdIgITk8pPh58KJTWRPbQnWqR2TQZ/DmdW8oMqO9kQiK2juvfVnvffcdrV2wja1U13WuuK6
hlTL+eH6zYp6igo4ENrwjAp7Bz0Exs6289Hazocut78EQSNNX+GffeIOpCMMwR5daExfYbOFQC+c
WQnWNBarjtB/5OUqLaY0cuMjtqHyrZd91zArdvbcqtoCqpjT7wf3gwf4KeurJ+mfk6Ye4c8uruGa
luvcV8+GhV643fHGCZi8F5LurMkm2cHtV3vtkMBt4Mr/1DibMqOKdWQldr5H/ihJDpo8yLWFYWXH
UsvJacblaN9e86oG0NWcfsQLwV7N2dzxWp2yxyjSinjqQ6W8Z+VlxxyIG4hqDtSlmg4zUH1+XpPZ
6piXqTDdfHuPNRaAHHshqpKh5f2Nemxuabyp543Q+IbKxVkyJDYapGGEqihvrqo0fU5hM6BGFctC
RqxN4RePUSr9/UEdwApMmH4fNjql3JLFtEbep+pJNEOeZGd8RkEjGlQvocGvRyTLRhh3UvYYMHXT
e9OjX6UWnMIylKZZyOKgp4HnKWf3/h5AvU9krzGcBh9qQPt2LgtBSPgWEsZ+D6Srd1D4sshcR4aG
tnnrlQgNybBubvIb9z1dQgCGn2AEn2mw/FoRo0LDZ8zoADHH2W1M6MQ3j6/XMlksCTfy7JdkvJWH
q75Net0c6SQTfkW6hvN3lqoFX3Ge1wSUDQVg/LU5ecBBWWu+/lXno0yT9djTNH384jHkpBDuRtYe
ip3OE+jR7ADE3cmij/an/d71iDjGtVsyb6GaeztjtYKzPu+zL+H/KTmxqBEnR9R6srw4pLwdklyH
oJSdW9unVpRi70KV+iEoLEAsfeyMnUCzo+Pvn/MqeaYlglEqryxxtA2tUho/Y7KWGk4Zu/to7N6F
/TC3/vFQrQN9ydU77rHKPaUertq/Y4dawe+6JVVEMjlk5W0AfbRtoziZD630NHVr6aXkJ1blm8ZJ
Jp/6Boeriu8yLdSmqy7Nr8d1HvdRuQg2s5PCuhPdcBNFaETquz0lWr3V2cl4w+yAqGeHZvgeyxKC
jTNqxP7FYplA02ec9JCs2Npis+cMEg6/AM9gv5zj+Ywcs3Z1T7owsvD0O7g+JgzvwtZtFGWEGl+9
N77hxAAEf3BFo8m3zqqAUTBGW1OP9Zd7belgWXgkktdHjgJPFTrRrPBypjewnRDVGfbx7x0f1jnf
tfgcZPSPWv4LxzYWx4r6Y9H4ugXL7imCnDNKMSwMq5C8TtFi3bpWoVkIRJ5+63K5rYSEfD2csGC7
TiYN88KATzzy+RIBoEZYJoFauLC0unhKQPWxjtQrMe3NCocA+877ZlqZ6jWVlGB+iQhUG89Ad09c
wInRTl+P8pQWFQDlN5wsWcKdqvj3jZkoYy9oCe2UG92YvTpBQr9Koi3AjjJEsrWRRyjP3rgx/Exx
GJT+xT4wMYFug+gTXuwCV+EA+B+cIhW5zLPOFeScEYSYd6X1e6xnZ8b2V6qb9KiUjjEa3+ttekfX
bZE3+dVPzU8ggi32tVwNA9CJz+CBa4J4Llqg7fLEqs3F4WUBt6QFe7hB5EQ2Za7k8L4CdPypiQa9
OgArnCoBOimxZN2JKMa+civehDAz0w9/tsWZsUZpEA2091e9/WKCkkpZQrif8KneLHKd8jawQxKl
irRzaJyhCiFMFaFhBPqTl0lH4z+PFAsbLh/WsTTXh0eYC4H6pBSXMXPU20i+aR8PlG6HhacViySH
YdzI+UCCi9Fc7qmfU2ckCGXCie4TrL/MuX2azJiHRKNNCVvxYgzEVSVO8LdTMn7Lym6wBED2sLLg
+67yoHSFmtjS38kRxo81eK2n5Yvp0w2UkMJvs1lu/LdQqUKzIkUPPX4O8YiakPg42IUcXlJQacsj
O/xlPDyAmNr+qXakOiW3WZx03+6b0NYy1XMt/VVCWtQ/yjnOanA1G8y/YC3pHLojQzPIVFKjnzPl
ZAGFmmU8hDU6QySbtDb+ObxBUpTWZQc5oeQYn3Vrf4AgZ5mUaDLwQNwOfCjOZmsntG9hBUdT2cqd
l2g+G7WSeK6B4mQwiKLiHueh1xyMaav08B7d7WLn5B7bQzOuFMUKvwOGBhmsHK9wdWkToqWal68H
AC1bE6AQp8Zeq2PTYz7mFNp5CFOIkUqgmIXdDGYUguYBOClmTMxds1HmDBfogox85i0newaZw3c1
8Q85GFpuEnWdZpweRDCpygSBI5oO5wTEIlSz0yBszYzF4B3chiJM1T2I7HDJHHegLUgPT4jAIdof
opO9cp9Z2d71tDxB0XUkzwjcYMDlunOLq5AFoVeRKIQher3VBzBelUd8XqzAA3o6Rp8Gemsibisa
3BIIQKP5y9atU025S9tyqtkHDVnVwGYRfydcypK+cFqvH7bg8xhrA5JFzI/ZLhglBVJol8Zhi9+W
XlbOOwQMaKRhPLm1n+K5BgPXmGuFkL59nK8iOHX6ABYLeWX6jI/JKXHmn9ctMnpu0ZthQso3mlaa
931mFDO2iPtEDEEThFbxWegsn4VMOKmmHQ85rm+Btl1kuzAdlfwRphNizk3ccleWK5Ess9y5xaPI
MofuMsWUs3NleHBzDqK0IM/aVNiFiQdW7FqBZeq8plIb+NbFyOb3cndwx/iuM9FfBfpckU50eac4
NmYHwRHNZ46K3CG9iHxG472HnjkAr+XXCg12NbtuGI+91SxZuydmwehTg/VdzuxSeOZynkqjmSU0
iSZ4/Sn+195ero6j/l7YuF5ikEY8kuQby3UeKU9FxBhVn+O/xIajXDfUcC9pm72HqIxRyqf+VdQv
2J9zUKtEs0+MNhW5bGoj4Z8A+TJbX8Xd8HzhCrufkF3L9QorjnQNvxZ/sMptmPWAOL2nU9MQGN5E
au5op1hH9xwXHv29xEF8CoWbx4TCBou0Uwmuk3Qjj6zTrXKSZlFtDnbB7Z6LQT2exM7vmT3DkG59
DnJqeTPol4lHdOBloZ8PEvZd/9AxFGD0YlQU6sp7VtgTt8Fms29zD41fyoZD8SrNo/iFHhmf4JdF
Oa3Y8cuajm9DwsN4tKJ7kkNsMPsndLC4tOm9+oTHLjjpkoXDDRf7tCOyWhs4UDtHkgf/0G744+81
ZD9WpMBn7XWIoiZ8UZ2UmmYFHL9jcO1uuULdBaujkgiL/hGQoavLSAU2G4CY/p5Wu1xSYmFy2J8o
Z0bEM0iRRMxB4egUaTN5TVogzxF0ES4tgd+S58oRj1avtaOGvja8aUw27FG7qG7J4ph5W5D/XLQA
0ArU4Zji0LWkqBIlHeO2kVo/cyKY7cCh9svWhWlDQbD78uDmGzdNuye+Cdb5qGR63xH7Q2uL3UIQ
HHb8OH9XKWpy+yKfvCfXy5cgFkblsnd0uvdj67VYcFpLEJBFxX5tDkj43T3WJ1y5HZ8++DACgYBF
UuRiqMsDKYXBvDKUq591zl0VC00RCf1r7HTbKrOcvMFIK262buAapGUbkRcCr6AZU6AAtiZqj0Mn
fNJh9+aYt4LbBk6WShwsJaYbULCvBDGLb9rZ2dp31rzDbWD8+UZ/kGuti3Xm7XCQMUFvB7dnLClF
rK7ZO22qO5T7+J0kgJ2oMqPFcimKpmwi7gc4vk/zTGDdQ5rdG45MlnC8GfGiDSlO7LYYod0YuHQn
efh4NEr1HfeFGLyKmtU9UWdnX1ObEuGVx7qXoEc2Iclhw9PBhqb2++/zrpjHw4JGM8VhBqRQoEsR
Uv22IVmjdrvAO7FsI3IsqQJC1feuzIsXXw1k6R9a1wy2WYQDvyt0s+kZX/6grxeyOT/wVvMkvR1D
nV1orhPU7kw+tVG0+fcsYdzUMmo3BwH3NUzA7xE84Rh656+GrI9Bqv8dDFEZdzv/S53CjkdgyPMB
JsXwUfz/MHoPIFZGOisTbFotb0cVREow7UBPcsj1MtVANseWChhyXqAuaBKMb8Xhpbfm6Q5ckNF0
hoDoMApDeWeGcQJhpiBz+JLUnf6NuXq8XoD5tPAhV/JIwIy9pImGDA7h/4rPWltFE+w03oJc5Ru8
WV/x4mwZOSsoGh7tHjUnsGT6BEu6pgvMezwH1TeTn4y9idmkgb6b24b56+Ll61CgKHlt6YSxQB9c
Tt0HtHGGqZYyBdDLNI4FujPntQLUrY7a2czA8l2IeheICRdrCqnQGWWASJjI/LgqKviV/ZFr50D7
Xj7oobMH6fCUEmMWDzqzUoJ/UVr9N0tiune7vASFXtbkVpwcZhms7GB2Aegd3y8Jzbu3nTyw/p83
cTj8RPVQw2BRfQsMduM97JmVk2mKFqMr8cc/9O1wGKVzp44okTz64uUA/u1MRVDnYuKSU90KsRgI
kz0UX65iUdeSX2OMqh6ywhOJvbd0IU+BHjKo5B+0luYZy7zPQjUlchzqzNvoUTPvRZDmYvIRskjY
ej/qMVXu5Eqv+15u4AmcpfomoGolid+7vaBoU8ucutO5jHUj86vyfKRUXUFUQ24NZ2bXoPfgc6tS
RIaLUtULMyzplOxzeovk8xf9lTHJG5J4ukiI3ZY4lQBthVRYUOmWCAnNIGoqlns7Re0Sk0YjmcnQ
GLZLGDoeHRiddyO3T7L4r/e1h3MPRQpcripRirBPY3dMu+e5P4/MiDa68pLIccI9sLIHu4EVvHuC
TDRK7vzxmi3GToJGR2lpymYi+HRgenmwjGK8vevKKMYR077GkvvfAhCZFUpvF4z0Izxtehf/R2FE
GwjpwkSgx4Lm0/7s6MUP/3CY3lVehd0iyTXPM6CAMZefjNR2S0oqwiniaIiK6oyW9FTVXPdY5RGC
sa6agd5F8grlYv2TrXFd3j90S2aVXb7WARh6UXbcFfLXb53C7svilhEZ3kpo0o/pHtwarKahvt1t
dQrSVwk/uLZlclFiQxpvodkLFWf89xZRWabun0kAW8LdF+/NtamJs7S8Hixbf2e4XnLROZrvKApI
gBG2x2pYvFsGr7W+fc6bji9mXdS+z/oMOCOJ1+WY1YSdafZ153YTpxJzEMMXhqb9qTv4S6nBPQR3
uR62Zr25cfn6Fhyv392I88OOEZz+EVyVHVwu0WVr/7vP6F3t5VPWFnp6MIvF0y/I3RJBXQ7U95Qm
kGTa1NevHhKWtOwzUzv2aFfS0n+7cIA7oml1AxcWycGxLWzKAp7tLWvgdZrytzw0YMbKQp40F4bI
3Y+VVltUUmJcI3JYawsVlSUR83oIkRaO0NCDIFdETEI0/L0ZQH8lElwbkyCHcXZUhMSSzkfXwSzK
ZRucUQODfszHoo1O1DnO5BlOQWtkwUb+hf+zSMhq81RS8giAmXgRhL4QkSizkL9HBGLCcRmomLm8
nENpsZgL12ue6iI6bSHa1PO76RD/StmVwR7cARLmiHca589KXLKWFwOnZCyZGEi+MuyoAVEu0XOY
QJXvWbNV7tKFnwalzFRkNEEnUUdI0OHj4sWRQw4Ep22LwU4y9rLJwHbE5YdZnvHoqVz88MWDEvFs
+3U1QHaBimHzJrkxHSyCLkLuuC55GE9/8QGpvhaf8qIRiCGq+2nIhcteQ+HFsJfPB9k+Z7idyAFx
SPVvk6sDjxC0wHGLSx2H30n68Z/ZohgE1aim/b1teIh6pncjXRREsYWW/INx46RPpynPLvhCZkNM
4VdWG7Eo5dkuN1mparHuGgO9TQLFrTrxwLG+U+zn8mrpfLcnIC24prGLlh/s5s2BlBK7VxI1HTmD
qr7FMCSfvt8d+CUjV7gL5j41dYbJDOLDMI98/5izPhrRFrFs3P/tlZdVwY1LWknHVzVi1ZPP0qXu
rxZwO7orlgDczjslHY6eWYRR90NxIJaN5EkP/6h2oZtiIZmpSIzfKb75RCRHX96ZPNExCvKIb1St
aH2rHgygHk39+NMVddBK4euBBl8ibpbQOKxq4lmFYVjvNy2NzeS8v9CHyYRrtGNm16WIT21Nc4A2
eBpqgZUaYCPlgAoBCPMozgVn1bwW8emrGji24di+UxdoEerWIu0aQCxT/AfXONj4hIL3Zu6K+60y
EWrSTKBmypGkgAQ1eRpq8ahxGL33KrxgAtRpIPxN363fkEcMcva/L0ja++W07N4D7Hu4ZITLctwq
orBWX0SQKNble6c6a/7F4T8UofB+0AuJXj5BMMGvVKFOUipk7u1oLV+s7hNCe1tMRWZkAhzFuoNr
HGpr5bcDi7gyP9NphKInIu0U06t13Kc/dT//uLBs35uwZn7SN4zEV1hOYGSO6N8/38N3fd0glDqF
ztld1oLl/FVSh64sV0v6WgdyhJ/y/nahyyY4eQjO30h6IuxuXolvQcqn76pa9NY2V9GoZ4fPw/WO
egSV1cL1uBKSP1lRoC1yboOQX5rpVMW+mZ76ikhXiKkWY+rC8/5HIhyuqWFFfzJrZwZh/g56pzz3
G64t5r6a3CFaJdL2uhmgXsh7ih8EJVDRRPzx8+/AQbMbPA2ji7nHhlJbu8wN5Aflieqwh3LplOe1
wO0CItgppkPILLMF7d1OQzYrs6fLN3hFhEjgbG/I3zcnFxdXwaoFvjBOsjUWo4Bq8Z3PgfMJA+4T
MeQ6VIpsGvNf+SKNQFbL4S60GOGgC/EVTtB5V2Bk394ZxZWSsqOnOMu243Gm07POMgvxvpSrVAaL
k/pXETeiR2CH1tiuHI9eHapjMWyj12p0RQfRMWlpCN1Da5g6FuBT5D9Rv06T0YmWcQXUvcihXr5N
JxGrjEctTI9I/Bf3Hq6X4oN04t7CTakA+TNlzzG/r18SMG3wpN0lt6GmcX2L4ayhBXgNO0pfqA1F
z7enEgCqDFYzp+JoeYZaj/kX3kBQSrS94M7Pvas/pa/vaAmPUjWMkyxac+4hg9uJGXfpzVI/maYK
LJsdPWZQyiatCe6ENo8WMBPUV80sCUeG2BU8kLDhA41S9PYFoeP6rZQ9t5ublstHCPojxrkp81Et
k6eVwuXENdFQ9WAOGEnC1ZKfirrfPimWvwnRqcgIT77pf3e27wrhO0ppVz/+nyvXrk3yAbrUZ+im
fGmra/ZLEXWmY8W8whg4+nXGFA4zpshXuuwad/VAGV+4bcPptuoipWvpt0FfoPVB19+n3FFfWZuJ
d52Rax2nYuhgncT08t5f8Ftdx1ZLqORAOGlmhiFJ0pAzQd5CftgsXpWE4K8TC7CEIztTIRcPg/9h
cuabSNswDUrw235x6VtZAp26igkuZTQ4+zQBRqVNmsE2fB+TgX8Ksb5Bp1jpepty5l6tD1grOuRv
dAdiS1tRk93yrmdotNtub6AbU3r/LbEwuPcaXyklFgMI0ZVGxWzbYk2MpsqAhjQ7Z9id0ff72j7Y
uoFT8xl5OvdFVzKR8HQpRBRGeFMKhE8LcutK1cFDbB0YZ3TqKFfQk0WZou9mY5xXFDxBulwy+JMA
5OSi0gXv6G4wniOfU6cIDxXgYMnyZpQToYGu9E5QT8RMTb/qx+8341TkOMAqA06MR/P3B2Ns2bpM
aVwnXo4YvSL2SLqjABluFzjO30QjB2378WZsTU7wA85Q5TbytZe3mEW84o+DmFVm8cTi7QzeGQEw
vlFoPhavGDhokD6J+S4pQWATEx2xXP8u12FjoK1qcSIluf7p594ngRuuBcuMO//j0kEHdCexhF2W
OImHBaEdKDCgugkX5X8UN7afhkfMG3jSSxL/PBFIeNJy8XLJjmnmSBle5g6+db+w1ecueHerfUiB
0kJ0Bp8sKm7lNPYn6Ya0g1HW7RwDqwbtLNzF6tvXZb9RpIPsyLoolXbqD/FpOMyVZlEjhw0HcMtS
6OBNLbeAzUe9lr6t+ziRTt6kQftMo5u7kakbjreEI5j0UjHehp7sRnivA3JKKnV8rFbYPebtRKcV
Wi4Nzei8GDxuKxsPSBqJVdzZw5abP7OB0h15y3XYDWZ/rS3peWfYBkG29M7R4DYKV/gB1mje31cs
5SX8sjSuh9uPVKmg2jHE1anDoZtc/seeBC1mO1/+wOd33PHhgg02gA8kQUH9qn8qZ4XLt6pOMv9X
ZVbiyIct2WmUWmcl+xlQ8QTM89ab4Qql51wpE8M2xzhFqTI4CWz0uhaWTn4F9kqPDb8F0+m/Dir0
d8SlPU1qr6vwvkYCZ+Tx/A6Ouyg3JtPQujqbq+0gyck/MbtNI10h9CvcELYsJmXyuVeUqxpZ0hpk
Rm0vxio8jWiyTo7o1yZSlE8NWusE4ZFlt8m/rffm8Aht/uOhclfYtzZUNSc8ooeTqzKy+PedcBxi
nmyWwDQC4jV1b1FVDNsFeAItZssTcMUgm90HAkTEF0jssLNu0xHja+WNRJwFhRrp7ncbtHyyhV66
cM6RrdROfAcibdsnSzJoDBxwsG4a7hLwFX9018x989RmTJEqsjQPapi5fCp87wtaq7A/Px9tApgk
DOQutO/CwWuZxAmICTbAdgmzhBnjJqkiZNzNL1G3z+0EZEQ4WubvXlPHKcir6bwpMFAmHpPftQPm
1ehxXEd9ZIPHjxIpD7EpbLBaAVTzYS9cX4IgKbU97yR+0VHGPURvCIFSxXSiXbNy49nDdxtXaMCk
JJkTmwfuL3vEbGBwbUqOQi5MoA18Oxr60o/+uw44uzEYVrgDxTA6Mviem3nJCJkjPCGt9Ts32Vvk
dBYxtE5WRmoyedxT2EiI8Z/yd+QkYvgned75OKY39uwX8J5By9KxEO7K9y4Re9inaTZzoNN30Jfn
f1txdvF3mdBPCBqaT4d/CrBvCbTMM8GlN5b0X/cWWgsM5uF0usNWNTF+9Je6mgYOrLL/T/4KmmYU
7THLh0H/0ZWH9AFW0/HHVkkiC8mIlrYnmkbSmsScsG8n1j7Zk3G6HZWVEajKd7YGtC8fs+kjCVwy
0Vq9vgIqkwbprxl+kO0i9NSFBb9Thxz0pypSIgJaIZN3l6Fqaqa2KUgmozFCca806f0pVZJyg/7a
etasx+uUvozLQQjqG1Zu6Fnv1HmqIyN6eXZ0VEqzAjdGBvLGdwkBz7/gR59X6oCNwtw/wtamWU/V
KEeN0q65jjn7Uq/5rwsJDLAkZVnqhsSi1+Rp9kh8IneyN9GB9S/EkdylYg4lAgV8otU5gP+2fknM
LxU8LxpKL/dkjFK5aAM81b2dVKyqCpXZPxTS6ngQA5hn1e9Ix0oJc00UwWyMHZKUG+4F3us16oWi
SNAKLg0wxYjykU4iUr1KtYz+HiJaHFWjXyYY54EvATjowrL3exuMvWkAK3SO7CuHO9L+pCO4fNW2
sbzcllfNwFomd6leMlOqTqTuXVsZQJ7vAVHlTYa+4Mnhz4i9CQfNHDcrY+PiyJITb9ydh2amtPvJ
7LMBFBw/ZFK2Mr54/wZcgh0huuYFHpRYK30efk9T3eDdefsXkcA47B2ORHDOFwn0rOKzWP/EMHYu
Vjq2tYTMRagSXyrFdJwxkHQD0tV4uZmfXH2w7wvOYr/L3oC9fsqjqzb24vpEKqdfgi2R2FY/b1bX
+KFbA4AFEDxiJ1xML4de5cIcl2JIudW9h7I48RPK1vtLxvwfh1lbihjtitmxJEFtcQanf85UebkQ
AdX89MmV7TEZgiF7Y+ddx+nL78CLTAKsOyTSj6lZEO8AusiXu0+9DUfDAw9NPlOD1A7MlcqGvXeU
J4JtMAp97etoZl/qXK+xlIARF+/2P+2hndpb3rJcbh3ctrqZxdC4VywWq8ZYSi6i7N+WaKzHxEzE
YQQ3R62ExmkMxxp3iHxDj4Oc36lPxer5B99IiEBaleDgdlRU4tmjZzdAxqNo7jYuiC3ET2Mw12/U
GOIxD0tTE2fhNSC9fOJUNqkJ7lSAuOENlWWu/qaUWBD/zGrWSbVN2bevg1qe6IwUflsumXzB8J9m
d/xLuYN4Mm9eDB5O+AcrmJH3ZKahYVMcKRa8ZKx6K+9v8qZmdGc3S4zu0+FQv5B8cvIQ1vWLeyT4
VqNRf2gA6sTJpSg5c1/YChDLZuz8CywS1ISPYFFvPQ9c5phDrgGDhEzsabfRQQdm3KXtfBMc5uIH
auZmp5WSd+wVWfBBc6hsfTl+JqNKjak86UHdgwtrQMpxxlOXcK0oOBp73V062Y//38/PVnizGMB1
N12Wbxr4QtWeFcQHqS/vvSe32daLSUFpN2ZmxOif1X8/iqZ+yxePOu2UM3fT8I0UaifGXcQ+/YBB
m0P6fCyuUWsqKNGof+N5KxC93DtNHfWDnyCOXgEAJ07tEAK/+pzPCAtg1l7dxnaQEgsGv7UhtT4a
GZY18EC8rd8eOAlaE8Ohiwe8Uw9zGNF2nKLPXUrLtYvGLtj9jKmt8Fh5AB9+xtMYQ0NoWbL2+sFx
7TLn3ZTPBO7GCAd0J3J0wECThufG1SJxar9A3wFsZSxiKvcyAAoj2m6m9l0mUWc6P1CV5usL7Kdd
AUBQ+wiKBApUTihjzaT/XuLjsv6HjkjAdsAAVCuPZNE35qBlZkj0CETHdAWs9pES2n8m2X5OXsoW
TpWhxC3YXjJjHbV45UvaKNrllyAfIk6XvSFS0qCNqBgr+ohLpYrRh4iPLD9J+KgQ64Xe037OTnpr
p6m9k66VU/eQfxVb0R2a9257XoSPEek9XPzk+Wv0ZVu4t5658N9/7Mb+cKu1PUSEU8RFuVATwwOw
txvWcwQ+o2fy5RE6ASJrfQVtob/yr4DPW0gz97ULOe0irgD9Pil5Gv3doV1ch7OqYtRdYZjPY6hj
UmU6VdH7HkBO4PIYmotCr8Vk45X7YhS1v46HHN3ZP+EUEOReBMmjXyA3xY5CKb4HNEaDS9BOBXWu
Oy2M6zsI8qQDxSRJPEuqtA0JFg5iwCJTKV8CnS/FDeKQXyArsU5rUFW9qZGz4rgCQuNbFfqj1lDL
tQ0BBsR3dg/yyMX4IkA6EynrWQ6fYj0LEaIaJQ/1N9at1BMae0ZwCU7VzJYbdL9uZVegwEm/xNTg
lGVyb5vLAg4OQ/SghMHdBdgTk4jumURcsGBn1oreqYnDcoAcfHF6Oei6KR5LwXDThGI+hNMgA419
q6ZaaTy8h04AxCbwhyUks4ckLS4MaYCDoVJASvyu4xmHJsAYT+nV8rpwM0EKvbeOK7kuqtiysZ1Z
Tjo4/he/5FaprKAvXdWHzjlhCBrT2ADIRG/UBwDvNX01MW1VQ3+bJrjkIhVLLng8hNJgvSUtcqQQ
2I6iywhLLMQa+HAVR+VwR52znvjncDvvb2M6hz23xW8vKXJU2B5t9JrhudEG6/k4ubr4Z13kJpV2
CPhHKAZqdVVNTKGGQHxmmui8U8ELnACde1JM2q5fXadspjzxsbFsgik6mSASBez3qcvp3QRRNYa7
BaF0HyykHccL/gQM4ElhZ1oEcAC7eW85b9MM8dJ4TFNzUZ41Vp6szOMYWdxZS4qH9q/4PSSXGk+Y
/T+Z0mg2jogSctl9gftTBNGzp+lg0YVmsW89YZZmO6OUi5r4M7C2g8jUhUqdk8s1ihcP6cIC9YzH
WAAcqTZUtfGOMp2pnudFkq5Tz5KeYiTTFlQY50SCCJK7dP1QawApO04/IOnM243/s24NYYxywAhu
jQ2RqXfcXfHSkRbnF5ekFJ5FGOcM3QXVZB7SpkbB7ERfMwJYjL/9yhkM1Zf7jmbamLTa68LaI0DH
zpN8jpLC9Aw4NnaZiJcANhkL9PI2lOP9p3Wb0Nr2VOlXOChLfxGK6+FDErlAccVeNoBo72b7jXwn
XrvXtBPMyigkAdupNSQg0eRuhtEbtcBaNK5t0/SgLXHOGew6LV3w+7o1m+IKh+ANZ5fWu4EgItH6
9Mnxa4yJ9xbUucI/deUzUPQNlUBhowSaOK1hqgOeBI1STb4ep75MYBAoDwHJU9ejovXY3EZR9Tec
bVwU7HZ6oUA6/aH530i+1az8whGZwCwq+lJfVmzuntwuWjxJeiYDvduHq60YsklhBAXz3zRzsRsm
12RITj+DzV2Y4oTzkkPRwDsJF+BpiTwSSy+2uwpEMafAwGZlrwfK7XcUErZewsrrExGC7HmvZT7G
8SCzgErYr/R/wHblelLb/ni/lOwCZNHuYpsnIQO6guxtntViP17wCPpxiaid74v/UVEfp0lGeS/M
jMWcc3Y9JHzgoXFogT7BmM30kGtY+T2Dtq6k5exCqGVYcPjLMc7MkIGX2auFZSZwkt9XLQ3DRbGJ
Be3n/+65sedJQNbzFLuarcGas9FhGXYMUUNcHjBom1Hn/w3pf0UdSOFLTMUUXLpBMS855YtmdSDX
YD+c9v/lM4xpbrkYDJgjmh4adqOkjcIy1/f7LJPLmOg8lKlFo4GD7xgnU226fbvoakMgbF+1n0PQ
AHhjZ82CTaEynAc3nbB3jq3hApbNCK3Eb0SVoq7D2mjTDoD38n86A/+A1KMR6KRT0ndb/8Mi0SBe
5RTfM7zZ5xrlAwVFwHK8yGpRWfeJV8I9HcfEmhhUM3jeYz2u8oOTHI3PiuC5QSq4VBnv7WvawlNQ
sWou68+rHz6mpqJ37arsKAITIkw3MrxHKs0nAPEjX+WFb7vHHcxSOk1T9ct3eekQqTorNHlE6Lo5
hPM5PG+lfiWlt78AOpCBZLbaY11DgMAnai24NL8lHuGwqjQL33YsgEOyC9ueyQR65weWJB1tBFoc
iNyW99JpSy9k+fIaiTyloVUyJtFM5cjbExRrroO5uVEFOzvRzaF99fR1krp1wLlmOU6WyUl4iDyn
QatcrHP0sq1X5oZDN3wrRb7eMcZ7zsUdFQtjd9wsewRlS8FVbl1ddXZzYvgEHak6PsSWdK9oTt0y
0DAShLKXkksUilvtThbimyXqUfP+dDOqsqvdQEzsUjr1Lc8yXm9FCvgjparu3I7YaCuAx34iUp0W
MJcV0FObLZNmSGeAGhTBrzobD07XyzQCiCg0pMooMLgPYCEg7VPUZF8aH4Q5y01VBx1/teSEU4Qd
H+xCWoxnLzadV8c+2YGd8wwkgKboqa9SQcMlA+ODGpqWD5P4mmAUX4YhjzDDQEiMyGZmSZV8n9Xn
S+xJ1wl0uOscXYeOJcv7V+gWMd8W/S9WD3zB9kUWYq4tWI2oxdsMRmQ0tSbRnG/ucYsTmpAWOAaH
eb+3N3qNq5aTAS47WJ+GP0NPYa5Lvm37pFPuAmigMcVz1JJbc0+DdfvGwlDDhoO/bZvb7uMpB4id
OBcIArn/Br0Mt+Fmj5Qc7OSXwd7bo4BioxDDxftsJX/8IcaH4gtO+aFofHZ0EWZ8xuaspueztKv7
5heDRbjw5yZ8CV4jVbawig1agUjjfnDZEcWCK9k9xeAgveSlK1gxSj3oAJaP/CjuOVPzw/mJ8PGM
J3kCTsYArAkhkJndqLVzxazM5uRhYxFFmGE8e56ygfDx+Z6F2pncrR0iUxeN3jt5MWgOFtn+FhDH
z8p7EaeCTSXZuVaVW316jEEQNI5GqtZUHYiIhYhP0JgiiT7/zbMmn9dh/FJdcG4xwmy5Vf2cHNx2
6ILrUvp8bms4lFwvekLHBgpFFgDarhsfyx0jQKBslIyRIhOKDbqggLcjN34LRsEwgYUZgkISMEau
/VI8nxpxXLTQA90ZnookJqG53eEtuIGECMVh88Omg1Tt/RzPmOiL2XeTqs5WwYZLs49DBToFwDFT
YLC4y2PKDNgknC1hjxJytVIN7cpGxuE1DTkThVVWB6uYorRdNLVNCR/lUQSbWw/Wzitt5GnZJG3A
Nj2iOoWAhPlrcplGD6mQbg167pGp51fuXIfQ/y8ymvVaef9Oxq6q2LQsOmtJUxIE/DogaNfgz5Rt
P9rKSry5nCGyFzDmYEHk99O7fbVCBSMb2sh0eL44Cfkv9IZVmyr+/8ho6kVpQnoIoDdiROhj3+TM
ZtDzOFAf4YexqpEh2/z7GjAPnxOD6AnEpbBm6zkIDw4s5Pnlj2vPfMOcSz4iRrunXrV1za4gphGi
U/aIxmia0Yscs56NnlnbGby8nk58zTt7U4mBEo4HMhoZ+bdQc4vvpCZdmzUf9p9Uw87oda45xAfF
83SfcNcOwdIW3F7laU5nqrPIz+wCN3GlL4WMJlxddZ5xb2TMzcVvM5dO9uxQGLbKsrD4NFcJaslE
C3poNEHCxBXkgJsrJ5FvFxgEai9P68anm2pGuclLHNRcErWp94+FIjOpS7or/A1MdKD/6oUEvteA
vsSwXI6AZTIkRRwyaRC4js3qwVRnr0ifXXNDE2FUdavqe+TaHSs9xY6fw9QSOxmGz1h0vVDNcQCs
dWrZJ4ODG+AwcnokGSu6tkBQAKiwJLgCH3pf5V2QYkJ0v3wr7jzKcf13FpS3u3BRc/NKOywVMyhO
He/kvQkk6gwkLFR6kPLKTevwPUCax0ClDHPEODWLfsvothcN9vJVAo4qHBQaeCMJj1PxxLZmNyMh
33u9jMHwFXgeoVIP+yMNliN8DY+MPTlWQhKwdw8d2hOUNnGB+KqLGFnHRL4NT9Gol6eCqK6U5Rxx
cs+xj9GMzIcEA+OygHtW23ZHEJF4qUKRig9Ux9QgRhm3cXMlSEing03vKH5/JJcdsCzgWD5OjoRf
QOd3E6M/LQMIHNC5BtKJQrFPhy7S4j9du6+L4paeetpD/szomzandmnczg65VI76Yki9kc6jjnkJ
LDQ+dQrxx5rt3rPLns5SsNA5iWjAnXMXBBJLhDNiwSM4qmA+nPlDNHPyqpXC3YKTJ0dmEHE97LlB
PN7w4FWwXdvQQIrAgGpOkFHvQcQzAgUggv9aU3yPjO/uYOJ0xLsuwqKM0MF54QT1tAVkxL81il1t
Rtf+S2iKU+p8EC4urDS3v+GJZ6KgdpoBW/oaxEO2kxxGhGj88v5SUym1QiwxrpEFmniiMI0J0fwI
UZ+m9BJWYKDReynhfA+ns6YN5wpXKBXAHpCMIv4KFBzxTWRyqm8ZbPt5P9/Aq8JR0zekrHVv5ISn
dIEmnsv4NEGxCROAICJ0Lg8yqN8if/i5nOeRwvNTqiMqblSl7XYD6RfGIbfUzafkwO9BWvWeYua0
BK1zsCHWxiIlpjGpsWaikKycCJhu6V3VcHjQP+U9216R9UEn37xte9r65EaS8Gd2oQVcwL4a8CKU
ZPra2Uve490XKguALbF/YA/pvhlCYClNk6IALTiQiZpaVXAm3Qgwo0Eq9JDZ1yWuFXUSTYViWjN1
GcXBxN4dqTC8rLbhH6/ZHqDYyfY0XuDeu2YO0uCUFgBDjJtEpLm1d3nOd1DaGjlWzLFWg8cqE6CJ
kCt+7TIEzhOEQrbFgtwNLHmMJ/hNuVwFVwWJFwFb0GkH4n1wMkS+R15DP+pUDCABhwhVIqcTVpKU
P94k2s7QfF7JR5wffrq28OoHAgdKFKbebKWpzN7PQRbl685yOibpRDFaN2GYrOVrxD3gGZbNCVNf
P53OzytuwMS1B92vuQbmt0eqbtILHp3k5caSrf0SgX5tSvvTPlqTEBOwUZEB4Sf/sENaQ6j5mqfw
VZMeEZCDt37f4b+Zmdsv6ZyZ1d2UdIpXXgPL6xcQ7KcDKFXRF91D5Y+ddseAGaIdvSrwiEgUh35w
QQStqaeCK3F//itw3GYW1OY1wlipeGcsMvNbIySmd+ncqBLjy/4EILWDaLd8bYnps2vUdzpEfCME
5alIA2RI1YUnmpdfmHKNWUXIa/UTNjse2PYaUlxh0sAirX+b6zuOJDQMXY0graV2jYDMVsOtpNv/
nLC7smdE+gFKI0d1eLtH2r+Gy9UecjadpCRgKWqJ1x5PuwYflfXwGwoJRU75Uz3y/e62CgEwLRvX
xYy7spO9gMQRWS/zj5RGznyneDgxjBFDQ/asYEse4tVoeBcPUR9EOpFO+QP/UeTgTQybi6pQ9vA8
0O860DpkEWG8Ptwc7auePP5dSoCZBdibR7qUMFqtPM1eU6/ROutnBuN5bhCDukkR8rtSnlD4LUWq
F5j8Bwud0T0s3DA88z3xR7j0c0OmNboEFhq52dKDMPDgv6KOtC1QPoLqO3cX3uLfqkPMxDp2O6gR
o+jmn+6Vf/VQYEk0XGQVGJM55o2zS+IPtNnRKZqZwxPMo/V2081VOaFnEnV/68DK42W6tVxKsFuy
fC6p85hh3Xb69QKRCbPOuy6gUnWpgcwPqyi77SVSwGBlAFzwyqjibc384IXWCDSznmKTQ9OxsQ8y
ot1P6yh6SMIP445A/sGQwbLQqLVp53k2HbEO9L2KPKzgqNyVB70ARBpWiEa4KtQSwl4KWYRDisZX
ciPV5woEVtQGf3f7/F4Mamjf2Pf03T7RUeJ9aHdQn1gCeVVaLuxeTSFiUlfBT7XiWFYPewc7D8Eq
LsuxLJqS6ySwqxJJLYUy7pByCn+EpQ2QaDNEljsA6EefgEqO6Ji+bxT9lgtMuQZ1y/1INDkz/eL1
df8+201Wze2MvfCkvV3zJ1LndN7tMsMlwYuhU0n9KTxeYnWkAw1ABdEelSnyc7ENWf+lylhIruUd
1DUIcDYAn2kFURXBrMNoqG25abVxTHevWGA4WB34Dl8hicxk8TuFAj4xhjEByLOomd2Nu3YSfEba
iH8fcxlhMIOndKpcQo/1aptShsI9CX1ZjBqo0+zixutoQH3jylBHPpzF1YDENwODtiJ8wiNv/9vD
kQyAz/Iw22ZgzlACzQ15epYrxiLRSqfGNwKyKim54OdFQrI+maLqqvNczwWmxvgBeSmeiIXc+P1J
4ckk3B5ZYZgTd9LOw8hNV4GHpMz4JiBi8+L8bjvhrAKD7X436qjNqg5I1Qb+PWRPR+poUj6VdsL8
+yIqgfDDRsgY27rKH/axNyNhXTMGAwrx1ks8c7OOffd0UaUUe0IEdkNexjXt3/HDAG1dcZv2oye8
e6clUWcRU7cm7bUBbris+xL4VIS427/8q1UtgtGXjGi7COBSfWopxgQ9B+u4W3T8WlP2+kZvb90g
AbgVZ4X2sms5J9qoNEoly6GlYH+Aws/m3B+GJczNQQGh69yK+BuYA4fF0Qo9lDR5EtFhZKq9SMNm
CzJ9BbGOUgI5SJ+Fyu6I6Mzs0jTGNPI71wFXizTzqiNAH/oMMuPse/ZQOc+SSFFXzCs1cIURMY0P
shW0lyg5y98APcrtPIdIJdv9bHG7DmD1g0Zk9zdfIejVdKsqlPekXYZIK8bwReouCtGGxXKRLx4K
xS9go3NnNzvL8LJIrKXMlVV2wh18XxLaU8+NzEwL8cQbortdRBwQ5EF6642xyYjRjcnTW42nrwug
u/ZBGSmWEdyqdpbb98StXDAq60b/E0UpMsB4/l/DqvKJdOwHpAISzHp+r/fkAHIvPnA2e/g5YKp3
ICykbYnTi01M4eJM8TbQDW2l4ewNmUXyoBnzXDjOp0TLlMYuVbtK6ohOV/X5gdOtuSNNzWZM8e5l
DbxZHOtKcnddw2gIr90StP0qm+2pUxrtRq/Mym+ksb99C9sD55FNFR5hfMZwcKDyJnciCp5lohPj
gYT7lDuc7Q0VDeBmUj90YsfRZW8y87/dqHW4IO1daZsyde0DPrNSa5rxKbW2D/tKI0+i25k3i4T4
S811WMi9cv2kpFoVbgJVuJOrwGWKxzwoSsCjkX/a4Ia9FnzV/sZI0HTA1bfjbDdDBev3GUzVXOPz
VAZw+Iz/zscEvDrbTHuQNWkX0BnMPZgfrXioY/gYZmrCed3B7Kjku4oIKpeAcMATYb96WR/t5ehF
jNeAEuOw4+9674IyvrWLr6W4IYCANDNEyGJg8vlZPGTo/t64gzjF5D3umzCE3p+OclJQAkJ43Ugm
ihlTbc9j/c40RWrOGVHLLZLzXgPuPba0LvmBg8uKiQ0J4KGKWT6Yk+QxkK4TMxgeOOT8Y212mWff
wwAJlkiGBYuzqEhd3wwvJ+npuZoT6tbycluLSQ7JfuOO3rX4eeo/YHDSx4Vlca+7bflhTy71E9CJ
f77fvQ8HCkWk9RoTHPZ5AH+dDQSw0RNIsTVSQqq9FdRa+nK5t/TcADBqpgv89c6qZazQUVXxrnkY
f+KNP1cY62EWmoNFKzELJ4zVC1+lCtqq3cBgLD51NCUu9UWULyPFf6FbmIV03ZWdUn12+0eGumh5
ZLsajtWAAWedzJmIzoDiLogA9nKb0Kc7yvNy0OEhyuSg/CXQ1U7STVwvtl8GsDvj7CJX8kIZLsZN
deSK5WfH09nO08YPsWQDVgi2elsjfjia2GBP9PPHAj2m1FQJwciBhC6mQ+6Kpakhy+zWT340IFve
3EPWGpylZ2Vq0nks2/+2MmauOtN2SiOsO/IxK7s9gBlt1S17r8tqJTKkaBB9URc3ZJDKstL/gzfB
PedIDrpMoh0uqRIHLXGbxK0fxbkcZAbx5pIyjvVxvWm//zjnLzKCmB69lSuYgr3D11FER+1g+4nl
Z902FyMbbcmGqqHiovqEUsBJptUOt4opd4PaucbDh1jh6GYLssZguTGgaO1u7Kyhhf0dbNOyKs6f
CvM3MXPBXNtxWdB4LmWD0JLlS2DcichxTMD2Y3vQUoIM1Ijlzi55ZzHEFkj/CYZd1xhdtCE7kqji
U5vVzf47zH8dFDejqoUVxB36mdfLXLAOgScawGcLBzwKW08H7kxkXPH3d0lXUOiH8leNDjY17biV
XbM3Gn/lVwUbRwGvRoNiF2UH8gf3R3lQRcuyKE3OQzHMEg5YGZhjV82kR59rImgxWu21BHwWPEZy
FpWUmO+OVzA/8dVtOJbhRY0ZhzSus0igR5SDUOoAm0zzZBPpRqxsJEGHxfDz23m4I9eqPPUWv6rp
DoYg0QGp23Rt+5N5PvwZMpsmX5rU53euoJ0kyC6gu598nUElB0yAfkmtFNLbUezoBPXr4VvyTCy5
HSQNAb/yE1G7RpErIr8HHXfKY+GgWEbNZA9+az5fyKVYMaBsOs/uYdeUVPbTwceGkwhvxePPABK2
qrHs3VSnBEJDgY1WJVLBVi4VHVNUMUUJUj2tUmk2ZYDqzCZBH8vy+TWnQ+uuvlEYaudi7eT9E/Ng
PPUW3GpFXnvxKDsz6bkJ/FVWXlBtN2mWxzfWu68yYjwrswhsUc8VErFW25Ow4WdTEc+tB8zKAPmz
pLy+pkWGAPYFyu2sMplBhHS9uRrTin5ObzVZtILOktbovENALX+4rJILZcQwOHIHHo163x3k3BKC
nLdAgIwg234+Mkhd9w56pfLT5BVtGtuN7jufYdTo6Xaulbr+//BSf1Fc9FmetQaQ6WHvIiX8N7nb
AbX6c9j5QvbHII9a15UgdgGjy97m2lGWf9IXZWdOvOEnXNAka2NSKm/B3tRslAuJwawyrQK7a5bG
gRM6vMu6sVatTY28spPAqrh90S145Dcd2bu3ITq9o323yhM/5ghu2HR5PSlqi6fGYPUI+6O8ftxB
XiPuaesuC+bOtp+kZF4GeYjrRNaEekIeFe1nmJRXcgU3Rubpb24US5A06XPi1SSLgs2q+ubsENMt
Fksx/LUQ4ObAKhRhuZnHoVRG7tolYP261K7FnNm5n99iyWzvnp7TC1w2mfh+nrPRq27rr/iPRa/T
xD/LuRv+Sh+wJrlXKXuIgi8Ncrh4+7FVmf5wMpxQlGw1OrdvNRTXea5yJ/SluQ8Ly9zEqwxovdxx
Yl4BhYktM68piV4TaovlhXemVry47LtRaGSYLi3R3wxk2cft/8nz6DVQFPAITCt6N3i1nOJn/56V
F4oVYIPIMMWYET4sgY8EsYz0xeldixL2gfYiz84nQ47bE+QSjM8r0e/cnWZlaiFotCyQfS4QfNP/
/y6sFtl5bE/6Q6lIQKI2phkKvU9ihaaFAZojrp8AOwpTPpAMS+G/4QZovjWfgR5EZkvZlz4qEabP
W1F1eWF1ZXBX47PTpymNugWFNWuUf9vSwCT4t3HerYq24/hi8W2DlYDwNmEAiem4FZgRBM5Vodp5
Uzk4o7/E810b3/2jA/2k+I7ELS8zpqgwxWEO/Q29ge0LTW3HpwOcfMYEVqEbtV7/QGoJJezYCDzU
rdghsXweSEwJcDeYoI92nVz7ZNZS5yaomMXbPGLO16FYnMAQoJwLAm6cIxCcp83+am5RW2pjQzy6
ZAGToQu70yj0BB6WPs0VcPB91+dPH2NyGmndpSF7M4AeMKfmp0CIJvxnzRbTFGENjc5LKbfvaQ6w
TSWvNot1kZXe/AKWj+SUXkdLoCEy9LW96J965qBDLAvQuxKFIo3EKU33zSL+w320nNJbM0UqAi2t
jmyfjlZs5+xzohJXPhdRJWhjTK++Q2Hui1D0vB+0l1gFe5CfRtUILc1GHwvoVWA3K4E+XrXrO9Uo
m2D7Jc2gT/kMqMaGA8y68fRVTUr8iKCCETvu9uoDBqvgUnkHIWvQrTMjrXb4e8ednsw+zAfAR5QB
7CdhF/exVM74TzSPAsGlRqv3vTdGgVaZdRJady7MSaAizfWZnqQeZ/WVpiF6OtHqkTUj8iJ+/Vlm
4C9sKrCogFJOhCqhVsDxkw439lRrp6qgCPk19IIxw8MjCR9Mf7utwYsaeyqHl4//ahkNWQm7JwTE
s56NV6P2PEqJvYhcl9AbRGraVXhURaM2Zrc7W1LKvwT5W5BNVXCIrOv34YJapmPhBQkDZOtqZpt+
B9Q0WYxg50Wl+F1FsLtvIKTAHTtlLMC2quhw8MN7fh25e7nUitd+Y32q6GZx5sda+gK/U7Yw4+pY
T035Cks0qHsoR6WEtX/7UWEnGkJ68zdekyEHJJBJ/nlmoZ8Ncq5pAc2V+msF307x9uLqir2Ik9xu
TmmBbBPpwOfRY1EgtePmETU0SgCXTwsZcu3BqD9tpT7d4k9oD8mrbOl9Ve3tuBvm7+HzWcck+c4Y
dBIBwnnOwLJ4Ob0P46VLW5v2zsNFEt/xKeP09YS9EXPQhBGR+Z9yiFhUatOZQwjz49xqQD9Or9R/
50oLjcnvwCek5uLIyrVFJa+efe5MClWTDip+v/XMdkcR3AliKFI/mfZSJ5/pDCVTSBia4enc/iUF
8MjD+QbUnL+WtNtO+ES10lA8phVcSOBJHt1hJj0pCatzBjx7wPeAEyYLONNniKlJujZvmEG1CNg9
5BD1XvQr8dXEAQ/fwdSF4pFC4k4gAhgrDvH+zDBLAE2iqo+v7Cp6PkwsizC5IA1FbjauSlKx8tqR
NHi65h9of1tY0ljqx4oVPVvNl1TiCly27X6GJqJ2V5TtCo7aqCv9EfPe0TtfaZocsoUS1I0+/2nB
xqL35GanKNJoGnapu5xhvFbooCw6rcLEwlJNZQ4p5Z8Fppi9RZ6TqrTZHl6TaacNWKMblsMJK4ue
ge7sPUIeMsMZ8Fhm4TvkDO0ybhJASX182C0o4lwPJh2HKGcorAJLBkxBYzkznx1mpUjKUwtgRoDw
YUix2h52qx0HRDlwDol4NWsW8/7V30PFDgh91rtRw7LmzB4ze972kHfx3xbAaUKnr8wUh016rM9L
npzogv6SIUeVKYVoNrP1nBUHVgfUe/aetzjRcybHFovXy+vLQWpBER5uFsjsAobL+Dt6PN/3/r9F
I9jPk/jwdf/v8HQndAbXYj31XtT17E0T4Y5ep3xEJICgSOy33ntOQNJ/dDbMMF9+jX/iOrSX95tS
kBkteq76tdrnVuYFGUlNwz3E8z0uWnIYOlMj/ILfR0uGbrm8FVEvZ3o9r89+JnR5eL+Msq58by8k
+dGZ25rYsnJtTRNUCzZ+LWI2SUz9Ow9nzJetEuWY68jI27M03tLdYj9QkBzwRmAHEkVh5SqTVeeU
CG2W1zSSBrT7AjaKRBbXIWof+IFJJAEtVNHJtdJPe+0vRt5qF2jcQt/9JkUbSIs3+vDl+MrzHymT
pyTpYeCWX+KfwLPGsYUNaVlMKf5ZKaUJszcqnzj/Zym+fcBntpsvcHoxTb6DZGCviF92zEuCByUr
9TcH6gafyITFG7/kmakCoYLBsuHuaIJ6D/6/aJ8ddDZgd+VY6t+q5bWwnXdu9Jt5jR4LkFE7hgVA
bZJJNLyuuBKerpljTZl4ZIda5aQVOsrHYl/TX+hLUI2t6ztHMY4qyp5+l9GmzSLgFnb9aQakBE+4
GA5URQ+UBO2djLYmZ7d8CPKOAETQ+8UFrOsIAwEmd2DFJI43hRZfOsAaMniR/9pJCRBV2EUG4exA
FjoRMcnhsK3wn4McYndn2EbHUfb0Q85GvowUe9QrsgVUxirsScyj8IcF8QJvYEinoVOtj0Csrh1+
tQXDVukSVyJ131gLqP5j6CdKTEkGOfiC/5y086sLaaH44r05DKUPlo2fa8KQzpqn06sfdiRj0otd
Kw1No7vIuUp7Zg1q+THRFIIlRARAfHf+rH177QMe4AfPQiXdwO7BcRKM108Fpje44lI6r92kS+Wf
xX03YDwepo5yfxxenZMoEV9Ss6vAhDL5aIKbIq+1MQXDoyRurk+ZGdSJROM+NGICfjauzZdeDUpD
dNRifWBwNAVjZZTuKJCbfcB0cCHUE5H2nSZOmlJbI29ZnILhXWya4EBM2n9MwvthXg4smHACR7hk
ev+2H0ugMYowPKIAuTj/1BdXL4qicR/PKISNuSc8qHEifWtcfhn56EAP9FRU+E8VNPuYFjKcuQMI
44lUIZzxmaxSgCNKyWi4VxxvsyhQGw0MsHEmnYTFRu0mCP0tqnOItgHmoQtEPGbbXTaOJ67NMbEC
MEB+3FqgZRrMDkN80CSKD7QGlWbIs3U29cfXp++R6YW414e2yKLwxI74qb9WczOX6qxx9H92plJb
P/ujSLf51jP58CxT3jYHh9zsnmdukRdAvYFtrSDNcxCGwdGeAPl9hNYtsTXT7WRfNRnTNJ21GYrz
4QaV8h81M9pM2vmyxMsDxy79Dcx4QPWwTaU6Ygn2dSsfcybN+8uheuE41UKZVr8vggymdZb3tdtI
1SqlAASWFnTUzfEHBw8ORvRmPwXk/HK5BPuvD/Fo7yYxGoLUzQay94Vh3sny5AIDUoaOxClJrF5r
e+3cWbrLyESL0NwXw1wctUPKoJKRFa7telFoIPp3Q6iqk0L1IwVStG+TIw01RJCxSUfy1HemymbZ
hPGGAXqNRWq0+h8MLrn/sFdgH06LELiKR2kjiSAWyrQmPVRxjbmZ9WimmaI5YaxVCzVC+aNV4XPk
JK4ek3z2wF6CWOALzQ91X3fprrJ0c6rNGiq4edBpXt0h8G9QHY5lvHhTjU8+Q+XtfK3USEg9zId5
bCmYZGlRCcEjCBaV5BSUckuwGNV1DcXrR7OCs+rnx9Ntmxj81jYeockP/XFSyGLYRcFPmxjktd9l
mvBYyq29f7RZwODusDsErZxJi1SHlD9gOO8V3quK/yOjzni02UUBXn6bADCsPyB9ACd197cBYVoE
Nq4MgksIrh2Jbx+G+9b+eWuFWzZrg42+J4Y2ZRdK/RnnjSqsydTwQHT5bXHAUiP59rzIfJwtnKdv
WlyP8kGwNHTZrn9OfkVXXQc/unH22C4/LytCwN93lcu7JECRMueuiHzuOOoBb/QZ0E3ZY+7cqTKI
sYExDtbryzt84MarxcGPckmt05cvFQGFhj6zgZ5wNd2fsG8GqvoBi6wugM36to8geXdxUNp7SYMC
H2FDfIWaw7NrTFUV3YMGs1SprJ2H+/i6hslfylD9b/SeuAE4aiW05CzPykBf0FOc0ZgQo5Lzdo73
YkxLeTbur2+KEUHxMjoLZwOkTwHHRDYKh5vomjWGRepMinnx2Xow6sqWY0N7H/AYAaXJyLfVg5Wz
/KyPgckA0EKGgSek/ETaxyWWRX/jFe5aB9O3LoshF7C0Ayv4qcy0OayrR+G8u4tRvKbZ+YSioAd9
oSmCuajRMxcCaq0NE79Dcast8gBJesJ7o7lY8Ju60vRy9DlcRS9utKOxoTwRznosslLsA5T9toJU
ie3c505gGeK7v8MyxDW1iGRGg+Uh/kctkgXKzgfG8U/1+YL/L2RJSRTUa8wddVk+K1txk7kLC1Bt
D/K1SURk2KPoJZ0iRlSlQulWQhxLONuDRY4qihGJKI2/jadA64NE1eXC/DcXeAuuklB8NjwV+r3K
ViJhzQnKw1C8RXVT96LPgbD6VBzN2KPGNvHfzuYHtDknbgszVmaAvC8wvZiJG42wDWzriRiUotGn
F46sgioY95fyiMUc2ZLMDZzmlyU/CwxXWG/BpmA/g++/U63dSLzcLeojuYFoTg3xHR1MbVqGtACL
2kiANh6u8+AAlIu0eGvNL+rUFmK9IwdW8FP7mvgtYKJjnFElAdp9Y3tgG/yDmI1j0OMepLnnczLB
l3vM4qE0e3SfuWUl4/SaOCqLStju9cbcyEmhAYEZ45d6B62e8fGbpHah/3Qjpi/rJggkQdp2/Urh
kEqtAJC2YFKuRHWKEKH2KraQojX/SubK509eI686R4hSWNvOykMadT13/hKP2fDlKrS3F7K2dgHE
0CHC5popSzUqJTIqsd5VLj/PkH2GCgo0MUncEEPxRyaIzR6u4sz3uA5yS9ymyzchG3cYz5rmE8Xs
5TdWZ3VOqaORgrtErJn0eVXS1R6ycYYH6DQtorrvUZzGaHrdTSk4XsQQcd07TlEPSZKAT7VUAZUd
DZ/PGX9+GcaWSTNjJuNxzTNb8D9YdzTVXXgPiW0eNPhhd7M1trFvbodFZCq+qXvhj3o1NRnmRaeF
dyu5iRYGIMrtow7tx0r16KeqoJZJS+LlLjJYKj1oN+MfQ+V4n4TFqc2zQmbUJGhxQoNxbUPQdMsn
/TP9BcU7NDypzvpoBlmXsKBzfxUtvcgc0TOCOzHRrZ5Oh/8e2QoxBC6329YsLbA+gfbMZqYRU/GF
0Fle5KwYMs/1lWWOL2VtdNFy/f9vRlfn0liHTFaZqcRNgnx4Qm+IO+XFMT1g3bWW5EWi0zaq2uFM
QyLqgoiZQtJyckSHj25YUVVzHgxC5lcR3TKl9VBGBx6HKjU4rt35jWwLTMf1g7OSX1kLvILeXM7g
l3Wbz6LK/FeiaYtb10jKM/zTmkFOe5vTL+rol6hfwREKEO/pkqDFcMkDw3IDtOVJiGzF4LdruKit
e8a0EETrS9h7WAHhAc98GzGuhpeEVk7EGfUKxMZS6LAaWjy3KRTpbEGigxVfiur6NLC2SwS5cTGo
YHnDvT58HqZp0EfU9kVlPjsdDF1vc40O93XpOkCwFHP1/ubrs+GuSAF2Jm6s5/Oh9k0s8N4HQvh3
x0t1otxpZVX2OS4Zj8wmZU+FOxgXWvt4TRdG0uSXIKAdU6hVybTzcWGpfBiL2AvGcOcJ6jKVfNSX
v2gZWxfdpZemWycEw67SjYCuXhEmUYPUFjYPhCtH34/HhXpyWZ+f45YH7ym/Fwe0amXDSwNlcr+r
PNtbZYWyFFEakkEsGkWKY6epNy4cCSU2nvuvRTL64kvlQK8Rpmof1WEqeNmifd3gEtaYciJZU4gg
yciFRe6vGDmp/JxvyBEW/bsTECnikWco2gfBhi8Tl+EYfcnA1OYkGilptmpNsKfQAARYIhxJWXqc
/ONtSoIDMmh9fl0rogeLU2dfPmol63/Npr7UhiiAcU1T8+nVNfJga2IHBWXx0DJe6NnXzwUgokuU
RoBrwJECI0QrLfT2A9rJ/KI3Q+jcnUT7pbVvBXM4wnl6POCbv0A+T5rJ1aHv0jGOlmmg9JGX5LrP
TSgboRu1wZkxFwQ0/ZSGp+lMvyu9mEFykHA1YtGbauHlPYJgZazIt+vUOdYKSetJ7fePbMniixp0
gjyoJkQ/dV1nlFOgjvqQ6OSg8nfVtroFpKITnmQzJqEwq9LerLPGuPqGdv6agT3I924fJU0kemLk
k9H+mIdqNo/88mtMSwyhb+J14RBn7IhzAgyrQOz/2rjO5FMaX9EptSG61Jjr1eIFtauHJCX04A88
1cWrJABmjZNhx2eVDX7wMOOVyAi+tFv0rGYujJwSzv7IyN7tfGQJQiE3rwe9tAaM+6IqPR2EVXbb
tOvXU7pv1pUxmjR+/uzRUhH3LJlFfZABjCcZJokjvA5fQi4wEBy1IP+g/qDYYhyZWDMJS516scf1
Zk4JB13HtMKehDoY4AeZfCdVUyLSh5idjUNtURiZZfeK1bgCnWZhNmxClabdK/Ma9uhoDAg27nW0
7YJvoCQ+sjtKX6Lq2joMok1n7uPGONTzz59ODhWh+kNM9tsSWPtzU2vuwB5x1ar9YY9M7ddAcaLr
XMmXot1X0vmD1ixpoWMNQJvFteHE/jIw+oqPv8RQYGtVOytz808dYT053KgXwvD3oxD1LfRQXnPe
+d/dZG9pSCfMNKukm8d/jw3xAF0bq15Z+mhcCYT/4CLL8isuiabRKzZOLFnstx6fGlhljUwaB9Jm
ajrQqd6RVgRo2bIVqQJjW5EUUm0AqJJ55jQVzd+46sulPBEO04qS2aQynFeqgDrt+db0UKMCEMae
Lv6JdO/GVmZ7EsQR9SuEwpqdghNrvjGVTnzoV2Ms7k9uBxgtWgyQ2ysXjUbhD4ZJovdkUCkvi9aU
yXLU6yob5nxWRydHA+PbxmsbjPyDV/z1nMOEEfboaUDI4etfrP92fzYTaTKc+JuMqhjxawF4M2ey
AmnSpJwOJSZUCEYKYcCccJlaEhOMUz1gqHzgHLonVuZxgd1pTC1yvgNG/5Lk+9dKVOcws1wHDaRL
DNR7pID74GHIJ4mRy0tDMn0J5h3AknEf0HMqMqlMD1Mpp4PBu4zD36xVDt2SLL5DP0j6mtX6yRPx
mvDvrN0kkoJkh85gd0QmtnMV/G0shVn2FVBcsJ6sBS1cLlgRU3Qd71pWMgdHutO6oPrfodJBGcmi
J8dcH4eSdBw54sW4RQs90Fo89gL0CHQt1TPobmUozKcSR+dPk5RnPvayusva1iySBlRj8V/HrrWV
BI4aSk1uW+5UH+MjpV/ALXXfuEi46+nqKAQe7HhqCtHIkp26WuzW4YzLI4r9vMl9ZhcsL+ZEu3aU
stcL0n9Q04s6xJKnLmobDZP17jWFy5OvSE8Mo1LkowNgmFuOKkAzHJrOM0SPq5snA/qnGbC8RRuS
bTvIAnN0HXDypt4LRVW4+5NWOEbEqnFfn5KyAi8wQ1+xkydqzgOqAx3QpxZvZd+QcS6h6Eiu4aWa
qiXncnEOFJd9KKh+nbnPMiCE1jGbS50nL4sKFO+uQTlf0UaTpHgqXykstJ30W+M9M56ZkZyA9Xun
5fpq4U3Z7EjZ//TdqVT3kyajAgyry40KSuDboRcWryUQD9hihIF1yYdRPvyXXo0JF0zAt5lU7tY3
QERpvgZ0LBaEnzhcIfh02bXcGzCLq6dV2rDoPbZNlUlPQ80/AvA3tUAMeb+0fDjocEtTTBfsXyAA
s00AaDkn9UG6Uj53edFXMTH4lOc6AA/QdK7F2cP0XYaEFlHyiiWJPG76HnvCcevi+t4WwiYaBdGC
LaUiqfLw2d6lmNEkITROkIOmc9BHuaPxWBq0NPZAooDu7A9SGlK44duFaG4TlxhnlOYwKq+06I2b
UKjxYtrlvrOVbWw7M5sfF3nDeDa9kbovxgtZ9q4EOitiznO5pqtfUZok+U7Z3x7HbKrWMYBgyL5V
YZCJGDix/VQZj0bd7XcqeihRCRA16Jo9YFK8BxeVJNpJrFS8NbE0XtLbMhrbawv6ANC36ETn1wax
h3LAfS0Moyac9M8iwQyORqcy8RqCHH+Zk5lMSq5Vs/Vw6PPNP0ClUjNZycaeOxfysxy00yiiMHtr
2HcS6SaUPAovlFig46YklSo1tC2pyhVGIbyWciP6EIXwmuBvB8HAghCbDfR7OJsObT1Ai5tzwNT6
up8ExNXC16bAsXesMnctStxBt/AjY6rqQ43Ghu/+zT2fQ6Y9txc6wmkebmmOm8aN6TR087bgg5+y
aqEdxPxnMatGCHv5BqRKKoVFBa24e1IytCkqDhiaigqq0h0EUyKb5II338EpBBB5602KMdo1cWsk
nd7cd9lSvzI/TlhaARAmfu0/MY752SBuROS0LhVmpdzAfL20pN77BnKOYRRkZ0gv10j77HQmCeVD
cTEww/7ivpGEWWkm+cEOTBzDx6OWiUraTJL59GFCtySmXTZPvwINYpX2dES/TBkRS52m/2kCYGY3
P7bzNCf1qWIOrb3qBfhvc7ZDdb7ZhZ+VBbXuNzZnI88W2ykRnUfFxi3LdJUNGMi0KOG/VjsVSXqc
7JosdlTeatYSYdxnD01RF7c0Q7MCbsumnibc1kq4BPO2jJRfb/1nZHnGKx8jV/3ajuMLJ9GLeFA5
auVpT03VjGLIsTz8cx0FD8vnp6VJjgU2oTzX929bPDJlQee5pk6xv5dL6nBQeE9yfLLGylj6BmMu
xDlE1NncsjpzwIOOfFyVtL4XljnMkvJyq1XfS6v3zkHJ9rnd/V/76rQgga0r/5MOPH1CUMP8J+RG
4ewN8qvCCiBHJZDNhwZLrmaC7nQzXDRzhm49HRr2kG/dEdmOTC42pei6w6EFwTvafkPtOzhphZrq
rB2ROr3NkdbnriNNTZt/TsXlLiOqfY0XVw4YqWTwG/zLwQP+1YXffXI8C8PlMjUEwcUqE6kWES8P
8VYuXNPP3pd9gu+3DEpOgAWqYGBp2/Xeu2oeV2s0uNF8jDuW+0mIOz1NEdvPhUsKD3/2KW7pcj3y
uNsf6kPibLvLB5yOQ4JcWb6lFkFmcduiFyPxfynHIMnlyjA9OHkEjCpJKj+ALMezuvoL9bBis1Ui
Mw/3v3lCT71d5sfTqETRyHfjAc1vFo87/yPzW81CwSOWVvQOIp1dnzzaOpC9Aq9hHqUul/ce2rRs
ZoURgfuipekYKvBw9PAEAf6Y6h9z3sx+HgkB7LF1t5PHa74gk4dbeiTUJ1p1CoBicJH1PrE05f8H
7dXQUgWAwfI8kiBVak4J8yD3GwksSUiz2LsWNQKXA29tsM4ZE1BTa9tNlRHfffYcaexDoEmo12hb
KrV81RE6dtRTTpHA2/n9WvBq5YrDdiSBcozcBACk3vZLPmVnXKIo9dzbEafblV4Yz/TvFgaHt6SW
dn7uxMvnaXTMHhAkhipd81bb16gBYaxAuSCs8hCIgBy+D4axbac7l2wCurhv7+8VLeelTLP2eYzD
e0Hz3gjvzwCBlu2FS7iI8TrOLTgpNnBzPFsdPnGZNALMAB0apYiX721GLjOw8wDDmwY12NZxRNdl
rP3MbSP367VaH7CazWaMsv6jtuUFi5pDvXidMIWRolmNvaIZJ9iRjvh+6D4RyGlyyvqiSevdEJLf
+thGKaI/+KeNIRFByoT9axacstOZAkqkgEm8/oQC266j5SpuSd7cJOwvqnqBrjdvpicDHu3h9ZvL
5HmN/bLQi/dnr1uibI2lu3byChbUrfG6nlnt6sofyW4kmpVZWoyMIKm/D9zZu6BUTATig6qYojk+
yIO6ZQTPTHtOCAbm39E6rzbo+MvvDOofnr+b8I8hRFjJucLeWbC3KMpmyB/JZlmfDtkT69rxcTtm
Nw3iE6sF22Uhufr16OA8XIvTKj6WR63fBva3BTuX8OjrMXlsRBqZmzElTGBqK5ebc/2IZF8ZUXOn
+bze4kCnz6fA7EZcTxdQ3pa4giGc4TrJirYkGlZtg2efvUWN5Dgv59+tuPL+wIwK+7TukdvfdyE5
YR8iyPUB+nEx5lxKo2x8xC+TRuz2SiyGxiJUmExq640kK+u43OTUL5rAFqp3X794e59ggvU1Y2VV
KdM8AOMQH6qpfDGGsGqXYqssHGfxXZcUS6DPPzDuaXohL5QfbpuGsNMGa1spfSXxeLkTCqGelsd3
1BCYEbDvkkTqYT+0+qlsmw797NH6ChJnfcwDGWFcgRC9doJpYqfpNW4GGD0OCngIh54rZy+9aq4S
ykuNaMWDWC6YB29MsllVuEE7w0GKMDSvJz549PbLFGYvVs4IkjZQakhGTL4kIbYH8tCzT28HM4Fn
R0jiqfUIfKCB8YilAoqbG5QpFFmTLlUvHAkTiSFXzdsDCgDJHQWQZDRSFqq7dTQhv1b8+0gqB66c
uX3tZs/Y4glj3lLBdKc+8vlSPWIBUR+8u7nGG+3AWK/nIQqai1MBIS4SB0efD23ewTNN8A8wEYC2
tUZzscF1wJMj20mNUzehCiZQyJmSlHPY/NpalbSGxGJvXiVYO/dHZBBj8JdBGtbLYaP1ArPaWjoh
sqskd0cw2kjsVVSZD9jWT/pjADR9f0FfuKI7QX7K1+n0rNsR6tBwTzxJ9L9YE8mZqykLDHKhC8Jn
4APkzShFk2Tu9kWg8D4zSVqUI3rAstA4D0ngBwTTknGqxBg6CKsRv2paRu0paP9elbgccYJdEElg
1D4s5DV8Zjx1FiekWN3zTWkK17qp5SoFx3Pja5kpiemEfLPKqyc3+m99NuSElxNSqlmyhYNH5ypD
eHA/b0Je1dTt/0Ue1fwieLHMNXxE/+hQCQdrjV7PQbiWxFlvNiWuhQjRElrsAH+Ql+I2nAd8YHwR
J3NlN5PmI/t2KwzaF8lku9N/mGNByZxhzHPnv2lQDatCOWWpibjWf4AEAtTbwTcIyZpmqXUwUDoB
aWjDRfGUQpyjOTIBFPBeDnmV4pMoV9CbUXkI1Kp5YTOgb3tgWnRHzdQUqsS/YAa6AZoZBubZ+chi
LwLxuub7xlkujKq/8cL4wZvREtZC18IfNHT9RsjsIQh6FBRgq/84eo18zuvOvqFiw8+VseXDIGrH
wc9eJWRwz3Dxf8pRNSBr87XncEq7GDDUS9HUynMHmlTdPgGkIpmAm0mBaYVOF402ZqCkM5GSddxN
3dXz9It82dPvM1SBhQRtcjGownPR3dIqrmNLuUx4BPBMan9I4Jnje7QQkp/WUb7AQ74jb9L5Er2n
wOlFLJBAlC+tZPF/ChPY+mqncqVvPXarayZZ+rQ6IC0Pfl5Viq3M1uovoxRBQ9YN3dOiZnwu3223
Ecuu1lPY4tZhfW2/P0FCpwteHVurYzoRR0EP6RmP/vDMPSVHcrDPd/GUMLxg9YNGwSc48jQgqhH+
ZCSHUKEAE8VErbecjSpGmJbujf1AUuWLY0sd43Rx1T/RB99z9HrpvRKE/W+O2Ggp+bR56QKR2BQT
gTh6mOJ32WaXOAIGSaZpfiu1Rga9zzL0eMKtTQkVK6Qx1vrM1LpHokGCUCMNTYyzd/J2Gq5Vermh
FzJVXv3mzcFiyG4LYvDtwtoQYPjhCTlA515dBfPR6jHFn/39Wc+8PQFygSqUQv9t4+VK1sQ4J7Ly
T7fhXLvkz0eb0GvBtR8GuWMmI+GKooGH1LYkttUzZd+f1n6+w8VBh9epGUTC7hdl5y9L5KteRrnE
zm4hKuCEjXAVUEdZJe6HJbqAjs+sG2atniHJErSm+8jks42GUvFpI0o+UL6suHEX0ey22pI13J9h
WdxdyxBpkrrfyXOwI8Pt7smM0Cxh/H/tnvQoUCBr+zqnkxSSYLHZyuOH3YkRkXk11N0jDZOGJSwR
plBoasMdztz1vNxUiBzAgpM39/slLKT2Uhfqji5oHOC7vS5oITCxhgnXHCrE6Cw8Fb529NM2QKhp
Jg9Fwj0QctgOl2Bu4la5XXrPVDtk9iuOw/eeHZW45BCxNSCW+AYduEXxfDnzvkF/xbyMH/GzbUJ1
ZF6Mzwfmzgwq2H5vWh9WMYhoXdqc9+d/zdcwUu7wvAgbB4eRIDQ97KZbhLRQnWX3MHCyhrhUoDJv
O56yHMyFPiXVIgKZ+7OUoPrgZMoufbeW6G9qNOGFNaDTNy6G5Tjh1OORc+b85ajyn5v6OVKIWTAO
YIMuVLZJsQeAg8qhBrbEnexMBcfPXdrHDdsiA4O0Y2j2JLruDCqaQB318hXvolxQWAYXsbGUqwfO
HWaOksulEh9N/qQrOw+2chnopv4CCgxX9AOJAdVMZGlxFL8GRei5cpAC11ilFRprqKB+eBPzlX3M
JRR/+mTbLofjeQuH8yxDSWY+UCDW0U0N5/ug9wQA6r0Cc/YTimOggExLAM5LaOVouqvsTt+RiZj2
oIa3KLehgRY6VOMavAzIWINVE87jc41YlKGWGaFOJ3CeXmR18HmVyUrZ5hQhe7iOj/GBAThzivIZ
25nnkcX8P/kq0ul4AQkGSWD5qPM13HtmRepLmIf6eGvJttF8tDAI3bfcWBw5KQrN+WKmYkdJxPa9
7dHnZbVlNipQu9PPaLRLXosriE97RwonzFHvdtU8Eof72BNnROI7uxyrvwFHkm8c/8X8V323xi0m
Afo6S+KuMMWQUFJ+HokTtuZ2QTii+oYl2c34xEC3m0cAge73n6srNuyimKelz/YIyyMJwoZAfATv
tSpweyJSXpJG1hOXcZISD5FEbWrULP/DdwZ5d6tVR4cRmBx0bRJS3YmgQC7nosI/073yef9Kj6Dk
Q0uQS4ajEivjoS5wFtlBasJv9jv7VsCW13SxBDcZaiy5iPLHZW0jRvhdZ9eXdzUQLO99zBCxBOA4
k6TwTb20wfnjYFUqPiMp4oul82CFsHIuxmdiWedshHNegtVEw/GHbNm8bs2IfNys3yqXSaxjGXfz
l3eqmSDK8PhXDODPevM5Sbb7l4DyafF/umFeijL8NWu2thuEa1qb480b8w1o2mv4zzd0OcGslUdl
rEjvYKKKNRabN/nAAefaQS2pAcll8XQOHOr4AnM2N4i9qZcmrea0qcx6bMErB/G+rhSiA2W8soIi
24XspwOwd2ZwXYkgw4QJWlwa6T/ozoAF6BCSzMRKA9oV0zzU5YVJ1bmj8LA9m8JWaFi/s8sEkT8j
u0t4sOc01/rFciC/qhDCsmWDndlt4ZFZjsxFnBzsCKWSXOLaqo6s5pDB/tCLa93Pc4QcvoNlUuUr
LqXm6XPTk4FF80CdvGZZgb61slJR3NOxGS2KPW1l4jj4AxZWYAh6SzSYjITrgZhEyMhqOB2i09wr
9G41b7LjyUfOBrUlu2IiWaRe1SqPswtRY3pX+h/omzfrvKiPBvUbtHbjSwAVondvIgD0Jcy4uOfe
SmhkQETVnfZIYVthad8R9EOWW2moGB7KCkzgEO0IA+UyF6KE9ocQ9YafaTsnA2pCkqhwnrsIO4YE
HDAyFtR7gcdEEOtZeus3rdgswSIqtlF8kZpkhDFzKN3CFZVhmUr2YKS5nN9T5upWCopOd28kFXnO
E+7DNF2c62OUNyp7YRiC/eUAGKgXtufVKbw/8A2qbkR+O3qmwH1n3qgNz4ENxWJ2Jg7pwWpwMA0E
FQLFPXMUX4ZZYwk/8UkRjwp7oi6UeyuaQxzewmNZRGYExY8tlUWAz2LybfiLiWG+QDr0T0jgQF2t
Y5PAwc42tdK+T/Ch3Yd577qaYVfT9u132ZpbAsG4jW68WR5wksZKso3kGHQZLl0J6SEh5sQZjzdd
rFj+XzvQ5C8s+c4nRSKKuajdGsW+pg5oRdU0omVqeHaLBNV7HuT7Y8OoM57WHRtHcqov2WsXvhs5
9LpVYSRqeq1nhmeV2wlMplkJmRSJsmwRbtAdkJ5So6w4YwFz8RiF+QTjqa5lfjenT5Aj6W3ybJVt
O/MRstsOmpP8xMNKXdpzjrq107MI3i11xVKCE2osDSLkSaBuf8w3BoP+mcBQ/8RJIFtgFq6qkIMA
26lvvwqmhGAVSQ8YLhK7yB0CVX+CCgClpgakIMetNbu4RxRleZr8rlCPArBoWpscwXVHvlzc+tBA
e6fa3UZT6BPPPwGnsxxBg03zORWRxGwIOACW39rbeKj/P2oSDQmFd7TWeFnSZ7GD95c/34okar0d
avIY02M+4GSfz97jsjrWJ1vQVMX/y1b7pRO7YgXYOR14+D/lxTZcAts8xSOnk0wNbOECUkQ9CJrX
ONKuQomjW7TfzmioXWdLuPXXigjmfe5OJFxDEq/dREIWvAyCemO5hpWraveChX5W7cxMqZxoIB6u
jms1gRm3aBxTggNaxkqeG9BPab4yOydKZth3G40xffFnw9I97GNGZ4mmRgJhaCb8dmaimVcrerI8
50c8D0561aNOtYAr9xzq5yplox/PAD2fUep0P/dm0skW/KGBH2lGnEhZ9iA3jk0zNLq2WMhS37US
HM4eG0yXW2TzbtyyjR/c+k7cs7X2HoXZ1JkvyYZODC4l/GUIueTZK6fhR+fsgDDruzBAd9aGyL2/
ZDKQKXIZoaRVazNfdd3gAqv6F2Xjme9aOAUvTu3ssfvsmwO+Q+sZ18G74ucsXeZVJrTBligT+6uE
I3/gviIf4xQQNgGhGSl4VEE+glAvs+s90xlBsNzpD3Gz1GDL1q0mNhxFiF5uTanoVeBRVzxd8TzJ
NMiI+5AwUSZOJxBmlqjvxS5mQ+FmRl3pKbffhUwj0rV9+ysN2g9MyrGzo+HMPDHzQBqHAc8W3poZ
8uZ1mgDUS7LVcHk+fMVaL4idDfFVYOzInq2piwLRh6VZjGqPCaMVMuT4vh7Wn/aTZz4wIGRXm2Er
uyfM6Lbbs16Bh9r37dwEUVgrKMCYGoWfXHHRnMhfh+sGYK+WDS15g+UP1Ba2vOIFcZ5XA7Dum6Jj
FRsCWLnVknZMspwKgQCfQnUF7bVXo83wJCAKvebtjSE2T6WXCsK4yr63G142CHhKDMMJjceem1Jk
p8ZFZX34IK+uEKDDw2ZAxokNvbolK3bF1t/HaU1lDFLmr8l/32Sz6sb5Qx/FW6nMyW+dDsAg8Guk
k6cNRoQwFjVN4cU1ktn+l/XufyUHERnU0h9tYe76JLP5kt5B+qLKMZqekmqfX1UbBjjPbVpmJiw7
35EmuTbRPvERDzI5DiFLiYXMwQowKh4s2/RRGct3eHvKIGdZQp7hc/ROx09dFkEjz3T/H1/qWKqO
oJAo6GUQMIAbrpk1QePIXBXpzf7JDcPVynTbheZaJYTI+X+r33Y8Rbelj62eny+AMLF4PFTGBMWH
zepuMmA2oUlZkkkaFA80paPKYyhjEjNFs8lNj1iL4u7QX+E1JwgJe8TCUUHWJIZQs3DFYPUxdlsi
GPLkCHx1TOMNjQq8kwrdQF7O6D/jDefAmYOngTjvUC9udnRF6glOWvxIVPXpF31m/2dhK9Cp/ess
CLMpTA7+YFKMqFrsGqZWx57SbdfAF/z3kYXmYOMfoLl3VV9RVVmbnl9NIX/TiI+hFzIgJ8nPTuL8
pGIq7KCUkxfxdyu4d00ShUKfQ9E9rQ3buZYLQK09S3rCcnrCimEW9CUcb7wa7Txhv4ga1QZnyVzv
8IV7GUsSykBKlZ4dT+uWQTAOnehT/BSMUCkm0FrdSGndBdq5i4vWTTIbwe30td5LeT9/qCXahcZp
ku2MGD8J5q1HCOwxNQIeqN9ndbSWcRB/cZKapUMtk1jeoDoHsgJE+SvhJ/UHVfbHmQGVtiQH6Mh/
IJr6zxnYHtU2cUSpNBACd9/XPiFiNT4OYM2J5SqzQ/+1Ef1q1Wx7FWzIMH/2/+L56zULjKViixyX
Rj1KMua1oH5dLvNVimH0ok80eyt8VX56gzJE5XJA7ElMaSMke0paV7auLaCrWVKIYsxGQJV5Z75j
UEVwHs0Zr0nQvr/kywgIpQVGbyLfrLFlmgsTyzRQWfLkIJ9BZ/F8QdudCdJdnEulWmto1qbUDHCt
vSmom6GWsfCUeEEtQwGWfgxx4wmhuJ7F+YU1FP+CqVXaStqxkT6yLPoarT9iY+TAGStiFprFF/Ju
qcm3jMi8EU3a4agWuw61G4usiqekl/82sQkvj4XjBGoQbO5bbjkpdOBN8lQJ7NV3HsDIwhL9UxVW
5aEpAyGFOdmNg7396u575fz8hmD5MlmbghNGzNCKVh6D6ppktVhVuxz3cJJa7gS049oMSO0KRe4q
0hfKnmCxtztyG3EySKruvOewuB9SlOktoZJhLMOP5osZXJV3APyATznXntADGQ/djH8v2HajJ9Yh
6XCbkEofzJQJ9ngHeLeGXnDa8+awGqpIrB2zZCYgR5LAdOdIwnp77XnoGIvpzCe7hq/xWu4ePCVa
OQQ4+GVdc6naKnBfYT4FDWy9BYtILM51Sy9jclW77lM6EFwjWGQQvCAeRBDefeZI0H0LOfaNLKfU
ZyCrWQMTUNOJC6Hre681kNN3PG4o6Rtq9SE1CECnaXGpPSi5RlA4raVteVxiyViDqajEzYJUUbvZ
ApBIyJxnIbQVww4wWTqCCroVLLtfBoiIzsjaPW6Q/jZJiuOSmUBggqeIvEu2hNzP4a11jtwGZ9wS
KfDZc7RGl/HeRBzGj94wKiTvdx4TZrb+xwU+mpMQrBocEYm1pX+8uB+tlxFCfJPfP4UkEebXK4a+
9H4kAWQ6dRzwv7Al4+xrwMssyQjKhvG9Ug2i01peTVegfmHuv32Fz99nx8rSjLDQnE18DEL2dr0R
AMdGuww3v2HHhaPjwZFiy6VcAi0OsWJkKeDs3h6z41rQ9AxhOUikrlxcos8LaEtFLdbeKg1F9Rgv
sRBbFqoxd0KUY3Cv9lYTfsiS5dPvV8jrWsmkTZ5P4n2j0CKd37+4ML/jATI32DN5rFLWCV4ie3LG
l6OKIB/Nxzo4G96V+mVVNGAmHSyfQvWcOyNzo39nSy4BVutNruH/4sqLsAjwaiLp1C2w/8yWbXII
6GKNgBkiJ+Lo1HAl0d0KSr5YsJBob3H3u2WgaizegJ4xUbtOOiau62MRgMa/DDH92DIcty+TPTBz
Jad34YZgkrV9wVZ89R7U5Lw6qCc50aVC5GeDZ+YxABjq4ms9ql2LljasI1pdDBfThDbJhCwEg0V+
d7k86NYoSd6aY/FqOqBX2VxGByLMR3Vv4Yr5kyphX3vpa1Fx8P4FJz3PprYyTfltHk10iN5h/5fs
LSHgTgf8IMZTLQGapqrszJjT6WH3EmcrXS/9QHgXmtaa5oIjVcp54k4wxRoIARRp+6R1vglDbeyc
7lR3EQriX4NJu0A+yidweBQHFVzv0D5m3KTiJuvxTPo67QxwP/Is4KD5ePlliRj9Qka74ckfBjzf
oNvQEABbBDuphBAm8Q0nxTfddQqVmkxHphbyHoNWF2gKo9j+6tASuUn6B+Jze00TWdx+mXtTm/Ko
LWcb+8y+cx0GnkrqkyJd2YZVedXTnyBMDbh92MR08tYMQLr7eanUkc39a4RqVXeH5Xt+Q3LA6A1i
wNUWj7uGjfImxqBZWpG/Dbxc3rIZXQzLEwiaNoWqvm+LQfk00ePoqvxoX/PFdvLPuxf4fxLvXC1y
zsWI4j//9J3VHvXerc7EG//Rj5jy0fjK3ouZ97th1+v3boFNx8aY0/tf3QtPaOcysRwWHWQWwBRm
N+l/gbou+U5xdav7EdHWP/Zd/Hie4/sCc+mc2RJNDBwHPErQS7Su6mj6+VjhUrje3kOteQdBtF0U
tHV4sYqEiQXLuVxV7RhbDxJA2q/P0bYFjCRhdka1xsoFpuNG+LwUtSJ5KV9mJ+3Udqf6FiepkwxQ
+SX8CKdEp9kIG69giU9UofHecaD8LMAcyzd/V2OafbS1w6Ov+mL8Bifv7Hz/q7JO3c15J2rsv6C5
c44ZJKViSRZ6pJWnV5i70xXtcxtK1QXPn3Rd2VGh9iluIzQ1DYPEy3K00fOwNbeSmMSPtLDDa0Nt
+7e9fUEs3wlGNdEi9QzqudazAifLe0ehR31KVLcR0tWh5EJq3UYu9D1DegrqP7a4mXauTTisWokQ
uPkH6sb1CAi8dhBI5YNUSHv6uZBNEqrHuVDvsD/SotOQaehuttrJ4yXJBnufqe5YY654Fbx841ZK
Xmx84etwYaqatIkCEKA++3D81hZ4tuBWcZRPfp+MVY6oi38C9p+TE88Uub601JGqsOo13y98DzSp
ZDheTucBkgwsMTmamU1oZV6BN7jS4gkKo7GFsLPOHBaHUJvTwCXX22MOaw6hvVtzgCOtmDZcSCMe
CmYrEOFMa30Z4b0Viy1h6q4PzYR0R4RGwKNX4QGD8ANe18sTZhyMe7JUvtqfln6Hl5zWqwzXVwP9
owzRg4g7VQF2BtDINBwratCPIwg5cXof4ezMGpXRiDW3ty3EXkNIEAsa4k5XVHFzJ4V6K8KQZfoQ
wGVhRKGHX5kiDVE/AjWw/11h5L7t4DjjDqUCBZ0SDgDUe4pZ+SpRIf1lkKWSQPpp6vS74RRD3sOS
/JkFsGTx2gUlQPFqBw500wUL/ZS32Lu/c1sCrwveIX4MNdQK3q0ykngh+PxWP7QarySWXdblUC3g
EvhT+pwiU1uHtzl7wqSNpw3lp+MIPhq566tC33roo7c9NZS6k2BjEHCdEZa9RWlvO8ahpX47UCsT
+JfalAnoe/urZf5hJx7r2ka6mxh45BuyYbHMTH+Rpgr9cRIOaiM+PtflMs3g+StMGWQiIKE80mqA
6HB80mClXYLDzt2jlmPGt6VOJcM+VtCGXDsAve9tgcNIw+Tm83lXUnhs2LolIrJoeO0YAEBzm5bs
SJjkzvScbMc5oJM+WKwMTUYnVs5IVNHv3ncZ2udqnGyuGmk2GRH/rJ4eEQ9UI7406QTzVmR3sEcs
2cKqvfMdoHqjkVNZhqw700CMXig2n9WO550hgqqQJ6rL9GqyW/sL/xwt85UYsEx2uIwoXXSL/3WA
hPIkhoYeX4caSW19PjHo1fAZkrdl3JQhP+CyEJPYkVsI8ybLmDY+lHKsbZokTUT4tqzEzQS0iSja
pKC/fC4zBBhiElOXxflzzYmrzyLaPQwTVM0Xx9jIeQlRgVsCUFYpTcdoE1CuM9WXruGfhWKwC/9L
7zxjV0OLbryH58nFwo0tkdCxWL8C2PR/kfAzT1AeUMgnaDoFY3H08Tpk3bb4I3ZDqirSM4M5J8FV
Dxs9PRrga/cmH54eZXUB5Fw7RRvwCYARChmjdkA2V64jRWXksfvvb05upWJaaQGv68R+Me4pGLL5
dBXcJaUOYeeTZpDdbMKc3BOBErTEYJ2lcLxQ/f6C/TszPHwc2UO58Ea5arjVMkhQPOkBTHblsEXG
PusNLvP0F69CAljSg5tFv2aLmuYdBkgoYDX0m9z3ZtiBKZKptA9WXHosN6rDXYXsG2+PT8kKVmnn
Rp1/5qhuQUvJEwK3FCO9uBoVGu8BpmMJZGKB4AGBO77Plf254y6pIDl6hcjb0MJIlVoxVM7Z4J6M
KSrHNUTdctTVBo395wVSIDU7Pk7wizmL9ar24dilLyn2erVwEUAURYS59+F+W3+hOzyz30bE2NKP
kJgJvKI0GU+6Aa49UyS8onLFhijR4jvgFKccOjWLY8fE5jBN2heMSovsco1Zc3yTtvwk3IeeJty8
4F6/pBc3L+FFiSlIek8F/OsAV91NrFuxdZfxTxsL/dCLC7cXpy6HIIQULKDETD2lOiIjcZmagIJb
XOQDnr31CsuHn/y9P8A0JjC2ilvEHSKEHkTPwTyjxAJBCOoIBqoGkFTZNhk1oatrnTbNSXDNFW/M
UObAnnGTSvuEWEWz2Fz3jCM4x4tVV5LGBOm2ABsAyyr+6uJ/FodztjP4ndOvakPXzTwkNN9/+uJY
XKkzBjDHel2o6wAAnhB4sjycPVw/xcS/zNJ5lYaVLzDGAL5ybfb4x3S+h0dV4CGB7INoFStEkquW
3Sq0hAlUWLIYdWnJOfR5HHzEiBQY7dgt3PRoQ8a9t87AKTvcnuPy0sxipKTpDwG2MG+VncKmYGHL
7IH1rMrnwSDceBYXbtl5vPjIiadClOUxGHVAiANVMiSOoE7lvCOL6Cb2q3eg5erO1sytq5VCDLKv
iWnJvB6GWvhcinsdLZm5j8xoplzJS7zhbAQiiC1kZ3ccoGoiWjO6lco5fQdJoAqn9iAFEUOqQxbU
HJt+Z/Hzfi1Xvkoqqn6KYXrXvKwpa/O/FhW2p1RiDx2nesMWtOzeNq9ROboKZs3MIEVHM9EaDeKd
hmZZzW69Gji4xZIijaQ7DxhMr8BlhfrIRX90uOgBB4qZDDtPqof6bovS0XbJ5A9c8NijmKFr5ldf
lh3GVCtNX6GnA/DGIWgDT0Nl+ovcs2wWvPvj+PTSqYCxkGZ7f515Db0D/g8hvR/3u4pmm0DGKrud
kCyUyUGHzlLZ4nI/wWHGnM9Md2nkyqvfb4lI7QkDc8ZYZu0QJQss+6h0KTV0oZKjdmYsPCrHb19l
l9hZvgeNr7W5K+QuZwVdTo1+BOzVUXGcASvgfng4b8fAyfT8LF/oEgDmVgH101KlXGVGECyqhylV
qgqRWIQF40u+fJRYDceKaz9QTvk645kKK724VvrQP55cPm7ZSpo2vV8rzbxyFIvHzIaPw5qEQ6ld
xV7QfS8RECZE+9u76a25xgGDwgv+dePvMQNJ+XagHKiop4EKN8BPm9gnNgPiH4ClLAYsRuQ1+IIf
rktozfTmC7FTR0QRbZ6TpSRL3nQ5Q5GSScWbNriCDZLu1dj1KJoB4lNBldSBhAnK3Lrat06fw3I5
wx4KTbKSRke6k7Ztu/UbAvGy4E9oS+lfebsE8xTSmZlfG6+D1xoGr+fas5hfdOhADgZPCYMZyYuQ
mZuQ2jSb+BNFuDgV8+NUnKd7r3cD/0eiGwWI+Y5TupjKzkZFzMNV33FlU4ofGM3tQ+RycvZEN40R
NBZdhyFrQuti/y5S5o/uYmyO55xn9MI51qudlQQQoE18La44pffcIr1eL2u/4e/L2x9Xptk/Sxma
6fqQfY+LIvKx7/nT1eRYUwPYANj/k33gDyO/GGZHzKeL2JnDXYoeqeCdB4rdh+s2NuFwu1Nl9bE9
E5VWLlJPfIaS2KwH0inINvTs0f3Zz5bJlhnyWct2zG8fwztIRiInhHGlb95/k8PMTOeKlenGF8g1
+8CrdG64+vtTd8kmiQVxdLhTEHgmYvVCRRAwTMKU+z99kQ0+UKmF4LIskvbOk0TkO4daeexjOoZD
E5nUo/0hexFtEOl8T13PdX+a5PCP1oZpjVopScG9aGg0L1SxAtZKMdWSP1HJmBcNbleO0xR62KMm
1lJQtuk41isntGzK/60nxe6vXoIT+FhMW9eCQZTaaCC+xqqaoAUDsydjVpzqiSwZhThCOb5OIthC
5dqf1rfi+V/UZBxd4roGqt3bKfcCO+J47i6qNA1lEpf/m+Jvw+mC8h1rEcsBK6X/X9stO7l0NKZu
xbKeumJxDnCS930xTlQ0oqrkvEEtaM57vs4IF4RGBJV8HqpoiacoaZ5AheE1N6IoXmzHuEM9hRka
ArvCjSUHBocX/wlYjUok3G8L449yArMos0D9jCs6LHXWxNyrKLYuJWhUVsQe3A8Z0Me8onDnuIro
0kzMcLIBhxggsFYd0F/LJepCNlpdauTX24a0AFVxOJbtBU4dR3AW5mQnWnfzZoK6diCfUNY6pf+9
vopNHeIYhHw8LfyoQ+CcUPOGUZg9/QMusNlU1QM6W6TObhGXNwVplqZK1mkthPnL6G7RhspoHFmj
Qb0WvvRADSMtTwFONKhCrnLx+LwgX3nFSSkfETDAQzc2hAidFqR+JEXgPtIvLHmn5a164cioYEzT
KxElUXYi5FpK6QSdRAazVnjC065E5yFyj10TYUk+GGh336w6fB0eBZsfFAFVb3GEFDrWiLykEtEy
LQsmBbBKLwh5HZiFY2KbClQcbSD7+YOnBplRNVLCIrji26h4H+dGoruS5Ds59Mhfo0R/A5lak2h7
ggYEd/AO1cv3M/jIMNgIvWDkrcPTCahZzix8ysSQbhADrpXf7irgkgBwUvoccstRdY3s0YDWxpIv
bQuvovJdINB00ckjy7/YFUu54WjagpxAPKX4C9zM1UhYNRU60S2ORwHx996RSy21ztggdPwqMhWm
T+l952TJSE5R4mB0nbJNS03i5BxJlf+tNISc2ZCJgTY2f/wKmu4oO1y3Vwr5+eZDCZgtGQhwi2rU
N3u0U78Aco3CVPFrpR/tTU4vkZkzw4Ij8UllfJmsVDls/g0HUXTq3l9L2ctVlcWVPRthJgvpnZNl
J2JCb3h4U13jdpXV3wfBIwbrqbpQV4xfPHOkyR/P+HqbSMRp3dhf3qaittTp9BtTxkb5wLJifO7U
bgk8Spsj6MyDeDCfTHQpuS73inLoELpWDk9FnRPIpwJPlE5Z7Fa0CLd+BC6ro0Z08clTUpfU3zb4
VmvBsVpaplxgL3Z3ToFN5LJ2ly/tKqwdJiBf0ToqtfuCnT9+k0tTBQ2r0SiKWC8v4czCs0FyjNg6
UlNCgSO2aWzHOEJmRXny39hW6xiKbvAn57VJhidMLEVE+yjWdPdZkMvhdEQf5FbSN1/txtp99lSW
zoeHnpfymKt/ry93joQJ9pOIlGriOeDSjJW1gNi+1Vjajk7FwAuPqnY8cl3gsJIYE5o7liBwG1Re
lSTf2j0q6DEl6xi8I6yI5IVikkQ7vQrP96AddzNba3Uu6h1dWFFs4FMJCV4/MvBIldD8uM76Y6qp
EwUbYnvOMW9iw+7FXNzdnrY5xSRQI4vtF7UqeUow6yQnUU5EQllgF9D4NdhWu2tqvUamesIKDW8T
uFfGq0a5irwikK56fbO9FM0Hrqv4634GPfL5dRPSEWflnv+nidJ57lRaQnHXfqSF5eJX3+j8Z6yu
D8fGm6G3DOFtPmpnPeh9kXekHqza7HQNeioag5MSnSBC6VmnjvIWXJJ4voFoehekcVROsQqXWZtT
8hxHJO0WvTHkiJjTPPXZ73n2ng9OFBWPEGgJf7kxiBUKdjV/mvb68zvsdKCvIP3SXHkVtjoNrD6Q
EOlHJ2wqoD+zz1ccgXrRMv84Bd06EItQf1u3aJdVb1dcRnS9r2GIO43g4x6q/NefiWZgkdhxf+lD
IKPS4TCj1tE1+2EkNkOoenCfKtQFgTPNM3bzJWxsZTZLyVOpQvEqpdC2eK51S/23GDpHaHv3yWmm
Sn2UlFfUpsWffFtpS46BkF4tqioyol6ZAWPLV/XlPWfJXU6o3WbddURwhuuVBwrrkzvOoJt6/zqb
l8QvM97V0H0ckFpqk8O4T0DlkNFx+BaLUtfBzEw/JCinSwM61d1bL0wyK43wjLlsSRxDXknJLk+t
XB+/qBcwEu1aixs18HEzSbF15MPjAjB5b1AHwliZDcJJlhNHvfsLzBIjCVqsTPp5HNMJHs2DJlP0
QUTt7NNXy+2Yjh9ZfxzhAeaQ4Er7BWg5dE/rFdKLCVv330OR0USFqs3f4qGfDrto0oJ/t+7pXEKd
8z4MnZyrpGbWWk4uJonlkZqUFa7gVB+sYMSkAmwNkBkg/1G9B+8wxIBqy4XiEVJJc2zlK6RSEh4T
yrTzL12r6lZjf9MGogxRfu7piUjTph8HLMcsCI/ITBHNhCM1r/9uilXcZHw8NQ9GdXtMGKwCN+OX
Dis/Ik0o4lu10Fp7nyN5Q//hi8UfUoKoIyz8Ng63uQPt4nAo587LJHhCib6C2CRXnyYqKK2FAdwG
8vbRJlR3I7z0y05VJd2gKYHCAlAgH7iBd/vvXDNw7g9FH0cWR4U/nbS3m5od/e85yYRpXOQ7/gyJ
/rXy5KdcoMpAcmIe1PU4LioOPosUnla8SA0cb7De8DjH9Jsi/TyXbM3ErEAroCkw5uID50lmChl7
i+zHbHEEQb+IqroHKhA43bKcac6S/p3/Ps9i5Qmh4iELBUgoaVJIkFuf2ogr/XVHPzPS6L79/qsH
zKWFPUqo6rIeeygenn6iEbqbQSJTayyvE2pnBih7imy89ePZ/jiye2OT3+PW+wILTMfujipJK3Qk
ouYB4bpUEVghbvm4CG7D6u+09rKBiFutd/wd8g9sz6gEL8txrnQImKEOWfMiMTYeItv7xNuurLzz
TfpsLL/jBwpWYsOAFiNDQyaRwoAnH+2NRRDNWeskeKtatgHn8X+PFfaHzJVjhL27gaU5EXI6TIRC
fwyOUlQteTQYUI+k4AuVSrdsW7yF/Vy+/TbaUM6fcDoXvsqHAkgK5kULDdQlclJMxtSiOqB7MOyl
+b10H9Ztq1TFz6AId8ZXdRO6M+NhzZjUOJWJtqUbay98UnKx5Blps0VS7shD3fTwQCHECrKZcMYN
NhrFZusp+F2fL5f6yWlxgCVpRZ375H0x3Ghswg0uKpW5NP6s6p2z2exGQT5yoF3K7BVFFzN1bgu6
msYYrUbi/2rgMwiZ2xrK/xM28UOtlx4c1dTf0ou3568olkAhkUxX3CallqNL+4QLFTl4SvY5f/Nx
gsWk+sugnFGx/+sTWNYR0FfMXM6ba5LSO9ZXpQb3ug77KJym6ZogdrmBWVO0Tiqzh1usi1RDsV4f
OYozj0ErZJTRbQ4Ua50mzMXKsJ11tPqGluoijkwqlmyKYawOLIPm5OCeQFwCAz2tEF7clSRJNTn4
8tCucQWBRSrfoy99o0cAKTGnjKkbza/BTa6OO08Yao6hVVSKg2LoaMI8+DSv3J4KvRAbudoz4iUz
DgCrS3ixL4NVftCyModuZ3Bkvw4gV7DD0/u+FjJlME6PvzCZdbvSd3iWG/Q0PaZNDz0qSSC+Lf0+
w+s2S1yq7QwXksclGFYSw55kobmDFyVCioLMpxiBIzL/yo7r9pQwm8Xe6uuRbNzsfZwPECTvIFUH
egxq/CFrPbGs6TZs08leOICkR+3oo+FAWbEL0ki5GOz/nnIQMgz9gXfIPQKGUidImwbpKX3QlSWh
csAa1Y4KUX4xXXgkZSiplry0NBWPsw47yMHKMcDQ6k7/nx4pHrYt+egiEMEScqVmESSMu8PJWkU8
/5wZSEdUZAJWsbVe1RFvRueDm6+E0VSdq5pnxP1lZljbwAYLrM0piIfoLsM5FsSfI4mO5hbQa3ja
6jGs60Y35mdv58kgzqdE4HOBY4sHKBD+OepoFOXjvP1h9KF6U34h1JGAUIOxpz8ab5E5PgYwaUkb
w38k+zX3P1T5WtwpcadGFUinfYZT9e8n+k2vkiayv0AGrr0biuWGf8zeD06p04osLz5gl1xPr9e+
hgYCz+xxsqGWMCGvP9WpTufpn6aPu16wzi9Y6u1BCYt75KLYfdz9wZ6ml4ABAOqNIH9rs6r8OiSj
8V6mqgbY9jAmccK2ZposRIRc/Jtg4BYmRBEO8MmQtecEoeg7yIlMroaQTIgXFuCxsTh38vesau9e
QpZpUSbCrD8hqptmExfJXGUay4RPbtJVXgki+uXps5u4lEHvIf6LvT/n7uKU/pxf8u3COZUhYkY9
sCwW6/uE5u4wP0id/oIjveASFeXD4T18d52HyzsL0lZkcPFCVZ5rv+UwCop7rEF9PZRtmC0e+ng3
Mzzias0wNHhT7niN8vnpHA615KyGTP0nH1059G9VeyXRUek6IgaXvFuLxQe12+tt91+AJ5PPRJy3
FMpgBYXPPZ+A3gqTjhjERUKQA0CWAY0HBW5+oxHi6G9FHGy/yrDSnTPzLbDZm2OEMuO9AE5jkpJJ
jZwD7JpYZQAbAQe1aUydhTFv/dIyC0olYpEvyQdOJq1NP4qQplKX/3LXT6gDoOll+xxuZHKuGuFN
d5iQOsRjplmlO93fP24usV7y24VdVnknSrfQ759BRzKXHZq7PKn7tqEXF5NQeUHMfl5NRs2O97oR
u3rn2c7A5qfrjJOJR6VYcK4SZJ87m0RrG9cY4EG7BlfLWgydw0ZzN8MmZFPZjyJ4R3+TkziKWrUy
TKdblSxsPtdfMnrkguPNWBWhsqlyc96iTQiME5/fEOJUBbacoODuqajbbWtFkVW+TlYdB3/yiYx2
p1PR7aO5E9Mo8p21ua/3/7pZ/tnBbme7n7cKpLv1Cd/m4b4Ly2B6BrTRmFkgWtdzWdw6aTxakxh4
XpfB1JElMjeekqRt9cGRSlY7mncZyGCeEW+AQA2AgIxX6DdgzP3yNFo0h1jferlEmxtkUnV8JyHy
d0kIIbVWvvznJti4GsPbrijjbOJAAkPUhHknTVi7UPwKb9+VR2QUehlCoif0re+m+QMsWl4tdq+V
SLo9lxKnhsHwMkM0pnIondYolQUOUsx0bXGUIl1oSTJ26wwBkPylcTspYdzykjLNTb6LFwcIfqHx
4bh3b7E7Z4T5w+X75lSx6i0Dv66gckdQO6sQ4aqQVhOid7dt2fEWQcrfZLxHI2/Ix37IaM9X/5j3
bhuZ1JgyBR3OhzjQVobDW3iLYxV18WsiK9MwCO1uClmfCcT5MREjw4Q+nNxjxFumKMfmgkjHSRU9
7A56uYSRuGHFrxkJPH10saFbI8Cl9uLot+pU3kcSm8F2YCr7dJip14PmFjBr3rOtUc/aTciEzZap
zNSg3BErCcmg8CWML4DNLHYHgWE2IrafVa9til+IW04+5T7KAB2q2YgqR/nslE1K4/L/JyW8v+EQ
fM2V6R2WcPQodxkkJZ4CMu73h+iRhiEDrADryUD09JHppRL9gascuZ582lTn3SAW/8TKXKG9xt4V
oPqZl88VVQO5lITCOG3S3omr0ai6khSK/TSQ4Z4CWSy6Ji6abFJDWjaZIsQkcUShURFl98I50f+R
YI2YaIlnRQsmXzDCyglOLAaGJ3yeu6+rXzJGqb2OZ0UNybGw28wRxkcRPCGFs0wdsMa1HiQiBzgv
BrObsQGOAJn4yj3P3jlgt+FaM0oLz6wf6ocfnZhCR89qLXh1Xruhlmeop9suUUVeS5heYwwIexOx
8nvzdMvbgDEw6l3ibF2KsrnfOu2fABVdX5cVY6vbtzD0+K6/C/IwTm3zqAB0eaaF2SE7C8NOau5i
JMX6G7fzr7oHBhDeeitCg0TU7B9QJ3Rm2tY6rthKRG7elGOs2NB/CtoQ5/9M/G9gP/Y0LTKHjSjb
YayPkuXwiJkMdSth/7gbTBRBvGTli90EO+4N3dTzDXs8m6lgjCI4UGo1uWDq6iTzwzFTS59DkRxA
9GYH9ownDosVWdgB5+FcLvP7z2xQweIVmUx+Mou9AkSKIlWMu2km+uCI0ZcmKnYwpEJRyUTAGPTV
WXgsNfpfFS9Ygi6rBXTsawY4S3VMTj6C12+CTuWiFlSbJ6BjdMjZm2eQtZVaIyu0aqqLWasOxvmR
6ZZ5p5p8gET3HxczMfVu2YXQbUF8Kh5O5KFZ5mNoZ1sPs2YUF+1rIxzNr8EjhlPNket35MEPPLjy
xT8e/NaGUnmGYl3MUyC8yn5hOWzOVPfsM2sma/gRcxbh8gE2z+xleSvIWasUil80Uh6io455PQ8y
JlgC0c5yXUk+oTzkFBcEssTDfWG/Qcn2CvXyBDDBDpEpxI2YQEhQ6I6kd+jrkAY7etvn69ZcwLHh
gBwUtKERfGlDlW8636tRsN4v/MD0APBJalkwBL6w1uDiMexj7S/rWgU1Bd24Fylt4Y6yayMQS/BQ
gq31NnqcbRPKEITA7n3gAK29LgqnN0sQkzMKhwnpfi8xech5YSGg/aLeN1x5r/znYJyey+kRoGd3
ld1IxMlP7xb1Km6ZpXjdRdxizdvAeHiOAb1wf21mNgrC2B9u9Wgju7OAw2VpySUBeJ9pDjgQqIeJ
WCQ5zFZZ25pGFxFn0ZB6UxTp+rhT/d3d/R2skHoYiHyU2Zh9AUqeDAV0ozK4DSVcKZ3mhyswLF6I
szgn9snJ9ftKamq74TvQYg2VPeOJ76/cx0qXGqSNMAZ32Cs5TEa4ZoNdab9qHwvwpgakjg1nMWUd
aWixjZIHWMw/BPbarHO2IeHAWNKvjc4COn/fb3mWKjQe8MRjBkoNROY4nFzrQ8Vuf/NaVRQY0p3C
uN1dI0XXvxN3Mhj2PGMVwj38KD6atTsQVXdbvpKNjq7eg8z3fi8k7Zo8xO+iWyrAiWOX16dAlwXk
9dKZB4exld7Jp0JLvQ/llI0QZma4G62u/I8J3sIRNluiQw8rDDdA/e5tw2l5RcPlx2gKnavpq8x5
257ng+AEwud8MG67lhz39tVMw5a7kwx1i1zDCZTGz/ONpG/DqCy07Dcz3Kd/SlZfP0SHX1eF/IKi
YwZo9VE3GAAzSfw5JobwogyJShsQZ/Ns2PuNsNG0/nyIzh4lRqan3NB7dOUlodEfdrwTNOBGFiLy
ejsnbScq4OxzngLLDB7NRUy1sFaThA4WsRtpro1ZMaXtPGaKGcSb6F7+bD+r2e3DUB/YLtXpxTV6
XgJs+crvYTrFZh+iFjQWi5KJW0+rQ6WyZejK/hFsmLfGpKf0N7dLjXflOy7pnNPJrxyit9gVZmnm
mhEyCjseqXnSwHVv3iTL8GVq2Eqo2iDstV/VOZYmDtY/Ch0Or6loBhRwIVqQQxxbuDLHx21jLYlG
0EoxqM4OTgrgC5yx4Ndoc99CmVDAWl2UZLGPg7lkawgyHHKep2qrCxHn1lyhESUJtQPgqftpPlDr
y2XGtpkBEXkfeGhn2Vfkqz0UmxZdmrbEdiYz4lKC53kRXemGCTf0QdQoEuUe3O2UDjSgyRGMC9TU
4wa0sLVse4TtARfNl5EByqVzZI4R5U2j7YcZkSdGnEuG9lQsqq5JB+njyw3XW9Og5CWu/WafJI9o
6qa3Ah+FzE08n+0PNNPd2hXz0zAYKrVVs2bOQ6dw797Ra7qNySmUh12KxEuGRy86ajNpkyG9mS8k
FUGtzmuNxcW1dGMU6H03ERxKQsHiCM8V1QKk+F37a/V84t2CRLtgysAKShk3QTRVcezH3FAsYran
ENrq7ihyAtMmAqw4J+iGLY3DDzh1iUqX46ZITnPqx4l9dERbw/AoBS9Pf4y+DCH4Fls0ad8d48up
V4E2+5K5nB23B1z4BK0IXNmanqfi1moGMZ1Km6UlXY25gYQBV+R4p+rj6Egnrk1Ws7BHfGWAhznO
qMFEg5aBtYUun5rAiAJW8FRyyHwVgzcQ9FCuSDIvEWfNmR8Zqx6exk58eaF7zopek2hdhSRJNB73
bpDkauIZQn9jwMXSkdfDxfutgUunJk4z7XAdBVLrOdZVkJOJwe1GvRrmpnN4q1IsgP8QW8Y2Zqfr
MpFEvQQc5rICFvW5s7jLj5duBBch92l3s5hyKqJheylV904kH8NT8Czy/4n1RhnYA9NC3kD498jE
g/stip0TY/tKx3wjThdXCXNwFa4MNy3Fb17St1MvOxRhRbrtFLnNabCPhdaf+Vc4GxXWWoIp2vEH
g/u3hNiGPTpKEF1lNTTIsSacZ8Sm7BRNj8lSyQ3p32Z8mifgmmq9HBFCr4uXe0jIKMgs1Ik834QT
GjSz9EsaTe7fWoTtnFMwgkzZjuAKNCCeRisGzn4lozV7nuScR3cjw5fVzGDP7RF9qA4tjHiMdAco
YhcImoiO9xKUOGE0b6ftwFcMaaSP1hgaUOc2telHJEBv/kRy3eQOGBLhkoqRJ+6RyAd6cMMrFM8C
wHf94Jv66Lw8zQ14w4YvtGE0D1qwfZZYlwzbZKdZNiGpat0JjXzP4XXEkk6ypYPsFaX6+81licC0
bxQSBKpn+qUuUIW1f9FFu2ZSGqq7HSQUGfC2wuWH7y5aJUtyOn9pyJ3N+BUYUhJdi7tdvOYMpPU0
1gwRfynf5gs94UYO9TU8D8Um+bn7RCqyEKlS75iNYloN1kY2CjLFrZWNXZlfhyjZHPydmy/DG3Yf
ORuX6OyhNQp6DaAoBrcYTnA3heGa6tsx1ne+8/vfTIo3ulPw/kf7lmkssR6ozMZo9iG9cyQd+4Ky
6MVJDkEWb5uPVij0Tb5puDEWZnfa+2Gh/wkdvO8T4kHiehNRNaKJOWrYFrx9tuSTLnK7/eY9jyuL
cnxuFBaAp1uVv5z3v3NprIOsQMhfDryUIG6LptIp4duHz3/EpFp2cNY1QXCSFdSolZfDjIvCxBkm
PmsWJPialWxhL6RcG/o7I5m0bpyJoGGHVecKVHagT9PhI2yLUcoZq8ahOaQEILroxNXqr4z8QUqf
6E82KX2sNDwh9Mxgapgz+ZDwWkkdxrcrGs76mA575KzB0FulOveBzvldh6MI7ExzT5LhfUKXesi5
cDwraG99LPI6t0VKLBmKx6GPZiV5saNsS7qgnfqEBToHWLnukUD5FCVKrzuWuKKuL7QFhfwEusem
7ZV8u8rRvSVRR+9d7keo6theMRSTT0qpxp4iT0LM+EmHT8DBGmDAz/rHULtWHD1nhHVfj2fX8vSV
2vJJYFPh25+G3qcW8nPwLNrdZWHLF1GoDd4m301x9K7L/xZror9VxxQJ3I4HJ1bdF6FFPsOLwZYZ
giKaPTnv52LZ1adqSdxxdbdSqZRt1X9hQEfa4UWc+OdP3BMHw64RBrrTuI64VGnS45zngsIIgSEh
3mCziaEu450HTM4mXHfkYJORt2AbwglG3sD8Ypo7glkZSuQbRrICk8+UVT4ctuw8YPVKdN+EVnwh
Fzkr9qR+5K2Ssyf+B3EMP9Z5W5bDngnnBw2zA3UzVxmcp4YPvvo1SsD41yZUPhw0Ak9VOUqCoSvA
Tz2BeTTGurM9Db8UWBcNrBIo5aXZIE4pUOB++ZJYDqe6Ll6JYqTd7zYTr/fWcVe9g5R5hDVGPLFJ
1gTosX0WxcuhleoPRvWf8b8pq1ipT8OBQx3mFOUPopdYOCq/5i57/I8YIbvxUdZibpukh02ze9fQ
GfnQx8L6QzDZ++vtFAU1xprM/l+m/GTooCI5eHkkmkU1pwdG4PvlRLYYpJ7iSQM7uMPNCF7sJgiz
GxpylfFOW8ABdJzNaMV8I9QQEcJZP42rtTSpQsUN45LkrtJ9t0dSYTHfsiSL2Tl8uT88mvMSBvKC
VtYY294//F3VMvYvmBDBv/5Oi9rCQqRdkLed9cZC03AG9C8+6Sel57AZFtwWEPr90f9HKYuVFE9N
gJDTkOMTh0wy22Dg5vv7VLRgN6bFdzUfpdC2pLoIFAKj7mxZiGHCGEYQFTvPw1FcFUkUt0PrcsRp
FwtnruYgaTZuShskrwpA1WwyHMT4nbXPcZy0jVTms65jHPEEt36X2ZzGtVDgrWBUcFKJ6sSTmdBd
9MpP+dOVHV186BVHLK4CgNojmJSqO1I23f22e2pMc69x/E11nk/lXiGq/MK4plNdjsviT3JGA6EW
6WX0F9j78hhkZiLFBgPynwgKUkiP7crTeYYwQCSTKgf0vfwryZLu9+7QXvakoQIps471XD6fiZkZ
eoAGpDiS6sEFk3qiSYCAQhJ6f4i6HrTwxJ4Frn7UF2QpYSJYOMIlHnvkENV2KySv+16xIYaLlNKW
WdDk0OxFgB3C3C3vNqjWOuH4T8h+pkOjQPEVwjvuZEJTuZPxRHopHphrUhB06OFIcmbmwvkrBF6H
3Lv8K6UjCncYwFdoygz4z/MvScGj2UkCdNXb+3mrgWFGL6fcJ2ptSXxIfr5QrtfTt1IoN4AoVJO9
OsAWC0QH76MSgcbcKxdVqdSdwnmQzhlY9TCm3BReF28OVG5ODawX1QApOIJlsuw8BySasXJ2jDXY
QhIm1qlbq+7oL23PAOwQ5UTH7IJszYg+X1fI63tSncn0We9IcBLh2b0VtNf1n4vqz0dXW4qJwsCe
FMb5ZVaj9nGpeW/OGtbeAZr1o7pdvXZ34HL+mxVsXLTHpWrOxRQP3aZjjqewYysCQ9ChjpKkhlMA
pB/r13/iPj5qOOK/KxJi0PTmSU/BJqap8IeaKMmE36s+IBOJ1kF1u0EFvieLYDEERil0pYXOg1fx
/67vy6JSjLuBa2xM+R3fPqqbw+ZnbYcSaxCryIvklck4zRRc3nLl+fdo8vsy6GAIZfkz8Biwn1gX
+12SXo+B/zDcrlX+Svqfw6uTZF5LzfkxWALDgVow9S00BP83Usc8bg+qhO+nyYi69lqYBceTIwM7
cGQGhhClDOZTROBnfmLrI3dHmoOJQmGhy7mQih9vCVZbL3yMsyVFNU0+lfWV+goK4ECEawl1vdiz
S3a3WN0VRRDOYJsm58sdwRWjtIiiSF+hEo8rGvExAQ2Qqmy970iqNSPkxpBq5ZvHXA5PfUP6yAgv
H1mrrvDVTVbVdXzAjxrG2tKF/JiUOO3o5LwWwiqI6PaPOH9+9umDRBDQHm7lGyJYLvHZLjaT05LL
t9S+ynGFZ9K49w04WLCR0VrIF/5Jt41e4lgQ3nqnmzKyD7GAjFtvEFRD/Ifwb5GPnnThibmLxrcW
CUAUGijKtzuTp7CLP3B6UC565EEUUQ9hnREBtlroOwmjrcFMv9iIDGZHKeRfjbej9stffwQ1AfCh
Rap7OkhrOmqJbRxdwbg/n8NNrwh+zIy26LVJIhNL9NVAUcD3x7Ua0RL2QIl3/4a5sVuTrWNEFkoK
4U4BnOGgdTXG4kpnJQMrzQjUixwt+VzoisWYqCHhsyUt28Hpp4n+r1T+EUdLbn+UDfIkm2g78uw3
p78ZrdPc3WF/++19UwFEyB9QmajmM2E+YV8tJDk/hxXdegq2pgxG7uHMr4IH151df+twVReMxVxk
czb4RQdaxKs8v0KKeuQfRiIEd/1hVPyarzCwAPKR6gV1FdNaJVfvnqFsnzZAOVxAqIWACz/aA37O
dBcjCHm/lKBdMkNioOVvFfLf/QlaCyVKM1PWIqIC8tEEKX/twGLqjEqypRCrd4ZHB3UJzKgQhzGi
g/iMcaEx2XuV78CYOxgPcx0eVOk/Xj2GaOzCEHeUcllC5LRBwGq50M1fCzzswj01+d3OD8GH/y+R
kjs2zdqdCFGvgAnQI/pm3jqfARRJUj+Coolj8qpoQPJ0p7cH59l5hZYfcJN73jE9h0rgxdfHjKA/
HTX5r9zxN7ULRVNhp7Gyn6CQnZj3pY300Fu34yVmJFZHPeE83bY6Br65Xv5idFy6E4sxh989Nwn3
0vexgNtjt9bH6+sUtIhGo6jQ4LyQItXMumYNDE74aO5GJnJpgCrFRf1gVyYrzL+K82D458k8cEI2
CCUJNV9pDDyUCc1oiKBRB++qsBRO4ALErtvhYF8A1z32ypA/YLJ+PW0zFD03wwhVurrjh9AQ9P7n
foi+RRpI3LIjEBXZya1kNxLZN3e583KbMsCsVWOAiW6PjV3fz31ZapMHr9s1VVbZhSnItgrCb/kl
b0KKetGgJxpzTJBkABTJTAIjZg2GdPGCp5IdZ1kVkd0YmHLxp6K7XlHdODuv6jG9RM48ByENh2rX
IOGb+xQV9uXg5+ZRG9FyoaJDcidAn87Hq43Ad2fx6QhK9jFLsLrCAuNzmxIDfCL9S3RLW6qHt26k
ZvguXDyfDYtwOYglspHVWL5GshwSlQmXLuUblVhdaOwuqdT1H5Tqp44oI7Mb0/YlRH8RTNfJ6wSx
buLflVfCqBCJvylxD5hJz1VecPabJlKgWC12xo+jtNMMCSIHkvFnZXIbQWSNoVIcfiRgj2HR8FhP
7HkPnUiTIwslsQYT6cqlsuPI1kuxDeNC2eJU5ZRy6vfwtRvqcjFkCJYIvkBTeTfG65tlfqpg2qp0
TfdiIa7kH8XZXcY26GHWFp+Jl1AQbQwGdrWtXO7aEv33kJgkKQoH2zMxKnzyZzW8Wfdzmnx+2pcw
vZLlFHyan1quC8V9HTKX/4v0ki07OlTHn71lAqg5w93FbWXN0TYgXQkJtvMze/pCs6jAwWrr6iDN
JPGFe3yZpo/gr/Nd3NGNfXeC3S4SNSmz4+WjKSv+aeliRvnaT0xv8jlsAHJ7d95mA7uVSOrrygSj
edHg/qGpDwwxp9WsXgdhkc8P1jm78wQiAQE6psO6CjQzi9MZ76PoAIW0CTy7UbZPvDbhHDNp83MF
c4wmUVYOJCUYBl60FPHG5Tc3qIY5HSba5FcR5PHX1NMpMTwsM76CyBKWYNlVOuTRffi7/aMt43mF
7OQ89mVjdJO+4PILjENwY9v2iDaUljDfRKQF82Vr48Hio/DbJbeENFIvzSRoUudy/BH1te1uTASY
xhmqNlDg8vhTuJXKw6M483bEC9PYwLQe+gu+Gr+E/I0SGPJ500Btc3IveIK03nDPbuMShNREvCFq
GbJQ4BeIsBTzb8Vp1HYavmfibJXkvypzAoSH0qfpxUd2ERnoLLYBzOkaJcuO+8GKlIrjaPyiPrBH
8AQHuS/tMzifjoNL3NhcXJx707k2Orqc8lNMnjem4bRlDbzF6oRJ4IHPdcjKmv/Burf38JPS6QAl
zELGLvLl0ctN++oytcFWO+6R/0CJ6pv47l+xGuZa8dNj+2Fdzt5Gm5PKryYESka/tYq/27PnAHaQ
Rnd5syKVwYE0/Z+kYJCZ4whuQTczADx2o3cIuEiuEhZaVSPpMpv8pIX7spHMct3JUZ7RVxzWc3xL
k2a/31Ek7h9eXQ4Ms/1oZ+FiKl+WZt57tGCAYypLKiiK5dT5v9e3OEfrIZfyjXrCW3JNls6rpzQM
0Z2eXHo6d8VGXo2Qyc9QnQYaDQ4VGrCMB2grcWHm3j0+KfLF2c4J8wZ7L2M6K7utMVEajOOJB8R9
Jz3bQZsA09r7Zq599g0ncNeY9sHP+3OJGL/JoxmzxkZwI9DyAWfn9gL9OCZrppjGfGykBTXkdeL6
0/JdReGdYrdBJ28iLQTKLKPdemQlhA4tTepTyFR7Rt93GbFpW2V9oPUuUNBa8TOJRiep0/sll1vk
FtwO6BecH9tp5w19aKhzadxwNqKPxNyl7zxesOxKAqSfYD2tjbSdjLv+vna7IFfOgpbiyWEq14ek
6RifACE4Gmk2sCXNOXqmkt4/TqGD0Ndy8ZL1Su5Aq2qqOwuH4Q71d52Ytv/ONgb7TtAi3UBiwiFF
H3K/vSo22gKzJiq7GYA5S2tRRJI4xvtKqttNbK+Z67owdwRcLNr2UolT85qfRSk4clNQea/+G4ll
da/bJ9CK4j2NJnPDqNyqY7bfdFfXF3eSsHzCU0gref7xCIpbGmmq2VC8sVc8IUfIkqAKJAMahTS6
Vk/9//rQIaUFH/ia3KPWLO6SC4h7SxKNJModmFpYykahN4TYcLrvR+X5WejXSiBcslVH5s5E6W6Q
F5TwGucGE+GDaUvJ0CiZGrfKMWaCH2Xt4mrDhN/RnZrAVXc7kJD+RsZod/6nl5xmolOCLl0N5VL4
ZRQCfWSrcWuiY8l9YFWJxJbogD40cBGfJKWOio1oBrRwdAF8KK7bkQGD1ldlQJdlvykMPcxwK3h0
rNA+qrmJgSnNNl3EAOygzWoxXF2lqnt+Mv5Q3zixpAfIxgLHnOHm8DvUg3nFzVXuh3ZB5443h3sy
huNKf2zg+RcNxT0YDKKma6qBO43CsgIofaA5tv+UPGoS4+tSkHdLHOMPTrqNlTuCmgbMAzZyTltQ
JcUvzQ4rHt+eBL5JTpM9U9ojRxhZOgI+A1u76jEXNb6stPf40o+dXxYM1LxEqN4rz3cnYhZs4B2k
A7qa+Jg/WXPdO8XEkasZQoRaohCnR4MzIx0G8LH948pFVEdBzvCoQbpeleJ/FZ+7HEIZzx40TnOF
2WnA0QHFLK4WOpRh2mkAJ2WtTNiEEZSq1tiED/s7XiJ7lZGAMXqAD48uDOVkqXA83lD5klCzqA0k
8v/sD+wB5/tAWCRCHc4Tg3RI1aZ+d832aMwMdbpz2rKEBLE14Uz75TTr8Du3K2wMn7IX4dnDiQE/
JsREjxQr85JtUVpfqof1kTXmHYzWJ3WwkSlnX9Et5ZqvhvVCu7FkUSfqksnu4QOay4/H021ydmto
6JOUVg1NmfoVFRu3HUhexQ4c2oj2zWrW+gyjIsYE4J8nmsJsrgylshqDNo2PGaGA+HlYbk5P+nnR
W6Vvrnj/TsQ2JcirDXg46jfbnOhv2N2hFwIzJQry3k0OcfOMOJ2NF82n27JKNN43VRWItWX4zL3q
nhy7guiVyaDYI6yOE8i/k7N1eguZ2KAhxM+cjnetAhxH0ZnF8SOpgPsGCUEQ6ArCcquI56X/pQmB
YN0Wi3cyirmJrV/StawtTuCz0SPLdU7cYsnx/vcHqiVZl5lJHbzq1E4Bf6wo1V5+lq3Xwu+eCQTP
r+agWLYb1y8yX8frMdBX23Tu1BCRrlXYb9nGgc1oAudqTHCOzxVMg9mrKElLDMj1QPRLcHkiUq1I
HGW2eEl1CCJuPWCmd1YnqbeKB2DqOZThiyZl3jIljEqC5n1kZ2obGUgVU0c4ot998xxufPsHybGl
PJavXxoEX/foogEllF4GgD22QJNVeZuQXFXkxJ/tm82D9lHlNy/7wqJtIDK8BDMVKNngy86h/QLj
Qmn9i19VH48+6/tAukbhjpqmCSRHRHk9c3UBPjS7Nbg+UNGAFePdgv/PjAXION1LOmQogyUw//Zs
iUiwJ/4qoUc6JZEtU5NPuhJluvV//D8FzdwEM1wR2Jket/WlIgg/27fESitFU1xhTzctPo3JpPAW
vM5dGKdcc0tz9DFXD0bemZFaQa+zg2T5DjbmlNM9LTqqhS4U74J4nnTSeKPIWSjs8LlQEuXIE9md
tHBXXN7+txIDPl7ctNKoICVKrRqzJt/Nyjl77wSx/bvQZsPOtPqsh7w/xw5VR6k9FJK/ecDrICFd
fumomBil5vOv7CnlUtWD9stuAUNAGuXOCEijxFQqRiWFDWu8DJHFCtuzd7QbTwMgM0zGiFMr7TNW
KDeXigMys60tUNMOe4gmE8drYb0R712Tyysh8gzkmpVJYEQx3OnAXODKtsmHbMVJF6FX2xECBItw
98r9gExCdaj5m30KoqeuBI9zqGLukZl7nJLpxVWSWozmRK/FbUHlXghtD+iJC18Pm2x+NwkpsOp/
4PR6dYbT1t2rWXNhFBWgQG16R9wq2SI0bkje2OHGndiBQL5HS0hwUq4afOcev7oTqtYmYq/izcbf
RqaNeLRQUvGABFmY5wNlS19JMIwdwwaYe7txRrWJBQjWI6h9xbuCDMOkj43Gb5LtPbT/ZK2Cn+SU
b7Jf0R7vqhUfxLOC+M8NnicFIWL2Y8uxuQJKJl50c9LcK9OG/0x6p8rZhnaROLRU2BW7W3Wnz09n
+Sle37/DkGQLGI7dpKOd3gmeZ1q7EH+NzMmTDTTlV9/+Jtknmp3lgsC7F4KuhzgrlVjO0Po+i4Kg
swGr717ibG8beslcM9PwOMv1LJN+YZSQ5wPiegzrAcI5A1sBanKhT/VFoSsnnHwmvvHQh8Inf32n
KPtCkjcG8A6z+d3reyJLPvSYWy7Qkg/rnq585qypM4ZDx+U8+qgThjn+Qpg2oGpZrud1EuM0DYng
Gr5zWKTz6M8R45AOzy+bHQvpPaq57Fzzh4N/P0FPuvUCBssEQLxUoU323yeUMbc2dlgmmLGwvJre
ZDjTZqpWC/DH5CdMcCunVHGdE20Kla1cWS7E05SGKFeU6SqoSoOYlf1wylSEaSvF7Z29pLOaA26n
rGH6/e2jyDQovHsAaps8xPLps0I2LhgAaRxaOsfpT/qCYwY1NEIWMSH6uCVUPaOZ3jC+f0+8d2j7
E+zgKJQETKU42ahTqrz9MvDKrGRI3g+p5iRBz1BOGVeBdQcFc/GheLgnF5TpzvhTwOHBGI5gU2cC
5rl2aUTGOTxW7QRUEH0jguzvCQV33WVKYWVDGFeU60TKWuqDqOYL2/rKV88DExDnjiT3mNwJVUmm
Q2lTes0Y9otLhN2fqjxtQ3BFBhrI91u6H47c8jH2zUCrnNCXPE+RLmaJR5CCIYtOY2HUEI8XEUlp
rF2aMGT0I2W8XMeEF+pGXC8JLmngERRxotmebPnLX563k7Oj1ZFWJF6Gty93zh+EKGsYbKC698UH
VJQqNS/knsRfI8nvdlYHhcTXzq6pqfQhKQcW94UzZsDSN/KBWVw/JKFTdfhAE/HC4HeeL/YZYDy+
D46brqVfCwTnRrgBV0diXDWn3L52Rzs04X/ss5x31a05vuOQOkvATnWpSt+P8/Se/DKVY3B/kwgZ
IfxP5lFNnhDNMcYp5TzHkvDGsM39lWWA5G0yUNf15/8Xct9lqBRYdZ+6hNnWSD+diRETCFIelA93
vm42lATNgZZPj2oIDGsrXaIwIRpwD93MRpUQuV+/HRf1wd1/9gt7v7UnqA7SJd1/d/YArtbeFjNO
eXj8UxVV93TaMdop8NSXwvklhSRFHFOuMhXpcPh5dannSfBR48f0Vy0xnemMXboqFrQbk7ERWmAH
Gu8Rx69mD6878Y1ck69GgC9q4C+mpnl6apUD6aCu1s6hNmYvwowgWHqDK9bBj2WG3We27zSijNRo
ezsA/x9oeIRe9htmhcEC8hECZM5KmNxwYUbNbp9QC26OFoj7VBMx5tq9zd4e3YzBA5FwyenCM1y/
SzfEVxYYFZsuDFQLvzZ6Iy9KFDwJj3+PZKjsw7B++7j/e1mKdMALV8P9WeVrXc20kgRw/ZUen6gh
VJ9tLyB9ayQZa8WNf7sKBKZKoMtzNppLYztv5vs2O5D+6Gh7L1EfqAWGsi6Pp0eRG7xPor3UvydC
jhWa687RFwYvWQyQOLEM0yl8sAVXV7TN6NhnE92bQMYDt6U7SWSHDU5t/uu85L1p5EWNHPw7eG3Q
/dYbDRPajXwvyb2RP/BptmXMJSSC3ar7Nmmvkq4Jrx6rGvkTHnt0aGEoo5iM/ypPDmW/JkT8UPeL
S8+rfo2hKTWGFOMkv47GFOlXYAbXdmAh5MfBS+S6iHhmXtZJNsoxo0aNnP6Vzi9jnzFcIwLaGkwZ
n63o8LYqzK3uecTIvE+4YBwzag7C8EHN38bD4kdns/4dYHMvU9/8iMQdxJp2g9V9H4c1CGvSOoyr
0L7HZxDvfGxsM4m0myTfyYacpKHqUtcCZ76OcN6+RRO/P/DkJBePUGeyNNqK2qMxas6L/D9OIe3e
qEiTIHE7mNtpopoCVcjAyyHkBuKfWkmmZ0GSrvRUwGFBmLRNjiEiZTDKGiQdbyVrRK0/fYH0YpfL
a3w86ZTXIj0FnwO6HL0/l6kBF1rmOVUhN7t79yf9EkrCh9ov4ZS3nFKlwPQBog3wWmyRmHkV55kO
PU9YIkA3iPG+ER866X3T9ZQ+LXWy5u5vZIsacQ9G/M1FaymCzaQGwwUt0LI83xWCebRTyTxnG+Ym
oc4TIOLyeOU9duPEuNny4XLwrkaa6QGjHw6jDgNqCRWeXDy53Y9eaxVOVV0cuQjB/uU7occoY0Pe
Ta2elljnbjuTDOeA8qbRf3y8BCAeJn6+IQw1Fs1ZPwO/QeYSs5z0HzQJXGLZMsmsFTVIYoqI21P2
eLXPW9veQVoZQQmH92eDS27yHVdABjGOsbuEynZM6dDSId/3Bt1BX0IPAm9CrzBElbUgDWRf2gGQ
JP6LtFfHf7iVQQByPtQHwyJUhc7Kh1ZQBcvtRXiwnSUYo+xMJKMqy+zVV6pq+0i3qvMqekWZ7dWL
wZeBgv0DQvQ5DcIY2IQP7z7WjYb+4mKliO6uulJyiNuXyhdQDet72lI0YcUliaILY+oRV7x+eymE
8IDq2ICqa1KVS3hVLHjtMueBFnxecRkeMaJ+xuCw8ruPLkxtg7G07owLL6KKf41Xe48665B1qal+
EBD+bLo9NZwPyeGP9BEfkGwF4LyWWE64ah3OWoUZAWZXafCrFzsiQWZgHx4Xxu2Yryh4I0CEnIbY
twIgUOIlZX4XzRneeN8Dmv+6MHDo7FQ2+o+dGGiOUX02+9cTyAu1kXq6vyAdh8dAadmjzdQsUF41
tUIL4qmeYp3YolgCsEFpV0Armpoujkj1XPEikkHPKAkrhlzrq4Bn/LMx5aaEHr9jNVQQ/j5rSLzi
/EBJ8k7Qt34OcDj90Rz5d0idDXhtQ/pcTK5rlddfUjEqNRXhTjz3CF6wm367AsDmRlvkEUw0CX2r
o+CV58Y88dcYZqopRW7DIUiBPPx6KyM4OWVxFHMe7Spi/KahQViC+2yB/oeu7zPt4Wk4PUgTiP8J
wS13KsKVu4lZyaX+q9CktS7k2YO/tF+C4XABV995AW6+M+YjF1e0WcLP4KZbo1ADHxfIG/ulJwQJ
+e3YhiUZ4tbyzJch3qCdO4HkoXRTp5EoNgEaqJcx6Q2i5C10NEh+04mWjLz/kd2xcTHZPCRQDG7T
E9S0ESeah7n82yl1paNpaqCiAkoedmtw8GMtqTlGllqhyNYaB43cMFQzopBddM0pnnrvIrFSY28n
PKulNgFUjFe8oracLeCwSMFd6Lf86bT1xfxOs8GxRAVSmAb/t+YCcQmy868MyvMwaIwXKqhEK5/m
RK1GxmntAtKw/3AfKyswQC6HVNKgmyCuA3r7wJ/PPC5SfBJ4Tuuy8KkA05/hx/aWRCaqgoDyFAdY
So9t5XV4nQTRWKW5GW7VHi1PkM7D13xvIIA1r4XkTxlhf0SqjZJcUoEm4aWwTzu2wXuJeCIwV7Cb
CcZ2JwYU1C0YQm0t+YQ7kGAp18cFRMKAZQ21ZKv0RjeW+xqa6C5leIEsI1afgdeg/RPiHqAbeVyY
eO7yp30L7vjiujDRnYrAVdLBAgIK1Ap4CmCfTlUXRDMVf6AeBRV9Ck/xc1Wl073FYHKYCMDVtASj
Fa9vsVi1jJqKeiKVgNn5se97wpzPIFwtr5REmNLHn7X03VXjmD/oOlLBL2kEvkiucGThCsOm4epm
l4vu3ypNKUJyrC4WAxcGwb8Shp5KN9uJi928+f6wos9Rtc9qLCdNIU6opEkLstmefGyHy1xcILkx
lAZ7oPhls2Ftb3SxFlNTCYH68c+XHGTc4ywhWqPGmSfIQEZiNGKsdkdgojd5JrtDfGpYRhoeQmTD
h0gxlrmXVzfCzcDnJLMgOboDxsVIFWxAIBxXBWEOkvDw/WXdYniuH0TSMgFqku7zHJ9ICGl/Fzbz
pj0zk/T5RKpwqiREkJeXnutyEeL2YMCp9YkDlULfmlcpFjrppUMNr/tX39vIYh8KsPC8Up55049p
T1nO4iFzKemMg7MyVu8L3sMbVdXxL2kdgSRvDQl96w1MCI1nUeZrbBzosXrt2Brp8Ccvy8twv6WQ
hfCgYnyaam16q2Kami0MEa1pJ8QiGGdxedk9vr/GaGaGCT99LxF4LyUkHZzErOILjRsKaSieRnq+
xZaJuCfi6ID7jDozai55vIi11X7YXGmS96pAFfkWZpr3gUTVAm/FHXDUPTdBrc1Tupxt8j2G5Y98
YyO2cHjxOSzk6/i26L6Oq2pG4l2WH4/8j/CRvY+BBMpZ6rN/IjF+uoXLFhTctvzD7Te5zh0tuCtu
a4yodLajSXNB0r/VHvJcyMDBfcVpFm5guN8lmZuIGpn5/TOUQt1L/kyA9AEDj7AJnOXSO1lu4tyr
Lhq0ClsPGZGsco1Wijb9MD3p4tQSIxbp6dKX+9jIqYYVHZ8AXtBkdoeO39IhN7ywd1M+CgFyHuH5
NwiyT9AoEKcfVADelpHM5yjabojzbO+UO9dgk00C9shyg0wV2QvvjTk1Act1uHlsi/kb5j4xpfe+
Hj4N5yOV2wQUOq3jEVr3SD16ILWDUgJZbjvNfNJS+e0FxGLB4XPZza+bYuBfB6y/T2LfQ9vua8uH
lRVzoXRyyVyxbN+Vhj4c0y7+oNoq4PxeT6IbndvmWyVjQYPNDaxkAQ3Aq6YQVnvd9CAiX8RT8Qu0
Kb/j+r8BgnOigEj27nkj8Ua9gIVozNUaNZofAVr2dlqky9j1KzNmhNAStgA6/BOwpZQwAEkzRwnF
ZsIei9x3L/ZhELgzJrDgypIW1osLL8ABXIh0PO6xLOOinILE8VdN/adwDT5N3oUhRPWSMJCj7ErJ
/nHj3Tdv+vpCoDZG6Mp3bYbuHoWtudB5jR+7IqKHwPVonyGWLpZuGEWErznebnUk9IMi8LxuDyLc
jNqxSQXUvPNI173xdRVNP1dMPNkCtWV88oZdat+gzH4GPCe/kxkIZuWxD0utmcBqTWU616YKIspn
6SuUPWh7Ge6Wg16MkI9Fs4bKaV99W0chLFBzqs6YSmJh98i2M1Q2PSn/U1Jci1Ex4fN8+RxQ3rSq
rgz1FQqIAFB4P+y9TeenKFHTzl1IuIHXL/DQJhk0WoPsYfNtLwA146FCAHsk9LZM5yUca/UiPJvF
0Tk11YbhlvGZ7z5eEESBao+k3DYSsKbPSNcVusHBhi3rbXjxWITv0OJyBrl4hFX/xemPenH10iCg
c3SflKABsR+A0f3A9E/B3FLQPlPtc2Db5xO3ZcPtf6KeH77J6JtkCUHIKmU0ljh2wfEg+Jh+YbYP
A52SD0gfbJPlOoeN5CjmXxTXQf2PZt5kKUqZSI/eqJsBg5u/w2+hhJ1GAsAWlaFBz6k/kJYPMV3T
vh1mHH4zCMe9Q4OiuYaXKQaiX0WqzWEEwjysmGrQYVcWEnM04Y4rH2DJhroFkVanqBMuwGKX8Fn/
1A7B2xsY9izPTGSvVhFsMnXRAJH2p484eUN9geaPahHUNG4oPa6WbGl+GYUMzJ3/G5Wunm5gDqpt
i3xxRvhf6ncAag+tqNQidZwN5SsXrR7mrnuzFhzXYjig3I7gqvk1/w3HSTtlmNpbbfHzTW1zJTV+
LzOpZg136jalB1Lt0/rQKvaLpaHOSS3jhNBvaAQnoBAgqwcL9k2TBsBuAEMJMz9grBdMzCVioeF1
6fuDfzYatqr0nyH5iDzcZtJlaqxMKwE6XRNwSTElQVqxN7rNXf5GYfFEPXqnRvVFe8aV4qIqzyrE
LInvzyCcSk5cnyTP4cTZ3u0OFKFRh9GqQxQYaUOr+XA6E7fnbFgza3YJFK6xYSKYrH7LtRKdz1bQ
cWCwwCBi1mx+dTpA/IU+RMFnFbo5/oCYm2I5CiPWKRRedaHkNhYYuAdfrWaamsiUcKFyX3mgOXRo
wKJNt533t6pPTWAKOIduPjfX/EsKAmvkZtV2ij5o6ts4IOguosWYNcHy6cM8gZYekLezfLmReuzE
njhMKq3/++vqhfACYOV3QjrFBCfjVr3EA1eOUD73iA/ZTBxUn7KlR8kgeVWdWcuDyj1vAk6TAH7W
Lr8DEBWblkBW1j68xN7DXSTl1aLgiiV1OhD4I0/0OpDcOcj2DYnQtVN8j4eihLQC7BxpoI2Cgitt
h8qjBy5FHkdJT73lBxUjA76Yb6QaOhgOR6Fkr4sNmkun/8nN8cvY4/cIgGMLBUTyq4W7GrzxDmJk
0CVe6HOikz10+zZ97FIhRXSl/Oztq+En0xpY4esn6NrkkRE57DQOIw0G2AB19lChhMO5U85blEiq
ywKLLO4Ll8aYP2ugM07UmKgohJrAu0ZZjTBZkgJbKLcvgettFwzlIw16S+od+Dd/UFTv8JNwDrCe
BkRYdRiSVsPm//Hk1duecozMIDOv9e9ekase4WzCodxVha3wjmdN0YLaPxTW94COXbnuQ+xwo/fi
3S2MQ1Bkgw1rUNo3AWOQFlZYZOfuoCVj+zijDcLaLwWDlr0WxtJAJpoIC5oCjh0XKGsY0hhOp4Tf
pmaO/wRNGM2frQXj02mR7G9+xzamzXNExVnDsz76MPw5M2DZkLngAkAjg36Fbfyd6RlZdpExZ6/R
wCoLlmhegu/Gslyx36Tl6bJUZn84/uTND3SCFVBH5ctGlEOxv/JYRyN861dzujJKvV6Izut46t0S
3byzcIWaHT8H4JCcIIIrueMadX+PCPetq7/epv/kHvN2VDUreandUYDM7ETokTglIf7by8qtBgbN
RY+JO83KWLegjgIwut461P8UYL/KWu4PUyNWfafGIPJx2C6e49gRBoOSr0xXSQyPsvNeTNLN1GNk
dg2GESe6Bjtn+wNnCs4fboIlaxvk2tb8DjABlCR6hLOuidcAUR4FJVh3ogXhridJANPfMvSC5/bI
40YEiCfUxlWwtsWO/1injamNp/pJxJOazo24UQqddOR5samgTVQK1fEA3rE5b55xgG/Bep3IQ2fe
o3EHRaIg1l4IC6GqxBdFASVTEykP2Hn3mutF3303ah2NVsFnlgID9H2kO7VAuFzg4NQ8XyVO/0YI
smEBKZfQrWyUESjd87amu35VWKzOuW2H4OiFuFBo2CmhTj5hUEaA1ONAfhgIUnRDvA1FtO5eKA/C
s6+dXJwo8Bq5tPCMzzUjienqb2n5CEHPxNspO2kX2onmTFRPMVesjJqzDM5XNorjeSF7rLhAwP5T
D5tXSZJM5z5tCN9OrI4jA+lhHYTZDWMOcOH0465OJyE6IWx4Y6ocfRIcAtsqvhioQcqeRH1Z3RbU
Umh/7npL7OGfd/97XtjxHmt/+eWBTqzPmKgcKhzFR3iVxZKvUM7k7q+zA4N7s2hLo0s8DkVF2xk/
1RwBpWYqjv3Nj3vMX193DsSF/yKRYJQelGShUDGlOlSTat1q4YQAyvCflw9JVT84LRukwZbLWoo0
sgmHNFL48JHh+TiQucI7RTzSvxhabv6fsx4ox4CfmEtzGTQWECF5iCTLqjTVcssFfGLpFANeRvSV
VPnHXt5LD2KvFd3Qqi6umtIOMk+e2tKl52x9MhYkmwIjW/jEHm5l4wZ1nNXpaRVlOFNgCDqc3qXD
n/SKzJnM1aS/KtTrLJsM1M95wASgVPFfvVUXfsEa6QWBqchaV1R7bDTz3EnLV2jMT2IZfXSu5VwQ
+zVA4kpE03V2c0eZxL5dHoxQPOgs+MEFeiA6YhUpIZrpEn4CSdu3DJPNnA5cmiCeBShdf2DhgSkc
WSfDdl3kcO8WkNaz2g7UTSS/AQmtlPWEqFVNXkUTKsYPJHQ1fq7VGuhkEGwnTPMq4KfwHvjzxT/d
8RYb7hWbvFDr94uw3gNNBM+YGNlQ/IjLrIQ2Y+VMqOgNqSXUTmZLfzf2k2+FDvUWIfKv8/9Y1UKX
h1/+/6QR3MlHTY9Kp4KT0nXZ/vq3F0QOjwl3/0bzSREOku1FXNJBeRjOZwkTiTgwgCs1odMzgOel
18oN67URvAtM8NFrM180vCtJr29XYyzeXB1iVGKEExvcy1SSDYh3CBQ6tiA0TDSyu1Zxebv2NjJt
hxCdCFGQrDyqKBHTjEXUCpjPvyHKkmXOB5YsoIxhVtgOt6ZkNZa3kPxs3jzZwRwf0Vq60n0gyQh/
c36G+QlDVWNBiYcaAbfEIYcImskIng+AfO9bnlX7xD+c57nJyfxd3jhnLAqMBmtt11BbQ4fzzSrC
wnaW48OM9mv1DA1bOxKgNk+WKM9jH6N21Se1YNzQpegHflFp9KKylgeZxpxbLa/n+/XSl47aQugk
xY2Yei/W7k21o9VOUpNJjpBePb2jGlWHFEwRAGsoQU+Af52WD6ex4x46jOveA53vZM6Nax3xuvNR
2a3snsOmLvX4w8zX36O6fFmLkq6dwIAbc3jiyqhDhEAWrABp4WyGcTYpvqJGlwKKklc/BV2M/Tnz
aB4+sy6rgJW7kD0vVePFjQQccb2aSCyvFX1cQZnVsqSTV54kVMgaIQj7rpQABPDcPuea86LlDUtb
dPPEJUi1i8x+7yMYa1FP2kOmGgXgKYfvSUoSXCT7OPX0jfGhHLomtLLeqKjGK069Zngo+ww4Wykj
YEi7s5233r0BWqzXeKMwkRcwhPxKEOVvxOboTha071xHDsUM8BaC6I5k4mxrMHc2SCvlzShRGqKM
WUukwH21oY+wuhd/mpuqOcG0+Fqc2w4KsvdS+sPOB83lIO60J+cpVizJqArTLb+P7V1LapTkz334
uK9/BO1qY8KtXEKKau0ZKWtqGxDDwB5XLFFbRXh+zZP6d9IWIQ8zaQj3Bxw+EEWOoD/+Wdq+JJ4G
vMFzfBhUXRR/ahe9poRRMxGY8ospgP4+78tZeu36rVY5ZD2uGt15TzMmcLajBALK5vktthJpCIWg
NkoEx7qP4lvZngvro6HDA50J6ZaDRPU2A2ZUyNUf7SZo+oWCJKVVE49OaCmZglW1EWR9QyoN0pOf
bTZLuBUDtF3zhfscjJ8wc9isjiohk1F4uq//bZ53LaZfTudlLAZ+NL/1kW2wOfBBHeMd9LzMftBY
F+bxt6B4xrhsfwT5bZNTqzOrwUtNOq0UMS3ZSRc92KJ+jBZpP0yoIBLzpyw4TlmF8A7ODmORCLcO
uK0FpjH3UnrY9iUwbk1goKcYF3aRs2Ov7gIpV7ci6Axc0GOu+n4R6W97BS8g0Mqmm4EBSIfnfgad
f5bPZuRMr/gHUTxgWP+GO9MZVKrN6US9Uaho6pR+hdOV9jwsn7umx1HaIVx2hFsZCWTRlq3OL3J8
B84anWT9B9jJ1OVRPM/7IZSD4Kq5QjT4DcXjASb6QZZmmM/RSNzZ2DnFDoY/62pLP+PJjW0XeC+/
JNw2UAPAiseFS8hERwU1em9ppTQdnHgc6Wxzfm4rzDhZyA7QCq/j8DJFnJLebzmm0T1yZtQClpoB
saANr+O41XVK3SxUcOpBIj86TV/Uzw5cJPQxUbDmmdnaSI7Id1W20KP9wriM8dSdva3B9fcZFXvM
FgwMHf62tIIqxMJHEBMWSJbcPEFSxpIKlszngwce4FigzUN7SGpvkhWollyRo49EOF5siRuy9RXI
BMWVoeUTKYtNZjRQVB7w61E482w80YGwo4CB80o9GyRWmejBEyn3K9u4Agm7dloBl14cWhl8NPr4
CfIfNI+dZfKMOo8NpTfOiNhYKi8IzEo0RMdave+hhMyWAfcbHDoaLJGs8edUb+iEimvam15uaL3m
zJo3rfaEoO90UfC1tkC2K+WKrZpTSY7/7PLNZ5zkQtyQYxqUMAM0+1L92JpqZRbWHnM3078XpEl2
UgL32ZtDOHeki8Xso8juubloQksWNKkb1M93oqWJltydJfPQQuptJr8nl2M8SyidqoZAh2vnjNDu
w18a/avm5w/1ytwpF4q1uRPQUWCcewZ7h/w5XkTuBqzqLDfmagWwl9j9qdwslJRDgEkddSZaxrv8
HpRp1V5oxEQhcrs/VtPzZumTfZtyk8JzkE6gY+xol4YFCl9R89wM+JvaUm3kNBcQQifnb8+Lsua/
nBZNli/PdEMGg7pS9X4sW33h+LmyDenrV2tgUia0ZK27UnG/TRRXzMYYZ4q4JTNQs0xEktZtHns1
jwbRU4GI5eBLST+vZHZtPaps1qLovIMNJTBUzh0CyodztPnWrE32R/Fz0HMW8t79DUuSxBYOTe/l
KYNX/txEmieHqdMN0JnL7hmqDvyDyOtmG5KiILRoY310/F4Rf/7ZH4QPWitU1WoOOfBU6S8BicX2
czODCMF/NbQrMH8DNUE3VNqA5kCJwY0WkFauZJH1XgRVgttddq1hzIpN5OGD3t7pbuxuQCAGhSXw
quXuUwWrOajOHBenOsv8IEWOcIZv8Pg6/p6+fw19N+ltGd8VXbtQo/LDNJ+69F1CRVsECqnsrOlG
h9y+HL47cH+uM5JruOoBc7z/svGWntRktCA2+JJ7D4wvxXs5bpXdVxVx9AOYclQUPjiY+yMM5zNM
lIvv7kkroEHjJoiF0V8SzAwisATatr1brJ3BJ01WrliCn+eiXr/O3imyiOonlp2PxsIpxVYq3h1p
xCnv5rKcg/orDrWDZ38aNk1LnlbOIwIaIXBOaiNY0qbpQsLGABaG8RWjH5DHj28ZxWQSzNk+aIfx
twkTY1dJ9y0S798UZ12RF6dbSR4iaYr5V+tvFpQA9nKf4x0O5X6+fR0+LMQ5l4tfuW3oQ+D5bort
QOwbu8oIW8Py4P8E8JAjWrwXGJfvvyep9Zj/ryzbSQtGcCk6S4LhIomY/MzVy0r3AC4fHlUUolN+
Q9BxTPP5sxmJa5A/s+n3DJRObIpYuJZqrjlR2DtBrbDZ+/OjLNNu9WEskT4XCMAhudNBBZ8PAiMu
st02OwsTdw+fJHgu7HFd3OKDHutvn1d9pJyAGZ+vmHeWQkWAdNzqs89Cmawf8mZ9QVq/ImOjykkx
H9YwjWAaaMPDDsK2+Akyus1hrKMgsTNGE6h4+4lRI91MXvf51oj0Su9QUc/l9Uk3fjZReYNQgLlK
Q1t4lfwHQrkf2IAfICPjmkTm2n8uakK1jpn0/WUzETQjdUtf6HWJ5IhEISbwOHjEk0f5MNDzWJ+O
1LsZOGxln8zZOHKM30Tm7TfCr1GVszMbkyNp+weVKAJlt+NMXOalFlEnAdUPFIG5pTowBAloIGBO
L97NGZAekOP/FCXHOm4ahjMDLzzNLCehXhJejsO0dxBhGkt79vuoaq2kzadcWinvhTFwoliFUu17
xhsiEfIyB8m9Jov7bnHFN5iok5JjLRVV4Ya7Fdx88Jq3cvnf9wE3EnH8IQGkMJ8lgnNdWDPHPE7I
LBMQMonaeAddM85v1JWYKqKmxdfngc07zv5NJsn5JkX98Hu81werEjaketh7s18OtylxsxBK7+lz
Z9u8NRu/3HWtb7IjmQ197KAVmFnObc4ABldI1V/PRh24xATTn54F7mFCX5kqPVXEHLuSrhNl219J
YtZ6bAw5VtU8Ostw24ldoIMq8KPjPG34TYAoaQvU5UesUwrIZisatMxkLigPcD6s7lOibfMuCM3i
eV73lWkuUKEHSxRMEDfIfn8Ll22nqGmImDMteT40fX37dscxwZe9/0a6xoCgWASK09bMyahNOtpu
875mTtx7/Jv4x/HVjwUyRe0cldS1PNmsdDb36GiNLPIP6t/vJ8emPbklDL1zW0VFKpNldyXuaBGa
VCGVg9ycx7I2O0VtZpulKdqfp+r3y1N4YN7NLLohxbg8UG290KiRbskhtqPKRYfbRTZFp9CT3oCp
iG6gSatyJfWQbC4QwrNFeK3l1j9e526YG0NGlW6J7TbBDp9nYyXwLFG4FM6oWGbPeOKOpgc8U4wI
fo6f5QoJ7QZU+nRvkxAswGCRPHhTJAwo4zbJhibEFMqmZCQtvmMrlY262+u+szDqMhj+D7s9f1Ki
92v5/H4MajYzsdUJC3bWpZhTEQ2rLsneYIKskTtGGC3X1fsUUZoYP52H0uHvyb0dlvqi8HT9nLDY
uj+g5Lsu0gtDGpSD9hx3paOLY304gdhOp134uoioUKcXSWnwQDJBIaJXlPr1SGYsfuR67Y58eJwT
3zYvPCBo4tebaoGDad7X//QeAQao0q5Ugy6JSi62vFfWOzk4hNQ8lnH65U0jvqXvfgBu1uBHdxBp
Dp5H6bu/cCh33t0QYxKJj8OsNpztb0jybFOFsQji3/8XeHXsd1nMyVuu9n7hVwFi51a2fdvJEcoL
FzfVag+NMlZUeyQtyF5H3213xxGg6/SbyXDg7DYA7xuNquypaoQWPgWyghfxcmqSy7RdiBc8tvi+
4dm+lJ2vgZmPfwUy2YlISn5/kN2ctqCaheFBlLfEGUb66bKctaiTsokpmR2To9BB0EIOYhsWg7AW
gzLWl1xrY8j4Kqz361+LE7xY452Rn1uKvLECVJlRfG0/O2zwK+vb71CSFCtXo/qIA6f+A3v+K/vE
OxWER9V4fPrj/uakXAr3JApy901jfE1WC/x5jsN+mKkMhWcE0OOPQW/hUsHBOqt+VMWaQPE3CkEu
eWaKrpQ10aBXdUTCupHSv+NavBWzQ8A8UW9o/ToikpiuwMrkopN9Y2Z0EnN54WGEL3LqGQXJZ6OA
ulIAresB/Va2+oShv3n4RmcGaxYYdp1P3/OTratMXox/Ts0OXPNp+AEK/kBWjQGLXgrvF7e7/7Z/
HmYU5JdI3kQK32FSV984HmHhCLfYN1mZI8A83FCJCHwfXJsOC2WHk/ovPt8is+U3oyrNefsDpQ0G
CKBP362rTl74T9lxk22fXzJrm/PZpPe+iDjgKWG9vrxDI8SypKXyK0GBlmWqxOjb8EcI9p/lugGJ
nOzrBGCk+sd7EPr1PcOy1AQ/qD48idzGQ+45JMckrUMK1JfymwtTUH5HZM69eg42VckzfFpe4B1W
Hcf2CercHI1e6Md2lOVjgv+0L8ATYIdxP16u6ka5TToeCcq/QL7+PZ69KqjsVJrr2YkvWAiNoUw6
TRI2xJ8GrGxXWdSv/b1kw8E5IFn2A7j4SNgBEzU26f2NfnJvK5C90TvsDl9iIvzHaunthHR8hcUd
gkXsfgaMcVTjbk9RqHfh7S43tRqZs8VjRzlNj8yyXARKflOX/araxwlNuFWMx9BwY/SGIF4Qo6b/
K4ySNonWYEqsYbBsKSk8Kvj9IoU7KQEe9q0ry4tkLrJbgoY1ojZd1AHZlQP+ocZFSJnnSUsYW2mv
6m7wAZZmgIEp6FyQSiynd3S//ap/LCtrX7eGhRDD7zHH/UPvoqntiotDor5o83nZmwdQsOE1c/hf
VmF5lq+bNLXhaniraxxqsusiAsQ6WRWmjjmkhEcIiSGLd9S5QXleqy5Iw/0KnJlxzAXJrwMn849k
WZ0nPPqRRf3bMLAm+zk5+9yZQ9ILrQ01/KSvw0SyogId77KoA+tImnvxryUcTc4Ekvq0yDGXQKG+
NnVTRzM6zcysdEiRaIc4yXOGihjxmz4HmktHJp7jLkRw4GTmxKzjDFLR7QsjmMunv1esYJhmKsXN
n02BSEjuWu6aHosDuUX1lD1xW++NnRePyeO+jSKNzERz1CjblFoAA/qmQUR4OfZ6VsfRMVGSAlFC
N3l9RIJvgbAhfroJrS2+RqEy+qlMnxwklRTdzj5iYKOaNpjpnEWo1fOcZrGbrJwVtLvTr3SG3yJM
MKMinSdcEBbWhC2GfZVEYCUaBwid7jLwyWtMlPQcCBZLC5A/FyUQBbMFo40r3Gs7LxtUhnYJ9GKy
nPRjizCDzPSPwzzD0boWzRNV4vTjIJrBmzO5xwngQaKp3funMDNCbRnGZiUYw+0CWh55e4lIwxku
Drp242+tRlQ2GbrRXBSqcvc4Uf7Bd1EyyUKfZ6j5v5Y59QWIOyEHDXqgVPuCk8TizG1zLA3tqSR4
6CqiZzFgT9pCuU4GjMHQcPt/vy1NflrnnqWoKOgpFhqu8il3M8wPtIUHbfYWSoXKtNKQ37q7FGEN
WRz7/A6+hVbxGFXnRcAY2c4+iZqlZk2WyiLjbb6sRWWmZwIvUCXFpWoJ/8azK7SJsmJNQezBIhSg
e8TIoaurrpQ3u6X+q0IkMFHP3ejTZJZtyodT6WRVjpNfuYeQKDjdX2o4/ecrujJ5n0Jfvw4TZJ9k
D7su+hw+Iha2S4BN/i4Ow1OcK23R31MYWLBB2uGGuGJDx8hhPspV6S5uJNNFZMTLXzF3UZCbPxDb
zObtyRBY/CPV49jxtX69wnIeQK0+ktZfIdNJoKGfQp9yhObsMebaOwFbMqnAyD3klL4n3+s+YS3X
Jp/Koo6s6NvpcTdehm1+s/pAa0RJdGnICafSOO95V5jym9iB+8qft01Y5vMcstPDpCfE9EqHRB9P
/PkqbkNBhc4r/pm9Sd03yuSN0G+2KC5dKSKmPJUdsFgCUJZhUDfKlul2/gJL7xt+dbl7kHaSwDBx
C1k8713q4aNUMNEgtiINb+ABkjnkOtWpYoNr4Sq5Fm7REtPfzj+XyEVmIaC+fHl5Xah1MvLgs28P
rMHAd736h1ez/e5XyOa69VMKZEzRxoh4DR+MxiLqTg0nr0uD98iwG0njyfN+kZKYHC5DpcehL79R
9LpHmBxA1iCRevC8Z/FpeYpXhy04ySp7pN7j2VoKHqUElhQWcKGsDKDm/rcpd1ht8VxEy3M3v7R6
dwHtpqF8yeeVaXhCamVaW49jfY/DYfwUjs2xQ+dRO7UAX4BuUq1rHlCuhQIzhwse035geCDNBI/R
Sh9h9xNTm6ec+2MbiMaH0hizgdYThZLsQq3t2laeiQL+kcGNZxcuQZQ9JtgCQRdS+gKlxKnHA3ly
suPDzM5qjWl/TnM4ciPFUIYWYHmXSfMeUPphjxLJ2jI0xpZij0hVL4Vm1rEYflCrs85cDDtJBKdN
egW2dbveorzudH+qJnoyDMseE9ir5nrsphMdUvTUnXCl4JjG5W3MDXwSV6V/4CO1u90ChxOI2TGP
+KmT1ID7tO+6wRg73UFQ4Z8sbTbRxgwMGBp6n2gXVltTPpZHs0Yxx8L/VpnxldDa3jjLhiesLnTs
upLbcHmScJK/DN2vOaxVq+sQoas97Osz4zTRmiqsGGQIDx03+AhVzUMA9v0QP3UL88Qelv//qNWq
jj9uVNc+fThpKJljHNNjWPVdTwL8Jl6HzO+9pYq2nRWWUtaX2Id+r5lEZNzjbF573oc1/hzRBCp9
PcRwyuU41T/6IafbGDziCMUFLVuunVxO/oHIj4/waXtSBOuk6f8/FyYbdAirj3ohrI+s2cLd8lzx
ULXTxPEGUst+1RXG5Z3NTjY3uU+qZxs6XT9munkbtnWzcSE2hMBlzagKjJdGLvUPaaZXrnXuggB1
H1J0BwDpJY/plFdsTwlyjkntfXPgRniTqZezwpKYx8uNUvNuTyitqvAPZB0F/YVYq0ykAAZx7j0N
SE0HxXVazOBscwY1TjFnYI5o9sU9FA+kZpI1oYxoIgrLhXRdLwxF+Q6TPvkff0/fdQ+Jy5nTLlz1
66GS0pflSnjzpdwIHtrmoP+V1a67Wb6N5QgBmfOjY7SL8QYEJqkw1yjZH9Mz9tA8De5otBHEZTqH
2RA3a258CiyPHFFtLUgP4ZTw+pTvqizFIjCzFh2Fnm2+9UKv7B5TdOCRyxkAyIinDcIdtefRvOMq
pqRK2uapDPObtJnQ2KeHikqbt0RyJ/xWeUINB+ImyspA4pDr4KlKlCCf6TsFWI5KO/L2KxxMt03f
zscR/nKAVdkT9quUxxHF6pPsm1+II/rtjWJCN07Ofy3mSVeb6Tbs9zo0jOs+Aog5QihodAMprPZM
reV7m6etMGQkaeSLHFrV3pgsBYmLEgJ1k42ez4O1ASTiEO/m42sOSuaSgK/VOASv0nfOdkRK4gd+
N6JXQ8/nl1dG8MkaQhJWDhYsJNDQ9lLwn8LlC0NxhTanDmhZIfLMjLErngexMhEaC4KaKts3vwJu
ckYiMmhq8yS0CunxyHvMD1130wUYO/myPqiMVrAAdkjzkiYrXmyrUuuQXvoDU4cpTa96MlJkaQbN
53rzIp7BAy9MgyGC5JH+AlXW374blG9gllLk/vxbRQNcIldmycRQIfxTszqF41Ikyjvhk2f00Eit
xhuuFJOFxw42OcmL5qUQ0zcsT+faMR1taMBwckJNnHRLPRB+IJ0rrX729pDiRGtKKo8b3AdeDEHS
rVAaqtUuKLNgl5wcED5ru4oaj4G+ycddJwWhk0cxqdEwk21dM8WYOpqeVrKaxpafX2A/VF5yp8hX
lRJI6XgW+OblhVFBHHf3lHozLwKGCfFzpSDQUAasjURFJZihhRXSoM3TUehc1UEP+OUcfIVqmZVo
Cb+uVdFop5DzHxh/T+HIGe142Sz1T3cuj5YWevsp85RVjmwCLIfW3kkH2OozhPUakoAbj8RoZKCM
unqMaS5h9CHiBEJaoJN6E1vjJiroifRx7YK5MkDai4co/RxU5r9ohl1buvJPWzXJMQl4aYO/8TIS
TJr3XfdZhfMJLxs0XRKUg7YdEK++Zf/VaqWDd+4Ip/WWtcRZ/GOr0/wMh2UYdGgTl7Z85DYs3WPw
H1Zr67Hv/8gydXBUYSNGnMoE5NBs+pZPhIMJJ6vBhGIo7KeodJS148Ye/ni/T21GIg+qwwwEQKpW
K7oseOTuHaE0wx30QI9RhVb/5WxFCoNbnFfvYk/6JlSNxFHtAGFKdnoE1jjWKpNxRg2JCzSlT+J1
nnB7XFn5mT6MOmdcTbl0DWSGOA+M8zkyaA+bRM1/q5fnHe7ijQ3fRXSu2boMXKcgdSBBi5Ca+Kez
bmpKjtHXQfUNjN6JqWJbdW4Yv1tCL312qxX7leQ1XkZEmxWAfCAHSFubU5i2TihQM0HkOuxvJlQq
fieV28EGbtbzXTPK3ea4iEwF/rguHe75yRJCmRTU1AGh+IPksWF3ATI1WZSugsfrjrYvg94y9Mxd
mIvNnkhvHthX5GpC1FAiZKFKCaUmgWd+Y2dWqXzYyOQLYJoOknVO39QnE0iiX5QRymGjft4Z268B
RhofzG9hljQnybdQcgpffOxtK5+zknmBo7ODDc9uQXRGl1k72CuO9JfiiRPlMU03+WO55bJgupEC
/tXaA/T7v5hHmJUvmotN7cdTt3umFbgh5aiLX3CAMX76al85yGtqwOHerC8syR8TelKQfwvV3xy9
FDzamj52UDkE7nbB9SRK1c10rXj1Zmvbi5Rxkv2QTg5kPWQJdHsX1RrqZE5dMUmCn2+iWKFDvZUL
JfBt4Jg7x92rqW9zgeLowfA9nb/LTdG77B0Rh3v7CdNeFs2rKwWI2JUaqSw0IEqx72ndei+htG9p
WsAzC0tc5LVx6ecHs5LgMY95PL5+viO7qhK73mYtRkKgi3/uZOQhe347WUcQv8GjOvZgfy0d2RMv
YYXBpsDY8gTTmiy/vTJcYslFt/ewn+ztIowQxSBVuRbYKzin7t4KrDoxs6mizA2IrjfWEayTziZc
P4Kf/KNQ0iAPIzzj8hd2IL0gwsLdYNLanq3LXgmqXq9xVqxjS99vCUoFJj0CCN+f7Ip62Z0S1CpO
Qtnm3HWoYRua2axHbctbBS+IjVTN9ksFQtdhqBKEr7l0uuOw6xN2X9XjALCb7SsbxAAPp8JDEDqW
eZiS5C/Y7SpY27KPCnDDUoo1d0fO+GPNDiO3EJ/DKGR/FTrFjayI3tsU0h7KFOfIR5ep7skwQwdQ
ed5eTZ0Jn4eG+5I9pBFwPHsJUDH5jP6ZAiQegxiPW85EGtKje0whV6Ip6fM0Nk2SXr3WBaJfkY+O
VaBivR6TMY2bsYywEm1RnjD9gBTfwSVeESO1+VmBZED03377d+WPrwifMtFIr72ozK2hintWAKGL
UWVPFn3OuRJSMI03PrK+C809mcx9/f028GzBPoBWOnokQlgKVTPmNLvrUbuPdNLrVrvYPY9gPcyg
gCvxospW8IiCt/fKMV222pXh32HlkX9HIsjXqjoHV3H/tmonpxWZ7kKMWuQo5tmAiOKSTqxObpht
hWB+O+aDxP+SIwGfQS6WNgB0MwoBSyVYLQlR3VsrVrNgCxVc0N4IkJGwusH7/EpzIQ8N7JEZ6bQt
oy1YUTkXma2P4bWmen51TxMgbFLFYe+L+BDKbPO0aGwWEf1BaoaJ+d8J6hP5xhshSUVW8C3+rKcm
fRPrs1vEJ85yG5Zka0MMX30Hny0DCPG4Lb7Y+62QO7dePEhmhI7uyRrmPwZ47Q5QxCngdwvnSZWL
YVoja8TRxPRu7FXoDNHMMq9TIxbE1iA5eRVlpxEyqFzcAArBbY9ydU9MjxesjyzjFWfDKmy5o8Rn
OKKTX4vnAaVvWem14PuTD8dUED66aNG+FT6lnpUIURRCWTQpqoin//eM5RleEKSAEEtIfqZdAQbS
J6tJjnDd6bgU6YuulV2hJXHYE7ahPydxFyjAK0iRR8UD+5uHorUNw369uxFA9a6dqDvm30VZqXS4
pK8qHpYbgmw07y1EHSfNMisA961Xud2ycwKhm25AkdgmbLnP0447f8f/ysYqpO5vV3f3o+dyWYs4
0Ni1M2MSQg8IgYfZlejzNTh+fzrGatvf8RaE2UfBggJ5+FN9t2HWtLmo3gFqw+SVtJGdnPGr44Yh
bhDdXyTVX1Z6pzw9mcP4PnQB/icy2VN8hSCareBFeBG7BimEmAEVIJuOax1F9BwCEBO3YSuqEZb0
aLVHIgKqNY542vFnSSU/Cu8NdT3w1MtnIrsvbbEtHaB1Cw+pn1KbnvjgfRm2wh66Gli0owWclcrt
qiVWmyKngKBkm7wPhmIdG4Mqt3n5w4ZQZ8/FMQ0xux66ISMR1JujJa77xJeR0+p3OOG6j5IDs3bJ
OrnX1UGcI76ZRILy/4atLjoUUOnrDOvb3MhSCjNdmFAgi3reTOrSsmVrV0YHGx9CkMvtzSXXqKMS
U1ncC1ErhY0AJlw/7HMxTaekx7UcUd3J1J6y+djOAs8o/ycFMfIrJ4Pd1+ptee/CBluEXKCNsO49
ykPwSWIJfnwAmT9/V73RdUcMRcGsZKDU1JqXdNH34IFc6d1C8V1Uyj90nm2JoigpuORam/81eeXw
7yvndB//sVo7ekIuqCtmuR3Slpb0fCaAa55f7n9S4QuPO8GI5zkBEWG+oWwiHDNPoScPZrTdfaSP
7GO42V2uwybTmo88qXPAfc17VbVGwIXufLH2afmQVgaqHsMa/zpsO1YVcm+wl2fzhl5Jlx/961dy
maXi2Uz+BtsUeU/NNdq1oROgn5pzsE9o/FJooTSWy3ZIybzM2ZGPi03Lcv9gsq9aEL3viN+ei3GN
XjS6Hgt64APtB5R9hKuMNe7ytpAo7z/82vbofRHXF1MjW0N48ItHqYP+DKkcKXE5/ORtS7UzqEXc
Z/tcBg9gEkFddq8QWLkcVuwAwfBe9pZRIvNZW5+YIKph9WSvv6wP3/VMLm27pjifWQQD0Brkczch
l+J3nPpgZXrYjGtg2ygQWT7lv05Jckv7ZZ9HBrtcB/OdBLDsQZgNy8YUfJVoKs+2zz4RrPJ3X8L5
30Cm+9yduWmwrSvv7YrPnoxM4B2MEVDaBJsOqUPf/8YUIw/8SyZtLDu6qgFmaoIEivkosxjTgbcT
LGAa1YOUnyOIAFUoIwHL/kp7lGUX+uvc/b9mKJiPl1STVQ4H2U9LEMxronRYwwOlFzSr7yk3ZAXg
ZmhoZeVF/D5/71PLg0Xp283QRooxBb4qECXRvxQdcNr8bMnhOt71Mt4PZreYl8sVad1aP0VgZ6Qg
yfgH6nYb8M32L0VbR3yyqqW5WD7cPc5MPGGRRCadfn6KGeGnVAkuTJZVisEtxpS8yv63XBm6k88B
nxTW3oso6+HUOkNjOL38YOdlGKvQqsUJOcpb+gm82sMps4Yo5yfv35YOtY22smvpQPzF0TkoduhW
T2s2bcr8AvrE/24exmUEs6QrIxxfjWTYWGWYtZMvSUx+XFkmIf3JEMKKNVA3vEy9Gm0txD44fLj2
Piz4up5pqZw9H9zTeh/WHLvyLKq3nwPt812J2bONh8MkDfaiz3fa+3JIj9IJaCgzFXz/xkUnk683
thSBlThQwRjRfIOhv6w2SDIKOsFij4whAoN0JpwOOpG2byMLoY8sjsDxrOMazcaCBmvEIW6+V+2f
cN4SGsJTEwBavX/4udNyPXTXEKavuSWg/Uo0eMU3H4l9t+u0QLTeaCeDYHQfuLduqvBfTme87kKf
zLAN2FpYoNlyX7pBsyQfosz8EbWv5VGeyJ/518iVwNFHwF9+WH/e8CM76pLBhfnDW4LJjhlAOjyj
Wkv3HXg4ir0hdBnIk5wuOU14QrDhOhGIvoTYe7RQ7aNtauxJEo3n2XZ0sGsBBlIcSeJFhgXZQUmU
pJY2ux3aalp7z6w+NS44dkCybU9t9Ok1X94FXlpwNfALdxBrJjPPR/T8+DYP9e28+B9ZeiZmhOXb
S8YSQCFDPlXmxx8R6EfjjVVedXAu9R6NnOtcyHvGBWDuZtgm5ldrjDC5YPPFfFDWopJ9HiecFDiz
hjPmBJ2Ui4qFgf4ucNYY8DIA396BAe5g7r22p768zk5g2rn30qC6EqFtgqK01PMcWVNnrgsXnd9F
avpQXjDf9Ls5OOyoWMqakaJvQdKQVQ0ChUfH93yrQpxJd6rZH0/2669SnP8UBzCBlJrZGinpUm+V
knF8DCBucU/FAUIqH9uHRDCjRMCsYxWdXD7LAHmBUam5l74l56o4aP1d93yHEgDwu7ByF9Eb9NLQ
/uBQv15cch+MRWWKgEGin9Iy3OrrGfvzi8OCPKDaIQn1q7VdhuHvaTkIXZqEJ+OFp7WDDdyt3w01
hc8RjHTflvlfRUHpcCeIvjmlG49QeAFidtE9Bke2yu4RdVYiArVFh84eiwtwGE2IHJIf1f+YSyC9
oQaZ+Bbdo1GSbfhxVNumC4kKCoNNdUeZW3+Q/iT2RpPnGJFa1Pr02xNMgF3wEtSj8zGthYQ5pCiR
r40NR1XE1ruTpAtVGfHBr38op/cIR0FL2mk02bFAB0DA1oeBWDQhmewuqP903D7R5AOFZSJV8mIO
aXOpaLvFT/A9kcORf2zlr3DDzb8HA0Eh3zgweMlX1YLclcpoitpW8brFbPwimec/J4fLKPAKS4y8
mPhNSlN/MhAV1LxNQ0W0k08ezWO2emKRIVGpCN+flYsmkOq2fNqnn1/Os2ZBWQXSwtzKZ+pe7rXv
Sw/nCaNctYp0nBc4rksVwLJZSUOqwHOvrQ472ofSRQDklcECE8aHXM5kLwTlXn1Ecp5vpFUsnP73
vSEBgDuZH1MDxaJxAPYia53JIvOlboRjCcFwPPsTSik2J979LkdgoTrIYqF8RSi2+ejvenIe/SGI
vU5dAIH+LXrbNvQUjHO5RBYPk5HhGCqFqAQYrIhKkR9JqGKzlTG8PWmdXgPbHvupK/kufeOh4mQV
5BnB2t7SOD1sFvIS6D6PMOMGaQbJaY740A5/Et8xmAlrt5z0coWw2lT7Sahgd+EbByyvWDs0/M7J
EQt/mguNPu3TfgViFftcidKx/Mt7wDHYEK78WGpOAglk6GfHV4D2Lr4Oi+NdnQCVuKajYsENJlN5
qRhz18Q9ifLx48dtsee7lzwM9bzAQyAuQMOm8D5mRTjzdTC2pl9oe/IoQJ8mdSGjfwYOp1mzZskd
kBxtzjukyWmutJWiH7WOjwtU8bxL6C1OFNLPMzMUEvIKqf+9bDQCFxQ0E2msnk6MaCYLYwORHHbZ
FW+J7/sidaQA4MJvFt/eRNGHv8J7KTLDVOTdI/QjUghI/xRNSkWCigvzbkCxgF/OStGPRcHnXM80
Rw9S5agwKV/VMm9BwKkTSGUz0vGTayJaRDMG6BlX6D4Fs1hnJNmf/wylKVtPYd/2c+5pyAgWwsQS
Q/wQDPtlONuDibnxKW6b2hH1rd/XjcLimo8rSVotuGWjfYHNzTHE9aChh58940Q08gcd8oPHEJDI
vjBA99VLwVKfoe7BSycIM0aAZ2BmJmI1PFLy5+P0FhmiuT4QmAj6yElBWS6MtH6ECPsmdrRFYio1
gzA/mO4J6djdgyhRwCScP2mU7vvaxisQj4A5UrRWqNPcQ7g0oyF2ddMW6QS8cy5MRZnfBfo7QkRq
Q2758LD5g5oW+UooQ80RRYC2KLoA7964cEQetZM6yuYf5K0A0lFL7iALW0SXk+HpYr518rX7H28w
zU6iI2JCaseE48wOqLuRCHv+BrmrBygTvWO4naQqviLPAxj/Suy2A1QGwuUlfypkmi57h8OUqrgb
YBNBNja169bg6hgM9V/EicLRX0/wBYcQd8ARUK5mImo3f1bkTsyVdm9OC1kM7DGLmHHI6ruU+uCG
/S3pE+VpnFmFe4mSTWhJYaxLf9jJg6jViSgLjAp8ks8tmlbxDEcGbmadwXNBEjP/GMqMq+VpKjTw
nBq9x4+Auhsi+svwyQPiw+hbT3QOs1VX4fTUJHVhnCAkkI/UNDEv7wv+QCQs8KjPe2zSahpb2oEp
dRVdH88qmWJYWmtL/erqwzQ9YP9TWFDryPrJqRgHCjeCucVj3nBVWSRDoH173/MQT7hfkLGZlajC
faE8FphPBiTwmZ8yChaG15FMEuGs+ikH/NesIMDtX/0B5gZv9MCU+eK6AiX5adk7duKLvE3hexFk
dUZh6Dsr1jqBUSeOnBA+6D5BfWS1O5gkFUNvLYTT4cRr7SPtdk8my9/OxokRXduwfNiK34MSLfR2
7lDjk+XR3o6mjnco7JmwUyEfnipMYocoz+qnhGZetml5RK2vYLSUWVRB33INJPDfNmjo0zZqGQAB
mv5Po8NvTUy60TCbqYZFAD8tAaGvzA0+X+rrazZXsTbhwMFUur8Xx2II8rjyKA57xGW0ACXgOnja
M1YmPWZvdHmyex1Nu36QeIE1jE5Fq3uIuw9pGRpVqbUEn9FMhaogjR2G8N+N/oLwZkms+Bdi54rL
kOHcrgqBIgpCMH/9dlRSp0aMKkwo2ho/1fWQyRfuAYEw4R9jUgou3xli/qUKzkQs5fVloYm46D3/
V/vVKLt6+6h7MGtTHGCiVF1c5I0YKPG+fmqclghsguXRDd77nLF8Q7hucXE9Eq3sx+d4/u2cS8aI
JP/MjLqI18mV9edt8tK+13mJAp7t0M6HAMWv4R9mjS985FBpoWPO7OW0ByT9FH4itGw9/BRdgre4
ZMSeW+sdnAZzZARDWbLUwk1/vEiCgQTkxRjX1Yuan8dIvndE9eewuK0+sEbOp+nEUJmaogvif1PM
XlmGDII3soWy17jf+E/JKdeXwVoh8jWdGyIGFfPuecms/Z2r0+7xY0lOjdXRJJI/lOvgZHN8IRzT
WI/MXDMux82FWqX6FXOX1KPxSpMIBh82NE5erXx7hPze4PnKhdvCLovYjLTXpa6WC5ALH29UVvcV
KPCOF5Qiy3qJAvnOMNtvcNQA8isj98v+Lr2mrTJ8/ApXOpeN1dMiGnOaatsqIQjP1LWMYZfmOTdq
xTtRG4+NJJ1bZygs0RnvcJ9Haph2vfWzlZblqN0R8tjxmoKpARWhpQVqP0ws0XskZh0smtVtrc1E
XNDBguTGTC/scQwdbe4JKPvOJ1OB6Wwkb5HqXGW3HkRUMY5y595x6PTax35k3mmi7wk9vYMGvE7A
xjLsbHPVqNlzXJX8QJQZisHiOPl8M//z1X1sbKtipPhgKeeD6xrbdQWo51iQTfWOYo86xhLZK6vt
XDtAXAp8/zB3MDnu2BwXrB4yAmATl6bGWKKNzEsfnBxGtkZ7yw6/qvJQOYAceGvHuL9DIo1KR3m5
AypX5GDNFpnYjMXATGOKoqyfaetBjcB52LnItBd+bQDGNI+AAx2uEjkfCcVlmgn7xCqUavwXkqXp
CwXU2fuLeiOL8NOoPBZeYBWaB2T8Py2yXaY+sIH6CNRZMP9VYbmf86ADx0jAe4NREoTVtOC2o1gK
tXRcED3atqWOz1PpPmjVGoG3phJuwYzFbLg4+eIDKhBiHu4fvXHPiO+R30B2yROTv+4fOnEkzCfd
Y+lTTmb2fFIHcpUGrf0OjoCOJ/0oJp9pKiFsZzX2Em8mcciOoeEofd29JLIV0EpyPi2BL5XwftZC
xDBH4vLOG02sqZ1dF6VrBe73oLBeqOFROiumMJZMw9PkU39dpFrX2Tf0DvE4HAm6SmRSka5Opizl
kRYBDknxHZB5DePEzPOK43kdMlUpEah+dtuMprcZeuZtGFp822VbEpkBMD78Rg4Ez6nyza9SeP92
AquJJ2Idu3p7hsX/rXF+wNpzqdf+NLRDfLpYgHqm3dN6qgVCf0llhGYAym9VLOuq3Lb3IwNnd1KY
EjoP8oU73yeQyOBkY++V6IPhUMI17KE4VsUPkXbZIYYQmeXw6JL89ytU9dOCeJaN2OCM6ygHXL31
fORZZIXeI+qctSCMbhD1xW3Hrf6jO0s6AuH0QafIH3NcNoH6UEBSnhp6U2prv3TT+900frBqESKz
goB77x+i1xrQYFFVhqtbWDfFH5uWwyBq993dphGsINbbUffXKMa4gXIQhG3yGuQH/Lxmlox1ac8d
1PGtgCRsil+XmMmejFKNpxBOWXbteJwQOl/QRb5vtWC0ZkCEgjsVSI3PdXHqC3B2SNYsqEuxthFj
aPJAAHBMEEb+myQ5sPkqVnmsCKokgRZ5gH3U8V96YCdReC/5J8P6BbffZrnozC6HHoZsOGxfih8+
SuckglmMNHQfZgf2qz0El0HdgW4T8B/04Ql7ITNdYtmXZZ4BXInDRjHJOyQ8B22XntWC86RwOsoc
h5Pd9NqYW2XxYKdfK5fJ5BWngsy10mzicde8ELC5ag6YXxxNH+e7y6fPEEfN7Bd9m+XNu58WzSyx
ueZcIGzPybmKzGuAaWZYz4zA/Bhb0H6S85QhnYW4cfBzT0dbl6FT3oB3ZHFUzg4YoR5JpspY93dS
Ah70nqw/WPxJ91hOihX1eqWlheVLgYfhhmSIlqDX8d6kaOY+txYJYJ+XLh38TbYkHCVp4diYNtZb
/P8SJpGKgp8x9hoGvsaPq91p3EqpdjLwvvZQMtBNSC7eQOKT5BTZQ/y8T40J3vAse9EYXoDbnQZP
m5IgVvC1La3BDQYDK1RZZUSXC0ghdQdQfoHQfQUkvjKSImisPMa3vrOA6GM8wclf1sfjVByDhZze
K3++ghoOMBsgDjg9/7BsgW+kaKDH4XForgYXUKKwF3owzz7xR1hIIi1C9FwDsaRyCOQylYu1uL2u
VKuqiPy1kO1Dk7Fyt6QW71FyFX4jEhOSZ1I7fg8bvV7YSQaDCvF1juSgZHw8XlPr7wFzZVjDDKbX
mgqn6ezriT+xKLuLdsNMOIulpIjyMpjaJFA8kZZB2dtpYfzr1nL39XzqleMf60SN1RVMzCWxEik5
X/wLdGGNOvLPvyE9tRJ48PQhVPXxv1zBz0+GFAji+aQzXZOeH7MwV3atoxZDSj5t4gkw3FFuwGAk
UQn3Tjq5nwCUzFoAQKXPmBL/icAQyZ3cFF4nQKDUhNbFcAvvBuQqVSkNE9va+6ZI9hU7uMkrEWlg
xAbOo/PeZlJ7u8BCE9twl6xmpXPcObVnc6JTQIa1b2oYaLrZK5r415xKfvQsJL9lJO/y1lBI0PsG
1CBAY4fXcfCYXtFtkHYeUFCFmCryAnkiCw49FQ3gPqe/izb7+Nd5KAv3s2pO2iDLnfDUUunM1373
g+aow1zvgnm/WGgwx2iS55FYt4eI9gs71Nc7KB/yNfurI79nviagFtNyUFUkCIeq5/bRi17cVQGQ
KSa9kjJDd7Nf9YC4Ld66TF96dIIV9k2uNv0Sq6f46ZwASwnk8vCgE+IzUxIbL7BR0Vv5aZNswPl/
UyvaYS9iV0bfxYzjD+F13YJsDHG2oUn8ysmdgK7fY6yIbPllZjUYDFD9Cn6Ynqi2d4OZsknQ6qVV
3tGzFjPjePNcuwVD/TJWtK7eGdEzcIr8qp9GI2ijHHFXLleLZ2FwMhKdJQk5OqlpEl9L/z5TFIDJ
Ah83v4MnrUOPz6vVjTwvpL7ab/ZgaLe1zkxLvVQ8UokaWND+xyHb1XPbjKGHCJKel+MZqD0DuLBQ
ZOcZMc47PcICPaQo6cPdrzv3SIFXA0I2t6dBNNOBGCSkgUY5Ewajr29jfgCPBX3KXfxV4KSQwicT
DkkSm0M+P64gE0o3ETNCQmKLSIw3szALT3lwtg95T6Tx0V3XE9D0DjiIq9Y4DToqOiFOB76BG8Bh
FBuzlW9d4r0oZqQzGvR0UBmZSCyO3aRIw4yU8rVqCVYLAaV/G7vcPhxHvA1XLhsVWqH/hUsVTpwt
nZVt10FLFJOh9bbRFjMchJniE31XJWG28g3RNBIQhqoZ3+rGRI4+Fq+qwFlmpDhqzCNCce7qSFmr
3l3ALkvNTjf48kIc0oYKMpSsEYUCgHFrqkj2YWehW2NKzuJnH3e/c8gMSQYijXeB5F8SnmNmwxAz
wRibrP3OUderJIM8CkpwB+M964JGlwn8RBjPjYYe4Ut9Hn8rJWRXDqrH26DvbA2WnHeUcUbZiKIs
9YS7RuRR/QtwnIpTVATwLZ8aNG3ogbp9BqTGy/Lpj05G13XqboZ1kD9DoUfCUfiUzWaOjRG/nE9T
5lR9H8rJhOozonbb54mjsRApDxV8asKjSgLuBr/SEn5k4y0FFo9bP5HMsOZ/7HDo2WYhqUkgGVjo
8/k/jv8zjlCUWqP73iLMrHKuDtvtu8sgXPG0M+qc4KOlW6xMm1a5MxMNqv0xlsFKjzgPDxso33Ms
4v4RlnngaiKP5PF55mxRaUqnAxKoIubCC2kUYbABSkbVCDbey4BpiQl+3MwPsiFmmkpIvBwamRhU
5ayyc3coqTLnIDHa04w7WTS20rSbuSzQVGTuRJtgC9u8eZrVLlwUgQeymxT+8Qpt5OaCtUAhr3rg
Fh4J9KCPJHJ1tbYQKZGjbJiSMzg9X9mw0bN2KB7hAMo7Im4n57f+av/G59wEjj0Kn8N+B+/NjjBn
xsX5y6b8NWYiM/eD1R95XUuCx61LCpU5gwMDGFemFbOlUDu2zD9+tl5FSg/ZQ85LdomOQiEp83Nt
VweuAAkfy8HZ2BiOpzd3U+L7rwgWjYvJMLXZvpR+ydFMpzVxATd0YYCzaxfhX2SJQyF6fDj4VfBr
oQQMOFD4I694LKcfYjp6rKNslJHRquhx1wAPD1J2Q0C2lezZrXNNQb4q7VZeYUzBkqrZ/LURacuR
LXBhg7un3oAc+4fehmJZKidNw9xY7EpjiuO/jWWmKHGryHFsXoLID+GRINyuwJiouKtBfebWkYUo
OTvPlVlbkplJfgbiKNIhxh125oWqbirs+OI0JGdKmKPFHHWeunnp1eSVhApXEv/etnAgTA/LQrYl
3gFV+l/nvO4qYWkAaDEg3yATFzOjuFt/TtBW/2P4/dBfRxdZujxQ5DcGHyLbkZyVbt2fOf4sYZPz
l8VHvy0UC/6Lo0wSZQGBUh1Go5oL5dYrES6Vp+MJoFsoB1kVAs8VOvVbHjLXEk2qVLkL9kQYd8uu
i5chOCBQmjRqYwWwXnxmdawWsL7sGrdGqlOYaOIjaLI0NTv5twy9EJPhkslE1DJkFFYSfK7h69aQ
LTXVI4korZP80IMu7Ahs3Go+uWOLgp84hkxZUvBrPkcHXwbfRX1J/Kmu1XAc/mVHQeOatAVj55J7
uhREWOFXhNKHFHi5fq24b6f1SddjOE+azb3YXZ3iKCE19lIHQoZ+ShbnG2dxY+vN2PfaPJrQDeyq
sr0qMeTATlt1KqTxgRp//4sPzIqtcD5YUS64+2UnqNr1NIA8nYQB2NJzoLQc43HtkhQWZhk0e8Al
2cOUEoETlZRv9vJXBA6P8v39+MgedU7zdp4pKMHF+O646bqzTs/N/8kms8B+C2Pz8EiU2a+3W/lD
1mDniLfZgWPQssCy++Afzs9ItL5b0jiSTfTDEw5kqoIFX46YgPqgpjOmzNfrz4aDNJHMdHpWBgYJ
sRJ9fM8UFVKlZQiLNxLktz67aRcD+RE7VHJOEOgudYj80Vz6ANqXvBLcNrUZOYgGLiDaJkRiuUXX
+XGDQfGYnO7vSWk1xZSfbvzAp84SnZcbTPxLJ99JdSHLeaulEP1+gvekyOMYSkFvAMyQAVX7eGwN
RPc9yCSVBrEmMKpAuHN0H6QyoKpHSwJHlIe/XIegZ/HtxpMciFC945w081OMkO0TkJKnhZg6BEmY
tabKSM0PXJE/5aM8TYfkNu0iG5miPSZHV5lphvZPWcJ0o2++CAv2rTtJK18/3pTzUWgmgLFZtVnR
nDKJ2N7tveS/Ime7RaZUIDlSDs1CDawbZsVKypUocsic1sgxFUpTpABtQQY3Z4EVmI2wlNN6zMX1
5+oWEFICg8b/biAnJtM1q+ee/fQlGWdf83d9sRdPj4PWHsrswOaJa7dBDGY8R/RFD07qQEbAdgDt
1bXPO7IT00vzKgZWUg0p1CFhqmQcJ8uF3hrmJ8JR7A1L8jcxaJBbBjl3alBBiXCD4gyZMO/0OP3Z
knBWPrhmdvah26gnBdUmZrFrSj7gtSNI3+sQdwHbymAbk55yc7yp4USOIZLqOLzJOpz7ife+8H3D
aiFYkT77+T3f4S5YY5KWN0Nkb7dQfiWwZc4ur3Lwy8jbuIIVtYurArHNApUWi7EjBF/1asF1l+VY
IBfwImnP+qqgCaelU9X0pdcJS8RtDrS+WFxkN0wNtCxwJLN7zCMfy1+OEhKCUFb8LRWpdZTh0Yw5
x7GFoZQsiKy7gObSG7EuGt4MRe5b6sFozujcRugoSmDSx6dW9MSruhQNtUnNohZ6DEDGWTV0leSn
waMnCk5aUR56SX146vRVakFKoxaEJpkpVOpcVYwOvo5c+UIUJi/SbSzpXk/pNlpv/nOckfOtuGu7
uO3nykcvgAPwWt3PfQpT/a3/q6kuG4TzksfXc+U/lMSSPbiGu/6I9krAklO8GdjWgjEOO6eUipz+
w1TJdCwAzoNOj1dJDrRaQIW9gHZKUK8xFLfOjlgP87IthoOxSvZ0LXsOB6wAsZb0FYkbeHI5o0sL
xe/k3vfX9pRBGPlcqDj7kdlit5vKKvhq5ytu7ZpEZUpCBunB3mCLvz+u/dq5Q8YVhV5duPaVkrek
vAyU5t/EWW3bhwUlHSuKM/TVWRTLb2Vnc4sPRZhPTZ+lccwL8cQF7Yd7BNauKHZ67D4mtNXeVmfH
jOmyCKRs+JWsuFrhPtzIJEeAzLQs85vjJHI40N9S1Y2KCAAoypOYLxBpdZdsdM8LeIv40Wh0QJt1
bCQBnu8npPL3XGb1xR53McpikgK1lxL+C7KLaC0mFjHbJJ+kaBbA542eR3Nd4t288lKifnOQXVxT
ivAEOcSaq/Gb4BTjZDKyCRRADh+DvHAIx7y1FlRuPCsKYw8p1bunWya/xOg1tkFMpjBcesxlmIbS
pkeOC15wNKZkxz9RLeZ1R+OHCVRAtODhsKzi/ahdhECLIvzs32SM6dsPnUVWOn8SXuNA3e+AVi8q
6xtfjvy3sl4FLESD5elydOVtjZU6TtYifOOtwXs1YxWeuram4jgPbPllj8PKMRe6B+WwQM1//2Fv
6fbi09zFzDcj9ztU8g5DzFazRroZKkWv8LUAJn8osgj//elwr1TvApkj8E9kZq8DWEUbe8+jpI+Q
G8otDv6LtsXHnSCJhKHrMdU3qLl8X7En1upgtHHsaUXdxKfPBYX1O90A48cnpsH6epkaPOWCCEms
Wj6YU7NnEZX7EDjXP6fo2ES+kGHdPTN3tq18Tq4ET8884qQzNjT3XfuMJutUU2Y97YN9g9MQW+R+
yd78TW2DgrKGSY3cL9wEzqZmSqzXK3yAFs1n4uvgDPzC6XFRDSlnH/07fSZejQI3V+6r13j31di4
BLBGEQX7fr3oXd7YbTVQVwQ+qtpbf8/PD3hsmEocBtiCfZjSC3mANRoMHEl9ocnOYRxoix4J70xW
+GJ4kWcUucskR4XtEAIY/rc9YF6Q6g6bVV8zG87w/mTTNRKQHl1/5+O4UN5PgthuAaChupi+ir6T
SvGuJph6aD9E7a2HCiGXHjaf9wxH8aF55oiVanXeDcq+o3xwuC4x3Zo5B9TfZV03juUsfMSLo8zr
AWFEYdSl+61XT9J7D7A7GCW5VR5geOQZ6TCmwzMveDdzYmoY+5BqpIT6k3u2Q0yo6gIpY3oS346E
QjDHO1obMYDYW8ruhVURwIOa3KBy+eEP0IUfysLi/QocF77e8kag+5kYerMjQIlXR9694+W/QBPC
2GjRtCWqzB+qWhTEkE3TCZjD2Ua6da+RBo+BUWyWLzBuaSai/tkjfTpfg+LgF+5sgOEeFmTqa5S+
Y58PbkoWGU+JWn2vI2cghDoTYGsnO+R8mK9GQ1D1sy0VDJwiBj5h0ZYdzJxNm8d1ltgu3f7V9Ynx
3Pfzi0gSbXNmOnjraN1QJiALtPwBjrT7+NemL1kWmU5m68I9tM7T6+nZQvcS4oWsCp69FX8nNfyi
H5MsDX7K1W4NE0MjyTEbNI71oLFVtF74KCdlL0eYC85UFxZKVVhOjV8XJeL3M6k11AXf2B/X3RnA
KlNC5D4Z9Znjx4A4fEO1R2aq8lw8vCZ54rDI5tq6R2iKlOFokSHiLLNV7XC6zS/G/PcUyxO0AIBx
2VAOzkRpemuQNCkvwdaL33xG7dK9W+zoLnrrwtHFvD2EUmf5RdtdU+fmi5SCcWF6cAUo2EOEJ3JK
/5hbknJrC7jWQIDeN0dZBrSwFG7fXZbSiLPPN1NJVIW0M6pGEERP5RpzuIQZXN+RwvD5OpoMuEq3
r9kRcJo/oSMrIZGKTrgFdWuABLTUlh5w5Tyq4ol9CBgZkGni7DICQmWC1eStkS4JpHZ0zM/JCAU1
I5hc6SmeGpap6ZhSu3KxpWMXQ8o1AP+1KHIkvrK1oZgvbFSUXBNbH6dCCNrBMp4QCWaob1oNan+P
tniV9+kiptfDJbZez4kYR8iuOEASSY4Suv6IccuidJSGOEjPMU2XOGJoGi8o6G9nWCeBi494l5q+
Bv+CCse0ju9zrAtGh27HSBgXtQCvT8/9OJXJPTg8Y2spImA7BC/R0L6+JZ3fNKgigqLytGBb8oKW
Ad+6sccntMZXTC1JOHzfGLBaT40ZBuXXgag18v3PhT9hO+B5B4KSOZp55+rsQxU5CpPlf43MJekT
YtbanPLlddGpOVsQ+7sdMT3uCWOr6tsJMn0FNEIokFHA1aVBpbAOX9bcW6gB4wjhodqcJ/NtslBK
YBOBLwNKzL5zg9ZfhuzmVPA+EW6VZXyezk5Aqqk5loTnbIOlSvpuhzfPw+AJaija9AnIVLj+7njx
fBoppAYxjtfmA2o9Q6me8BkF0SFEKc+aoxiOtn12hISkcsLioo6EtE9Km6xWslxgWXKFj6M/+Iec
lEFblMip5ErbK1tbWewmIRHwZPNLnD7OxmvyzwgJ7Jdoh8C3+RJ0GqNV/19OVC4pjX+wOJo6hBwn
RBNIilJ7muVv/1cvxSLHgsH1oZKJ+rDAdPiY7Zo6er42LHwN0rRYrXa40bqmveCY+EFLHJ3Xj0TX
r41M2JdQC7PdGlp6z+EfjzFSxCAXWo1tTucU18MnaCE+L4Y7f3Ugr0oLL/Rygiyq0JtSu5QAtAmA
ZFrCpnDqggdmXe1tFFuWBVHLuM5dyBSXMeSAFLj+HF5ApipzovsDwYouHn9rUz2XCPS0bhMSRzID
ohuT5XprEYR4jC66Ybs+ypOHaI/XGyhIVP+/ie3U9QK6ARS6gjqNFQ9OSu6Kgb3Hz1PlA5V5zsaK
/5YnDP6rgN6gs6E8G3X7i5/R5qOA4tah48PLV1COpAjYMKNcLdgo5q4m/ugRN60W1oKkC5sgGaby
VyJfK0aIPHQ1aMMgGIOvLtgGdGifmgG4f6n/HpZ9IsBvLobyCdfHA6P0yrXx+gsmlBI1DC3BAIOi
VC6UMHAjne77Mr5OEzV5X6QTWPxaA2TGrzt9JvdieVYoY/8dWgAMUQ6hYBkYJogmgQEyuY3lq3/2
JZeXsi7vTza50GrSusTPGy5fGCRkpDzlvHDHaYZLAyXhyZYLNgiq8iXcSsCfg6SxLUbPumGcBvtr
a3pycMWVnWG3BJLHdF+hZ5Bi9ttAg0VTYVlMtk3EdG0p6uHPCf7cG6LZDwS8eAFHdf/ZkFaNrnNE
Gy3oQHEvpr/GwlO38Af0L1hpLXwW4N/qPStrZUD3K33ksHJ7IIU/5MxvtU9JWhI1ID0n/hb06s8/
8oZBVymyUm7HYoDL/tU+8OQCfPNrKq7HsYK8qpLh9NpC0puVnp5U9OgJdLP/wfQWplTBDUU0eyly
ModMwX6pNyXa1Vk/l4eE+FO+5axcoc++nWEpNF9LVSUOSgoWWcDLHHrZB/z0z68bDTpm+TfvG35y
De2/CnSZRblYJ6IIjeEiG6lZkMTOgRAFZV39w6UabtyhzZmJfICQBfAggDaZHZEAEs8UA46FW8BZ
jVJmK4EmhHT5JpJFe12j2ndNmBs5oRPjl32v2jnvhDHcfHEsnE3zNN49jdS84v2yj8qzR/YuPPJ9
fdQJVrRNoKG+9jxtWGtQ3ilZZNyNgV20QbFlXM0dvSaccDj53DACjpy1xCmHPtabm54ylqWzfLbE
HDeCRJw+JHeP7/gVREb86cLTnyLj6UxywxdFsCUXoWZD5NpiSTMMo2pjjd4acAKvnFJfWanqDB9i
wFkDra5B4X0bFb7ZC3VN4rbwutSDk+BQss56RgS6cC6OTYGObDExfrqmlLQmoP5DP29V4TPtzGTW
UfpefKsNOE1s7Y4Nhgm9ghFeADLAr6DT4ooP6YzmfJKKhiLspSVsACvBbIRornG53lfE3NHDmZpv
65fTJg5ld+mQp7hj1wu5ffIQnbGK6Wlr8uQEKeI9qc1+dtAlye8GMYvdc89/a6BeDWtCI8NQ6qTE
H3pd8TKSWf8g7ZRzq5ArPeLp6ynoofZTBD8GYc2w0Vhe2mIRawUnuPnqWBBY5p38+61n39Ara3gd
yLSmxxbtFuc5HXBJyp2Yo5umZLs9hcuWKVgBqr86/LEjQkwSIy1dvKOwiIQDoIp5Qlh89WAC2McP
Xbn4SesdEZjT60gr3f4Gy8ll8bA5xEe+vyKBp2zCLUIU9OzZ2Vb+UVBeNYfLuOzM3sJM/jPKqlRH
GnVv2l6NxmDymIAW72rRZbxZ+5sqMkCO3NpwJCBu1CSFIuCfUSI/PG86k1X8qP916YNYsISipNfb
GTlaGy3zXZWYO4WJbl3Xa/1eidyrtEOcgfYFl5/rMQOECXbqgPvUlOUQluPuyuX9SswltSw6NNFs
wNBF3bKf+Z+Pk/cOcie75jlAOGyKSA4jjmCH//bmzPLf7WRyTz9ByCb5PX1nLWNXSsq9vOiKn2ZO
iffWlwsin0bdrH4mFfn9iO7SDCQ4++guaoXvPGoUpksh99vhE6iZS7Kwr4DtbMBG+zavkQTG+A7r
e8VJs9aqOnFrc6HF/e3YKS3b8e9swZ5Qqe2OMydQnYtq4jdY2iuT1qVSsYILyykn/7DIKspPjdre
c5mkjEQ1/U5J6TUoxdKApUISPU5aP7tH/+U9iajW3XBBbR//eyLBffljALsWIUPMQmFHZro4VX+j
sGT7W0GtlvxeX50NUvsVmMBZG/JE1h8zLWbdorRFUZNdwO1HgBKdAnzucKlGx5qBgqDZP7X9bcYb
Ad6Xx3WaFJP9L1S1Uyeq1BBPy8/EyuIPiQGxbXpR0Q7YlcYT4Md7avcxBofEHMg/HtMUzjIwFjGY
pyifQny7+gzOmSY8kairZ7/eA/hmX0ADtCQPnuTaQMqPugLdcvz5Kg48UIOVYfoP5hp/yMBmz+dn
8JUiBqwKziXd/DNog4p97CN3P14Yo5LqY+2hIqRyoTlo4K0zt7v8oETIAz4OemAXa8E2XdBLq/Xz
ECvQr0PkdUtHEm9Feg3IT+RH0MRMpM7c1L6WC2ntV7eZz6yoVDnYroYOmu9wh7HVNZgPRRE+X0pX
NMo1mUAb0ZrzJrcDRIAl/L4cFibVr+m3Nx45kHgTlSDdoIpguNFXhM3SxYm9C8KHq/CVJ/jP9OQm
CqYlpn4HgYEqJvP7MBSF/AlbqDUY+s2jMRI8vGmcVg8JhWYyKr7pIIdpWZ63gsucLfaL8xCdbCMY
xfO3A6qoesxNjDDRfTGwho/Bs2oHCswuF/9Cz0dN1mytycntz2hNEDCuq2+hnRP3MEinj08z34bH
ZiHy07FcMECN/ulGPF5um23FeN/NER5DoRuhwN/xYc7/Os7ZdR1EJttWiobHnj1C/9sXyAz0Id/7
0YUmhcj4hnbPfQkC85C7XVcx4zmYUJHwCwT/EO7b0dJIdHQf7vW29VKdRQMwL5ibabtDqbdofLqf
Tp1oGgucn3B8nqc+ir6gigQTrJxpUzSxsG2QM3XXWbv/bdUzhdNB1Hgx2S+9QMLW+3dvAo+3L9z2
/8/D7UYAfyu2KrHC82WWF9T5aqQJtn/m+KcQvG6iqlhd+ix8Tiq0kRC5P4fieRb7JjXLBa6HBB8e
hgBbWTywDrkPazq0reutOMKLtdXHOr/opfYkluZzvEk+EsHjPJDVR23Za9Og1nmlL2wlqFF5xuCO
O5NUqUijRnsGd6bwTyHmvwphaqy9io60qdF9MUsiOsf6sFf79+1vntkxGweL5gQgT/ans+doXa8E
7Q9kQXns0hQw3CTcB8fcKyvhNXs67VJoByCZ3B5p18sqF67qr40tejPeF9ORxDSnag4I6e2cSzjY
K3mwff2a1L7LZtBVc+F1gyWGwHJ+B2BkB902AWokfk1CogV9gNuLaIz4j7FQ0lSEQcmpzJkh9Kbx
oeNCcQMS/NNyZCUKJOaCrCpSy08D0SIEBRsFwMDJ4e00eEd4UUlP0z4so90GTPcTOE7nl0391BfF
41DkDNsqJnTh4uGVFhLRAnlDLr4qG0Ms8WqKHdF1HgLXW6d/TpjCj31Da2+aLBTxjlxhb4iDlRxN
oPIrpquCwenoZznBMoCi2oIHe4v7yaNEzevEtEEXSbceyUPl9OLp/UwV+dS6pnO0h/wszjf8950F
kxUjprwUMWoZ8GXA8HPnXdYKNiZevllc8z/x9s3y34zJmn8dtNe3uCMOyUgetxjoC4PQYfDs1qaJ
fcKDj4aJX/rjuCanxF+oGq96DkXyqK352TPJcGeSV/N5BYqcrx1P9YeopNeX40+Ct3jSR6DmLxmo
/ne3ZjAnU5YwvfMGQs3nwCdM0vbsJKqwBjfuHv5ZXjCL3AltDD0PYzDlJdhUljHpQ75MklQvF+op
QGw6QqWo8+EsqRi48m1P+blGa5QH0T2Fmabe4TWxI78eH7iNZlDleD8vK/yHlAyxWq2QenKaqrpc
GxrYTbp8OiBkbDHF9wsZZmU9siGif/8Lk9uxfITFa7VJPQr9COqG++f2cjg6G19ck9XK7CXKUiUV
A/X+M2dchEQzgozNUhOcJnH6yzRdYfFZmwTnk06xk2fz2j6JU02fDHeBDj7n9DNIXNdkGbWGEfT7
HKVrtMptkY6aZiQeeV7qv/ipEaSFE3m6kXR45RDjf/qdI5Tk7QX6SJ2vJAyRhCAzKnt8KWXsy7pO
3yDDvZ2bSw7S60EC2eLUBNgKcmD1tObGnpGACbcNyQ8uuNFVNVwj7TntPawadxbJ2gXwt/c5VXSS
cqhoZBTP1+AFfD2Jx14aVuYXCstWWODg6MFgLp2uW8U29kiiCantXTJ4o0Z4PZP2SAQYIfmHRitc
zsY6we95lwoXpNvmC/mAvYYcIC+LtmGiAepqTRBuZjxm+s2BN0TUMHJAZjx1w5Y34fgDUiYFEbqc
59xc2Bs2VLhotq8VbRM9wYY7qBsBSQZui0D0fTeOQK2OyV6Bo+vEfExahdN+NRBk7cQ1FytCG3Bt
3a18d6tQ0jASUtjJjjJeGOxa7A/BearrBhI7ql6bsPiWntir637mhE7JBbPslFoipP+wffGLrTuy
P8xhXfO3EpdRlrRlyGiL6Oiqrfd+ikxo94Mjk1pjUh0fpqjhUhhuKiScKgyTiGbwbESn7iHYtP4m
L4j4WxPRv/3WutdzPKrhlPaDYX/nPPLqvhD3ucev2FRprhEdP/Q9U83lIdt4NPO0ROFq5KVxtCp3
AlHKZdcyePBM9UFRzZJWvqxUVSCqZrcpelEN7mX3x3MRb/zjRDCFH+uU2Zj9vYkxLxXe5Qwrpz+i
V9hAt2xbB6xYF2EW7EIYsfxLwidB1N4+2M4r3x0+uiVVOJNaonA/1F+u/TyxYbOC2eb2/gPWuXfe
9ekha4hnF6QKpsmPYxeDPxJO0rQ1ptK8CTY28wYXn0KuJN0lS25KTgPdD/+0uLm67gIX4wRXvFLB
JQ7n3aCa9AaBYAvMQdf9aB1gKe3ctfHD6f3Y/YBGD0jKksKKzx0EbCW0JajF/h8jTeaL/Z4IckZ1
wpTQLBStsV0Yx16GhFO3ccHbjd02SjiFyUyJspuPSUDweMSj1LMQ+8sF3B6UEPlrvUeCepxDbcjz
lzjtANBZgzGy9VpBGQ7H7iBvuhNP5s6lTU3DQ0tKAk4nBlk9TRmDGJpcK2r5fwHvVcpcduJzncCK
hMbBfYW3FST7B6QYK7V2VSF6xp5rEoapNvd5R7y8Sun5sntP7IwXLN6hLDBQjoWGkQTJmZTI6Vrh
yuF0iU2OMYmAcU+e4XHMQkcBKw1nHUe7SAAanpvcl9Mz1nHmcSDQvee9U0ZQqQr9eHelNrFBhL+t
UROkCF/wpOlRzrI511nwhfFp9x4PjR+Xsqe5AEMA9iPj5WE07Ndx7VDr1SJ6vkNrHUTEg42eoMtH
qZ7Yr0zojMt+4OB9wwFZQapXK76OdN7+SGO2n6i/W/8vC1kNfwzRj5J4dbkTGRAxOB9wte3aibJT
LBC6lCiAZPbJ3GdNxMwrF1dnn5ASnoCLGmTQd6HifOmul5I3zHTPeI/VXRI+BIBX1i+uZC1GMPs8
b5u21ofdVljaJEKCED3LqBj4I1wqpVD088jOLd5MF27eTYIFh/eOWEN6fKncGdr+B9gI6PpygwGT
Rf0rq9K1w1YrRDesBc1KPfR2XrouNgs6PZHxTuDuFOPpbrLc/y25j4Qi50xRHG8u2qi70/cyvAb3
Dc5kN4FpHvJewdeCLNgnIJseK1PiVNeo7oBsznsSsifLQMFsD9TDqXavtuo2TxECJfMOE7ECoMwI
KINaXO3gU5w8r1XmwSXVHBdSWB01OiJcvwVegRNjajEqoAedrFrHWR9EDT7xJMoVOF+Rz2abJ/Gu
xnjICtAKZa7zimK14gOkYOUd2iVHj9O4zMXyy9kJiUN/xHXuGfCjvlNUHdy6Mw/xpbYAgdsuwfue
AEEtBPii+tIByaw4TXAygXnqC7+wk1p4TUgRdjzm7bsg1aI4cNBCc1iZX89y4WutIUKsYn3MOjUZ
z8JNO374Hep4w5CSxBQCkfxeITlAXxtHzI7ayK2NmuZ4Hk3fgDPh3VTuN/pdDSJ6YEqZ2ZXZa1QG
TVlvmcjd+lwgsJSZfwCaPQQXTljUv2PstDt/c2qslmatK7D52+2BJA8jdiIi5ugwenE+alWBcKY6
L0OKwmcLQHtLbrT59rmX5IzIeG7s1/LmDZwSIpL5PxbJ56MA/gA48Nxb7n7hoCKlDXv1wBTpPXVX
Kv/xQqr00JQyH8z1t7VwZ2DclLoOGA6g9e8QrNa6crDYyGvLw3dzL0uHNf2G+TZvEL6i7LC4xqSK
dsRQC3GvbvGvXI43uyHbLoOkCRUKUsrDUa66AN+FRcWrmJV4usVu6DcqA+c0AyrPTn2KiKiJa0rc
z4d6gPOY9o0siXfhuXmXda5jlalkPalYSMw3pWz1HXwqaM1pw6irO9WPy8gfJVlvqyE3Iclv009z
ivXM7PLLqy8SMDq0Iv2e7DZXZDAyg3F4pNyGDdrGsRfweLtOiCiDWjQR8pf+7Lpm9Rnlch2vhjDJ
yLO0NE3SzC6o0ClqsxvfdTaA0zBu6Zywz3lGJniJi6kWMUmAMwapkcRIuVzyCNEh9jYX4TW4NS0o
vrE4ovFj1LVkwH20V19g+vPb6EYDXATlKCEHZFa/9rbnFB1sHBHuaeKCuaiOLYDS9wJ+L3fS6BEh
7MZWjSEcAUiod4h2Is5W7+7v0R73q7OesOh7ORyzzSfhpncTRdXc7mLn9HDlRsw6pLqvOtr6kDs1
OQh2LOZmAnMxB70ggguGEuP7bgI2r7K7bF4IVEgljh7qWuRvSYcZKvbwy2PC7pxzha/Iv7AT36BH
GNOh5svcsq7BDUVKk9/5hq6GD0ecmkNfN+13ihZTr4RJSp0A8HTrkcn41RQ0165WidLxOPY9pkaT
wravlBq5OTPccogZm1F2j2E04SY4TB3iN+shZuQs4ZEY++Gp2hUJMUbVByY+MVSmSnTLqK4QFPQI
wtHaz2vHJGwQszTExVpgYecSLGUdn/XV4LKjs/gOd4QIw2aBwo77AKBccp3z23rk9QSP4Z6InxNh
jsXTABiVkARIf/X0479nXHlxV8+UpBicy1tqgqs+vyqjWotaqmr/cxI6TZ4Hq+u9Lm6UwkeiG2MQ
rH9tBEJGhHAkc6vqkZZuwcE4NnLyAmK2VS5/HTgT64DZmfYc+xhjnTgCDXEaueU8SCzBft6uaHiY
mfKBCNAdVcbZcLDUF6RAzqENS3+KcYuXO/GI0ysFhmVu1nyFDnC1P/SjPE8wu6kG/nZGkd8uuvNS
gxoUk6oxINUu5dRoUnuQAZQxd+pwGO5qY25oVJCbhjJCjuqwonBjHBltxgR9JQQoQ9XJz38xJNFE
oiiSthoSRbwfwTs8agfvp0lximyTJnAz+BC5F7bivXQGH26/QxSPmxV9TWvoQIDFrRHhjbt26mFu
5cpoE1xkBRxxIbFshCmrwa8Rt4B9iEHb5l1oCq2X66g6QP7gtL9CIXiclV/yUjsLtlVa3DO8Y1x1
atDWiZ4x0ZxLultgToU7wkpo3xl2YY+HH77RjJwy90Zs9avQdsEv4Hc+FazJwejME9KbhNxROGwi
dkXjFosim6tMfFhaBucVYMcmgcLTA1ZvPJ9v0rDLfWPuS0FArzphRcXC+EDWvBf4edduFEBPBHKz
P3LD8y408AUcNjglreDqp8TajOkVg8C7CiDMUsXG+KAfBSFyylE7w10SOUYhu1IPOTZ4hrng80iD
w+l2FjBx84YWyi4J5rPDLXdzWAkOIa36fnn1sBWWJ2+9b+0VhylhbS9lSQUK9+4zoLSpdpKQ3Rk1
ULdM+PMuyohThH3gVo8MWTViKXv+urAOdTqV/cUvLdAq6bCLBO1nS3r2f136iSDaFyrFdpIIq39X
CASLzbhZiF6eowYA1b9UenxMtwUFmmuF1L/5tjjTXM4PEwCAixdz0gxBzgiPI22drJXgSFd7hiQX
FBbllzfefmiEQFHDKRphCRn7rLf/Wy/+ZLnQ2XJWFhr70JRJTZ4nIToTQ9BpaoUrM6fxVjTbiaWI
UsIhPheX41aMIYMh9nsxXXax3nVWm1YUa6aLimYvbW5t9plo5k8zWRLEfvG1+gAr14dTAM9hZapv
3bVkU8jwiKDuNUunjfSVndHcSv7etVuYPfyVMzOrM3TsMi/iChlN38+RLgJ1+vdK6F/8W3SUakCH
n74nEqvPW4R/9yeQpCHJPrSgu7Ps6J0SaGoC8M81Ho34AVzDkXI5yfBQC71kYMHj8vHZEL6putlO
0y4VLFhgVmM/8hGZzZh8ltSGPhzl4qsDXALgWhYbv+oWtr7TzobEaICutG1lcvGBoaojQzHeE51y
+t5pav9orElDrqfZ2H8HiI2Bgym9HnGoy9QVFuRa/DZvk+spbE497EZpk4ULvhUJaoQQko1oWajh
OUXJ7jzA9IKQ/M9mVmnEYep7wK5diUfcCQGZewYgK2L+toGqvd3IzVYYijQ+LeApanQsmUkiLJvH
U5VHvNMrcCjn2d+hJT0I8+kwIG7m2S0un6J1HzurcxldwranftJfrg99dKPBJy9t78AeNT5P4/fk
Q8QkshaULt0KLZN/lgz54qdqt463mDIvtPaxU/GRhrwQFPt3zMcNpk2Kda93PCfvDin7QXPH1zdX
xm2GWgLjb8B6M4EQuopUxVrvEP4VnAKh3QTcn0TKf1L1zghgHZvIPIYeqGJR1bi2emJURulJlDB1
+GMqo8RMVJ3r+Y8/q1DQZak+/RQoaSb5tx4x6ImQWC9SuAgI5WhfzkbmttQlBrHCSiK9TFdjju/f
qruY8BsKdcPwoUNXUrvdGalmaEat5BB6VewFnAIPSSBxCaoFJG+939Lbi4Be1rgxXMl779V45yt5
zg3FvKop3rReoG+cfNfcFI8vX6O3eqRCzpCClKLTzYFer8sxIbEWYO0gYhAVVZrmmMNAeHRLqRYe
z5RDBO5PimA6FpjniDUiV4Uusibn8Re1mDcLBOoUtIv63AWSRq793OQmm1hJv2MZ58C/1fEgCs8Z
WVWSe4FWiYSLbgix5UIMllqkdar2CSe1WtcF3pgcoABNjyP3LpJvmy39rFVpU12i+F28MqanAoQY
PXuHGxy6t7R3aOed7sHl7O8Qc6nbDDt2++cQcaYC3Y/k1CkIUCtEcgj21L5zNt0ORXzy3rg7LGvL
IzVhug5WsQWocch5Y0Vr9xFmtlKLFh4urJu5D/3TpC/FlKAvUp1Z7Vy4G7T2Zp2N9MSq+c2i8ix6
Dl+7/3qYu/PZs92fP4zULqdpFAVf8Fs7JmQ38nHjcIQYXSaiaU6npqjkMjzfZSb5ESyCT+ljWerk
5U2pw8FVSwDtupZRm+ApN4qcg+bK1QB1gXP3fwCwQ4dJcR7TKFGAgu8Hiip37B9PZ3lyui3Q9J54
2mHILuDVNepEx7TWqUOP45tUi/8DHhdiUXGF86g/fQoWLwlM2b2zeazMcP8QD4SxMa5qXrVThQFV
Y9+OvHyHuQNqoYm8St4kAy5k1XSCAtXETpHoojDAFRcN8nuQVntb+FlOUxLio5QcvO8DHaqKjL22
hZULmajQMwQabDCxVYcH1lUW35hOqVP7se2njvoSusipKCz4QO46qvqzCk4N2m3x4Du9k8OKPZn1
PyO58G77vVPHABBw2TvLbvdhbbN6i/FU2uNeFvNarZc/id9pF31wWuItO/UuO1JwtS6OwUVDZpDi
JUmBSn1fpvEaOlWlO8OII+bQrXJZakZpQfd2GyMf1OK56HR8Jr49XF1u9WGnVrqqHty3WJkJxGpL
Xz1TTxmiB+DozH8atm3W8w9eC4AGW7xzF9zgHHbvOjvTvEs3tVeD0MssjPSbhvDM4g0EsUFFM6AY
G8SagPcJtBkxV18LPIWeg1uytf3SUq6AE99Iqb2GXPNp50Zr0/ZN107CV8huSb87Ox6ARdixmZX4
dAf93n/5MVeRLH0zUb38ydRkrDV86HyPF7pSXk/1cvsiCpnCt8/Jat6ipNZb8M07RO+LTBeglGBX
+HCouWmAo/b7nltaMohBppgR9LzAgeZwO/BHbOaL0eesaXoy7RICD8PUkl5y6pQgkn38VLielG2/
M0TJ0PaUwe5s8Mv0AfJWE9z8GDHE0kkQTk4BXk3+ROn0svCbhvLhUjP0DI3TDz4zQ0PI2DjBksI+
vSTZTpUYB2X9ZcQ0QRPsf4bylaqJe0E4S89eDMmBweptUivgofbTF26YR7oaeBfTzi5Bv2WTVJ1g
kuoLaw7NpHvlPIk+fIrVOarL5huyFK79tGdAnfooRFmAnKrzAQUzEVuaKxwBwHqEctJJXAD9HSOU
A+WP+lTdljzdJwqns/Htc2qmOiuKnoiDVbAZGCFcPlHZbcEA0xi2G6I8T0FLIJF2VPaiGECI7m5P
JWi3UsbrONyekksPraMP+iUGscWR5OCqrLQNVtfzdxkzWkQAH4t9oL6ysan3BFJsh87h7isWxtAO
sQ8ncgMj3WV0DNAq1/jIALEy19gzGko5OgvRIKpCC1m9FETIkph+5Kol57oKuS6+aDwjYSLtTJMS
XHMTaWJR6K3iTiiNq5U+aXynM8+mPhauHoXmQuiAay9QyybtEJ0fn27djhNFY+pvg9br4UVYhkby
EQ6MrkD4wTHPAwU3Jy2hAMc2eTRK6lnnH5TGmCRQV6T4nTAaCZVL5n2v8qYh6BdaMrqNY5aNgyny
1TTR18+L1q4lS51DDBrF+o3wlINV85XEaZ0jnSXu4U1o0hHT0KzJPELiDg5Qy+D5ZZlaYReKn7+C
Qt7Xk+w5XfBTV6MRczYIi+hI3DKcfMFH/7/emPU/5XmwLXC996SIIqDY5zZ1S3nds3X3HbiC1RXf
7dIvqUGGW0La0bjldXbbxN0Dv3/n9u8SKJhliq6o93A0Sf5wJ9gcx3HUdbR7y1zDVA/JDccytvFL
vpRxRnQWFdB5yF9gtrlC9gVFNOL3wAxRvq4edRV6j9rY5tOS2+yyP8ir7pQmu9hodzIIHr6rrjio
TPvde4OvE0Et0q63t64WZGSn13IvSuZdb6al7LrXDforetVyKuODPoRmogrgzeWcrSWj5CZbAGJf
Esr+SMKiLqumIBDDe294sjb4YO4CVDQiot70JQTbo0iv/IoUmxm1E8ArDkqFuRrgDzfq16bADmIk
xwIBZtBRx7ZW0TIgR/bHzb7VAqvIvEc6vu0z0r1bvPwfwc+stLfccNCWc7fYEt+vdsu3qVfn7XjP
zlVOZqQ1a4bVqjOfrNCX8Cx/wsdqPHPCzgfLiynH2AvDAaLbNljX+522/RSj2Insrsxa2HOFazb7
WgpL1WUVX6kNXk1ESyAuE4McdN/lUCoaQDCvd/9xd2p8QH1s4zxVtkKTE7+SUYiLUggRpc6EssHF
6t8GgxhRz1UADljGpD2etYYPEfmB8sxqU5y2eZ9ahrLqEmVshqKydN9TaE4a/+gysvxcn/Q11ggT
ZColX1RVl8QQETm1fv//nsGODNwsc+CqvW+jHvqyqI/B3q0gtbK6EFHFi+PuoQSfrwD7FXjNaXSB
4HHHINBWpJBEpOoAvHs22leOUvFS8B3Iq3ah6z0xiIeeEH2WvvOl9YFibJUoFt7WkdRjy6h3Jav/
tRtBfcqCGIbWRjHLIaqzhxUyDrTo97mrkYQy0zVYclB2c8JQcUzoAtF3qQ39AJD6//DL7Z8CzC1s
hZFU4pr7SSZspRskCH+6r7hgu7z9com8jkAN20ZVQrMnVtlTQkzYIjMDOGYjIHCHKpbS2+whVmBV
oWnuOQjIPpLo+yDsbakIPU8+h0FxSd4XkpyLHEGruUWerFgI7+BHJvBiHKpqcqgnTqU8jOAQQkHO
VjxpcAZ6DDxWnHHRlkfeBRaMqbXCDFodMNHW4e13TlqFZCgUGyjVnOXM2EFbVG+TUXtP8zjBqwa3
EYlu0G3pezpLBvy/VCOpk5sDvoOG+lQejHC2SIC2xBDA8bYkb8aTXyXFAOH8elPa9Xu/UVK5r49g
6q8KNdgNLenGahlDqjSV+/js799JfRIkM8Vv5UAxxAViYKN7KV1IdwuKxfI0u6QUsxD/yOoblAXZ
JgfU60EiYzXT1u4jrByRNo942C7K4kin+3yxJ57GjtCn8ckAxQd5COp9WM/15F13u3YcYWxkl9aW
AWLSrjnCLPlZ3IttOwy+V8liI8vLTkzT3YF+mzq4X7fHZyjqWH23IksnGRKUckVUTZxamm7GWq5M
1RIrVOS42A7U8z4AkYygwAq5H88+2SaZ93IqiPrg2I/kEPpqgmGNsPiqXp0CBnmTSQ5eEb1Ai3OH
Xwk1VsaU+i9WinCucZQGN3iRQr4i/slOL2RFpMdCY6PTKDkIbsT7X/UfFTmscGqNtlYaDJ0Carmv
rT9BJciKNkoM6+xgEVjVSkf+6yMM84gfCEQmz734YjHjetF11lk8DrwRpqAng+SehDrIcJHeSi0m
pUsGLADdDXkiCin3IGKkT3A4426mS0ZMETi4uYFkAQgLsMCzVPhLbCtZWYl2+6zEGk+w5C5hZyt2
QAyn+81dxE0nmMAV1as6pehBx6QN13RFlOc9079KJnoDnSem5pfsS+jkaSCZylZw9WyOM++lzyBQ
ARUTU4OBwn1cNwql6HmapqUqe8SoUoJKjzvaFoh3ApyBU6qMhQwTbyDzunILEykv07mmGgBzN4ho
csfgi3py2mxC941bRbGe3Yvjy9zwkfXHu/1nNytQcwcWIo/HjVx4Ms0c4sc0hngo0be3fE3PLAMK
zMk3AgvAWpTYxPnhizERhMXM+or/cr16QJFj43QbgQ7dbPO7BEbu2Ut4v8ibsYJpeYivK19RXiDT
SHh8wt0O8PvOD7AyVI0Oxa6kfQRmaY8dB2ZypMj9Cda67uDqUqtf4etqHVfpD1RI3Xt8t4/ki44o
7pPmspV6BdWeOZPMGUYUrDkPXZIjp9uW49K8bVZ1/zmEtCUjxGi575FuwbTWNS33aEWgqetu1tos
eRjpiEixekiAQF1htKVgrdB7I2YFO4I98rxeLHgXCwfd1U4cTdKpJuiRS2E88ZBArgSPxr25GJBg
YRGm56xp7anPkTRs2TzRR0uXR7xNuepbBmYjL7diP4CFCVYuzQ+Swu8ZDKy0ulFajOqzjJ3btfS2
ilAo55CIdWuX1QbXJCNK2/7dJPtUObVZnUw2aKzS2T9/WZJ03yW2qfS+MmaZVccHZ7cfM0EZRHpm
W/zAGXEYENmOHmRISWcoodtnrXYwyBrzCrb+kJPMzM7Z6h5TgkuFnzyrkVo0Y6PAPERrTnm3w1WV
jGpq/r9mVHm3aVzAgjiqGa44u4YNQLAuERyLiN1u8OnujaI7wgG9c7K3ok+yTEUQ1zHjzdJZUsN9
euU5pS1jKs3g6RI67WLMQOUH8f+nsFsQM5obeauxsI6HQc+ZPA4HnClFCyWer50zDjplLLToGjKD
EEr2sGMf8+sRHFHwvJSxxpMOZIdHQwDUi9WeNvlvkmOM5PEGVhC3sDyue024tRiL+m2jRnGFiAiu
B3uhfUvxn9+dhSAHO+hs0XTsR2QEjxgmxqP/XOu/5JT4zsnndhf/M/ZIsggqZH0BbcgeXt2hDZ4P
qFyPVwpv0hmkmj1WZasdkTDG6EeBC3MwcJBwpszG7A6Wvb3OAHv603MtH8Ozi7flDspAshitNsU8
BippLNvAPwc0C596cH40roYdteHKx3BqKPUCOESePUkl+VNWuEzepEVboDlCJlB62hlhBidaTmQO
Z8mkWczwz25okvei6harW/HLivliOfVpJ1mazZ2X7p4NEJRXZYT7mkA3Ul1dsLjOC/TdyFmjVV6/
P9ECpdOP7War+FrF/z5fPmKsqsxAdkink3tz6PVmSMNtSbLxfU/GY+NEhUyNlKKHejIKpo4b3JkM
/5B2X8Rhdfg5yFOd5p0V1PNYznjMgjqK4p4veq9HZRv3aJQzNZmE21tSPJzb+zqrjAkqIPkaDYdw
hLuQG0g0fFf/ZuFHoYuD6hr7Qqm8Sa+tKhcU9BgeG2fy2EtlSixjrxHyUigP6a05WwXf958PlR5N
Q1vD8JukdSN6Lc+weSm2zbXMnDkbuG3KAYSqiyF5fsMxvrP1oh5aSuK80V8kvz9Tk5QAqnjxWPE1
aoyjzAynONPxervGEd3T9iNSVjuorhr1KKeMbhvurLJT16+nDfeJ4P4oxNK7PyMYkY/p1LSSoKgK
w/HBLWdNyGjQTJoXA6Urj/rpN+2Qd19kkyPIyNx+3qjOpavQrkisi0fnRm/LJAYCi7VmLcH3Tn4r
j2TGrnSTHJziWVdS7kcGxWErY/IuqldFbQpR5vDIkCNLO2xv7wztN6/MmQ20XR/TiS6glj0riPcR
I1zd6l61wXB/fgIkSphN5Fcd9zVMYc1IRfMRTWqPl2MS+rzoJpSjROq1x2xmEThszBrj3KckJ7Su
xR2MpQu7NG9bd8Xj9KNr94EluEmQOiK3RIV5se2eqYPDlMf1UAVJnupKUFnQHI4kCRv/y2kff0oW
Ay7qWX4/D8+ATtU4AlC3oLaQuKg5v7mCbHnMWSQG2czb8/mvitsn9/PJYOCEIaj6BMGWO2IjccZv
TOrYXNVxylOtQUdYPUjNJj2DAOpn97bLlcrWm0D6fg6eSQGLbVTWZSh/1eyvLke2qJw1cc70ThmQ
Vb5DHoyQDDYzeENFMqPA4CwklfFoXaQx5agqmPIrnNjYxAPSi13720L0h64yGAM1yfbgJqOFQn/8
t9lArF2vl7UjxSS7PkYqRPbKBiHKj5Bp8VcDYlQQDBabnoBjiLZs10IAUN14tme/fZ8Lrki7qB3B
AYbYQQL9hcwclz+Hpjo6Z4eIwWn0GzJoZrscyJKZ/wnRT9mH5f6VMtBh/oNcadJ85L8M5NB2YRSH
WtrFgKcb73y8bXpQLMF3geN+PQMHEQkBhe2vnzNmwuZ+5bAWpN7hZoNTH6k5I6e53saCmx1orzUX
ACR6ZJpZL9j0v4TN3aVgzBpwjAfo0JBd9PRbw6/7O7qMw0gJ3Rmo0AUplsApgqytGEX6QFaYz58a
hVpW847yPqm7hUf/qdd26k6HQQdY12LiwQltkuS+ZiBdWbIbj9QH02hpIPNnbf7SmJPaTCcSm4Pn
nuVo4YPsYNeNqN05JMuoRyiaAIAegMEvXohra/xokLVvDUfA/z8dps9OUHEoYyTv3cWUX04wDKmj
RX6wnRjkdZKdE/kZzcRhbdQjWmOYC/+SExNxIWMAAgniipSAIGIhwbW+8HLH8+80oOIN5ICC7Mqf
Suu5TujgJAnspoiT67u9kVbVqcP50D3IozDZ3YWwDCV4fxBg4rOSFGAmG936s8jKIgv8RzX25MSG
DQA8nYYGsJs7mfGJCQ40G53vC76sa4RGJV547MjxKXveroD2mfEUxDi4rcQNgXO0JeadKbQ431nA
qmdyx9WyzSZSBH4rhGjPTIacQgfIlV6wdcHSIe0tFTUsfWdMeRg5VgBYKtMyzISkS63sTF1Qezrc
+ywJSxGz31PvQ2FQN/TdR39ut1LbAO8jiqaRD/s8IGmw9DqvQgsHhbs1umGH8xdH4xiAGy9EJYQw
qL5Mhbzmk9gIm53Wzuzw3GPMVIDkzGY24pgzxYYHmxKOA/JH9EcFMJ5jNE5wYWCmtS4V/9Ac+lEh
6E6Ftgaj3400kXPtEuZAs2tiZFSgFPxtahIrfa4ewpF4E4LWRb6c/AWmb9Q+Xz2UVoI8yDHBoCpS
QsicWwhZAxGYsh3kurIsbYsq5OpIv3ItejRS33oh8/R+qs4CrN6HxbE/h97k4KE5XXAH7qE+EOX2
keEu8RGwvK/JvofHuCztTzrTO/cVii1gePZZtoqGv8Wu0sPQEwuy0qFWkn3I1jhgYAeGF/IcwHFq
uhaD/9YRFLVUTSBhYyIumAUquJzHwTIeP62S4dx2Q0w79iHpPYTYrP06RrghoOe27AbY0V38Zv6Z
JidJTmqUyyMmnd6gfnGG9FI1nP6pHflZdRu5Vk6XDvmH4aesMZC04KsAZ0yDi+hvBwMl73kMwNJX
/ubzPyapSxnq3jFzB++p0NJO2MXgrGBX82YdUnIfPUa7vgBqDOWNWM4k35wO47B61GESfyrMYYIh
93+x800raD2g5aNSf0/hEBO8ym9iW7cXKmbYrVGZ/K5dZOrDyKUbzZ2eD4bixCHeBQ9MC+nD+Gx9
USGOZR32b1W++yLK8XzELCGiElR5sm3OVosOmobJfiaAWBXPPUjRO2U2V5NNT/68S7LQ6HpC0tld
qyDjWb6aD7A/TaRcC8mMM4kRK2WRCRUuZ4RW4Zo2T1fp7VAZ29VmpY3SGo20y3sxPYRaRvoCMHkU
c0UNw5zxElWOe8MKsMnndDh7z+vBsG+huqu8gENAgCkkaJ6m759Aph6lYYU7wp/MOKzPRDtP45bs
EykCK5vhND65Di9WD7KwoU26hPEd2EqkK4QU3YCrRQ226nG/v8q07HH117X50VrwNom79s2ngEfP
eAztMqqpGkyYH0o7/zZhw+M3dnJejtA5BQumJTae6EppwA3KdN51Oyu6dMCLL1W9tn1oZnOwRrnG
N8+COty4eEcsSZDM0lOycAOLky9gmZdkRtkwwZF5RgSY0LuamjXOrMAhwCfSHmexGFcDD9N9G9oH
PolASfcSTG55mmK1f1/Z6savQmcjSEnUk5CDby+i/N1z9JlbKMBpovxqgojV4gsW/HJVFtZPkTkc
M7ruh0IExo9SCDSIonQOsZbQj9EdTN9Ib9va2T/QpSeRBaK10rWqa+RTVyyHWy3wkGPgnOoJ/aEt
crpu1feiJuwZYEXQFPt0qlSSztUtBfmCoOzTJvcJfeuIYdo0HmJjshD44ooa0Jl46ivOLK9swDME
PEXWnXdZrpdLylLmrrfC/46Q2bh4E9iYUe8hPOCDBSZrkSSxXoxxzRMBr5W+gcLF/51oUPI+/GFj
UXkCHpWmCdsYvzxwAo/lD20aILh8tHzamkgmLeTGEtcWaz2KCZWEatF7ph0kAa8sc4gogM3oF0lD
jWcf6JQSa+Z51HLKMY66BxXAK7oVU8CYqRNV56/9fbAH7Z6Huc5QAdr1oGfp0filejhf4qyLkclu
D+Ndd00YLceh3rKL0zBafRPy/vddweQjZPplpD15l6Wp/+Nbg4k80uYEd4TIo50c1yC3E6thbKnA
46jkSbS1DyTWtbvKIfI/zeH+gaTDAittlQJK0ZuwHpgCcKMk+JCvgr/CCeC9jsx+o7uZaBZr9sTD
y8tHfe/8z1N813gLc6hKPdBqJwN1E63SOMfioGeXPZCqSBa+SH+LnH9a71yqDpVtW+qEchzNIXjJ
xAzw/1G0hNYTRxJJvxdESTpqoCS54bf0uO2EZ2UXXIuwQn5UIJ5R61kjWrM44WF4ZVSi3tXN3MUk
60Hvrg8WKflPAN+9kTO3mS6Cy2g9jLQGp5gzzK5FOJqCZrkIaizIQb5T6nvTx2Hu7L5rTomTGkod
G2RjCOJ0oZhC7oxOPdvu+v+iFi6umdZxaR53xg39/NBhwRXsEr6xRSfXRwfsVYLcs0G6b+ti0Q5T
+FjHn95vsy1X/iR9bqQ2M/UcfrsYqUYLyEifzDhCO3BVz1QvyJXFahtyTk18ofW1ScmckGP+zxAf
97hMonKwdQCVCWuJX9HEdvKIYtEyLyT4lI2jUtxtgt0s3AVnoB7aoQynoPojIFwBA1xDIezQ2VQS
RDlhfVarJFaGnXp5O3e1+cwl7yzdpQY3SVpnm+nKJ2xG2qcIsR8qcjNEGGGaFcMbN/TirT1l+nVg
fxg03czWpo6ro0BId8rDvfiJ/7PydjpBT9ThNrUc8s50IydRcNN3a8lFigKb/CYc/RunIcNtvOFt
bedVv66zqhkW4ohBjdablLt7X5MvoIs5AkkVPxB+7NkEk4alX65AZ1GN0n0Cd6qv7XIX8yMgQnjq
NHUEGZg3oOteH2jZB56lJVRM80BKPLUJC6t+vtrjILvWVpkgqonmZcnZruAhPKG/gJ+FYO0kVso8
wOY9QBp6Pf0zAElu7Z1lbOq48IJk0xz8gemk18yU1CXi+0AVnim+cUcUSd3Xy8TOPr+11a8YA3LX
nJ/Nh9f+8WbSSK8GgGaXka97SOVOIcjGYH4Uyq4tRhqbpIJUGPgLMU4kIbCsHRm0kZzKKXjXczeQ
GpLJzvt/eCmiIuzNEakl4/wyiQYJYF+gSNK0EbYB8aBJqx0khgSU/duWWqmamNB5PpcKjri270Qx
NOjgLTFyUHYWwLpTYb1U9OiVQg1KBNHqylXAiuEJ6L0tsdsdUDq6xqyRHQLJd7/LqGZVfCUmddDQ
PdRbQck/pFQn06/xVZbaI2X55AIUs/NBACfso61Bb3b1W8dSOlaFhrgL6FklNqfKWj6Kb+ZXyBOL
QhZk7VYMBeuNt5frX5AhcVEk5MB7qRWcuj5MGg7BNVimxBV9DMn+6Ujs+WEVVGEffZAT2HFirIiQ
s8C4cerK7QrbU8qr97s9IUcHIssFWHpvzMy3VmwzlEI/DIHOwvaokCZRERBG38/uHwSP0WTj/BOs
/LYl64C5qvSpRS4RBklGIA+YP2myxJUngd2gic0X4DcGUbZN5XtIes1oR//dcaAMaRr3jJSwYiOu
m7L2erYota7B+zDi2l8yDA0+uRzhZ2LJmx8W0S6LQr8/Se7mZS6hMETHtXJH4P5+WRGFj9pbdEU6
YbkNQoUTHg8EsNxs3QK9LJWJVF8hKa/zsm7uPE6fq1g48ZqXEuiVuhHG3q201lbgaFwh4X23Ucuf
7BmIFjMtqT+Djm3g9M5gteVKhuABpdwQ7WcrqW+PQgkdWbCzKE20sAoO5y510+jocq/977z8kxPQ
YGjX9da/kK7cNBZHbKlSOj6/pxIxyjKnsxb/ZuUV389tPNMf+vc+NgROHdqflhJXLqIVqCzd55XM
jhieMDGWsGa4x0/2BLDJHUUF4qL53Uvq5wpndmMHpgqblGym2yBP7JOJs+WvtS+RnFmz4a4bYF1q
Ja7tdnyQB4o7nJUJlBCTaRr2zPEBwm1p8vUSYvvFsx0shrP45+eToXqCzd8rYnD6/V0yGEPjbszH
YpFaGiZnam9Pt1corPo077UaJ5BL/MUUhezv/xuYKDVMZLDQZiAGSwapDecmAqNiFkCVx1CnZtHi
TFUAc8Y5qey1BrW51E/i4v6vP7ZWbdIJxZMfhqwDCvuWUSRZwSQdoC66Nxj5h4ZERBhOC8CqO1VY
fOoZuCDchrdTsnXUjumG/N/f3JWud7pWlTnEilyeCB9GAlcNNJ7KdXPKH2DKCDZ2/c1W39MVC2Uv
rAswYkeK+ycw2hXhAz/Qm8zmrLTPQtN+2HLGCrtl7p9VGbp1ZICQLf6ZPtW+2/yciShEQfAprUoG
HBWwA2fItgcjF8pkPEMqnecDml+i2AHqFSz6fMTwY6/T8JmexFTvvyzmzEIhy3e3bNu5uGb+7wUs
lN5o8IyJjzdZC7RIlf0sYX2wyu4f+Dl5wtM0FGmB0KxC8OJlWi0lJghOtP3/66UZzpX0jEPJInm7
CFa89s63lruR0QwSP0MX+nKDYuRGaLdbZPfgzbciTYHc1qnAEAXdZEPCN4BBGGN7YEgXX8IEJHMY
VCkfL/sCs8QmurpDq7hRDiuJiyad2qYlOZOUrRsvvdwmebeqOtZHL+j9CaZKtGTVaxYySHv6NEHw
EEjA28osRNGCydimE9jfiXQAwyAoYPOmwSyOFZxaIoRkXtxidp8wjhlJGYqhE7HgoWwjc3P6LSu1
9YjZ2LL0Jm6M/VaNmqGRuus5La2pzhMWhpSxd+YAJRaa90+PTH/5HbWG7kMGqBBxJ71p14nGNfIG
hL14gxRJsipafG6DxYzlyQdwlIzUrzU3H61nPW1x7Bqx2MZWmlxXrJj0luJXZjNYDXUQpFWlAZrf
B5vkcH7NYht+7kJ6SlEvLThMO41tlSZk0zj3cKlgTI35bB9RcJaVHYGzLEPc5ZfD60ByZVLVHNVM
piMty6xGQkpbqr36ycsdm9QNobxsjFab+j3ICkHqVMJH3+ligcBFziFONgfk9SQkYIdQTiSBGANJ
+aUaZI1t0J98uicPHRUq9HiTvA7UTXuArw0swkpiLdbTHE5UBuC7tlNYDRyFt3Nxutxfa92bDrD+
e8+jBW9yxNcbcCnoZtkeiIfIYhwW9mRSYHCHQCzGVjCFo4RuYROLya4iHBDz8P4neqJHmazzCqv8
f5beh9r+aceLUJFkcScFlMq5qa06DUFWzcekGxZRFs3EGI3JtoIhA0tJpG4HfGuo3aLDtR/BtqBN
Ou4Vtez8IvF45BBN4ZMY6NFGX+lGqnEdDEc+S9iQFYSW7r/JddgBDoJxQbG9DP0795qI0DGCI9sp
IjfeoRZvYdJMKu6isB96iTO6/2LcniHTgqcydmMN8LkyF4FNC8PjoWNnPV3pUHv1Szu3vm3yhs1E
/d5ZU033GxsIcOMyfx5EZa7pSn5x4fb3NTZebJ4LT3Wfb2aUs4i76D71rNtMKzy1tPQz9ekxHHNZ
BF8ah/ErAU/E0xbBe4345gV2p+BBl1BsAYr2B6xwUy3UuBao2WulF1w/e/o93+CfGxS9QedIarmH
TME4FjBt1x05yYXF0APuWR6k34Co2qgaaRIsM9Tai0vt4n3EBNQ2hhlXoDxd8TCjkbZfrVtH5N6Q
HLub0SxcxaUfiygpDDmMfpUQ6BbkhgP9cgWIz04qKl/OQvjVr5V5kVctHX6mv69sHOEROUluN9ie
+pqYLCmbKHJ3kevFPy0ci48/3UtOKD2vtLbKwyEqJK+rOUrjsc9BHUfOrVbBX/9Icja7m7br0F7+
2RZaNrGtqJn/MYDaFPvDoVB1RVX7k6eHlEP98cdox39LfsEJ075PCrPLmJ8lkG+o+qBO4/pMUWHm
fxp8zkH9JKSjwldnRwFvmMpWngJr5fDc8yrT8l6hrpejIgSWbnBm5rXrCwjwU1gmIBMEP5dRRXhd
6ZtqFfsQo7Ax9iklmBx/WhoHAJBY2JR3RBQAaJpfwsxjpgwCInYy0HLq3F0NL3piRGWYokCr08+i
CwARx1yFvvEAQCG3uOfmB4fW0qg6nqi9HctRWs7EQSMPAe8cbc+DsBe3PWjb6TrKpYPawhgUoRk0
EOHi3aO4nSeqyLDtKGOfwwPEoqslamUFmFc1JtvEYfrsrPD9n1Lf3mk5cPpTFrphsNrqaNl+bUWW
qEboH78o3qIoqtrmyezXfc7Xz+tr9lVNNm1+e06n8fDM9xn0KJvUrTedGQH3oM23ryT/Y0MUw63u
qRpl4mOgoCSJRgCCab/wOP7IgAFNdZ86wZwiUKwg95K65Dooc1pP354UxmTBcz5Ifu5TzaE3bY84
bt6JVYy5ZzIkx18b0Zhdq+dkTgQAbo41NcDQLub91ECBL8sYbjJlXI+0RFzBkWl2LqBAeQnvj2US
2d/idKcFKxoWnvl8lg4y3pGf3xXPOFWL9tUqpgFequ3I43eceA4LYG4HMhgYUcictuLmwNOUSPC+
iHD/EJ4OrV2YBXXoGyYECeFRFRDFxn+6/KzRUTzapXNVXb2z7JlAlqd6+Ca6j/MoySNF68YpQ6CC
9b5gkrQp0dRolo8xXoNcl5+azbxELDrNxc0R1qxCL9xb8Aal0UKvpeED6kmJbVas9CaBgMVOsSZr
oK1zAgoqaDR1MLoSLxa+N5mXhnr/mo+JR53VL4qspiK/F05UbJP7v5Tk1dvKetxvrN1Bo5xNU2fe
HRd3eZ++mGHHxpfOu5CTCnFTfrSUPUKIXZHHsOQV3Jtdj3d6dmIqUpa01qI+4wBFiSf1F7cT+8Ee
hHX7//uuwuLLS7McY0PQWi4OLFGfEHFZMRBNS/LU2sYbxaoErKhAxUH7SKbou1UBvbF7Ze3WGA2d
+mt1bb9OMtPkpWyswmxQNOktrJ1eBhbtXSHoANO3MkkLLhI3L3LtdDqqDg4D/I9XG49LgAqHBe4g
kKFciaIsy7yNckQZ3n9Kk+ZmMJPBWGhrMz0o/tl1g/MxFuX9OVTeGjztOI0/sWrWigojyM+8sVpx
8eRMXAJWQgg6TlD2zpnmjpYVIz4jBMLMcMCOdw/Fc7lmEk32yCBMa9+1z4nqT7+ntLcIY2/v1548
wtiBuC5WXMbFoGDaiWKPf10xHySpg7z0Ef35kC/gaJnPsIcQmzOesn9ll93Js4etA/QfUwmwyDW5
1frmta7FyTOx1EZlwuCPdaoR01bU5+TBqxAi9J03wyHG2ig+kQQtLFf61IH3+jRp6PNmGPQiHlka
eHogI8zxl6ukgyW2OBzdrwf8EsmCRNa4uRHW65A57QeJC5TQdq1adFr+31ny25lbH5IJqgFH9wjC
Ck0JPYtQQOAbeY4Ubn0zmTp8FXEf9uRW2DEEJt3ohi7vcU+SofYxtmzqrpgyCw+MuA7THcMUkSrh
N5/f/pRvJBMp6y9bC/ocw+q/HUleA2FEUWSPLT2uyOpzNaf30T/tdHLCEMCWThLAxRAHyt5Q5W6X
oBns0yrrY2t/kxntpgNMUhI/ydFUd8eDYAoRv7xLbYhW0O3kz9j9UD/lL9fY8pWpFITmhdtt9rUE
Ky+Noh2/qOWxhKICLHB2j9eFH+QT/9IxI1JJBEjGIP7bTtWRA3tKCZsqKGQROwC5sxCv+gQGHbKn
/+qM/F3l5truhSFydyw9UUbPBv9uworbDMrXxcrhvoyFM31iVcKCs3KPaeFatue92L2P5nzbIMNy
+80tiqqyteSuXWgL0JmnfYnpEENTKbsyidgnqTncqcqCUqGeAxHp0PTjhtCy804nl2CK1Wwynnbg
hcSgyL0OJBxC4GzmDxJ65/JI9tVwVljzjhONAQ1u0/ZnkrQ5UiS7qOw4hETSqWipwD9laRDRkwEZ
YOEIN6WC/BYOPYjXHlinmQzEunS7wFJEByaRCZYKr+y4YFSMcfGcfU4VmK2NV3PLGM+4qWcV4IrH
CKNvdyw2IFclwR1tNEWWIGlyIFgeBaI2xuKHwzTpFNvpUuJ4LlCgpWahmYb8tE+dS7qaYnMR/lRu
pVRz8B8Wbjh/fAnR6bK8CXGgrJ7Uy1Tw5LVGllOQB5EnZE9Oip5J3CBPF0RpLq9uHkRMfVhTBEhN
ItDwIGFlDlnK8h44HzmabQTmNgv1FiN/nMKKXvSstLFqyG/C6tmgsYEMkP43dpwXcy5YkV2gMDyu
B/JdH2j3gc0P/k34rld8RU7lwwqxrHqGf684uiPF5/egtN5Lmp5GKt/c7OC1a0QdhM9JnvYqsaKW
86SlUhjyeoDVXeEwUBDCHKgP5WtNybxu5zWUT5SskRnhwSc3WLh5J7Xb8zFq+yWmAhA3989k6gnj
M4G0GGsnvUnqmUb0rMBTu0Ckp6x+UhwIFsWQBJaDXBgTIoRzoWKgiut20810XQ31gCeYvjh56bBM
QxGTpvbgiZj7AnJqHoEJ6NifNT+fv2VMzA9CzmAU/py5PHNACixUotQdXYvx6fAkYu/+rTSRjsI8
ED5vT+66cReFUsMfkiQzA34tcVdnb/jux1JmNoAdxPton4cW1Sy0GO6qaaWtinxTsA+VlIvB146+
2fgPLhGT366JLrUsGZwlr6XN4b9xDas/dJJVbIyJOKgnTW/8Pqf3HB9YsrXyjcVHDtshIbVUwdxn
UBsd/w85aDLuI6gwXAPV+IiaTCzv/tIaPqnI+RoTIoe3YvK8aHkmb/wHLpbxsjs7s3f3QVMMaoP/
iAqdvVuh1Cy81naQQZLyNG6l+Rn2lqvqAFJrPTBhbo3xONuTn0c7bY2uDvEf8GCbcbPxfgsWL7XM
iYSULtXr4uFRwqgjq2OytydwfvavfYG9vASOcEf1IGSnysb+W72aPykt8Ll9M3b0yw1vd8Ih0noV
3gYLnfzEopeQVdShrTYBlKbo8VW9ZbAfJLi4OT4wcAHEe0/ataAu8bHvBhjjsQuNFg1VVHwpLAli
kIDw7xITDf/4njFbhHu33cgZiD4Wr3Es6buj2SQL2dJD0xckyVQLige/rBR+20fyeYQVJSQPNHz6
XBf/rWnUfwr6EFzud+71aUBG+BaAAlfbHZaIPySxFmvPvYCPUelymYo5vwc2+qS3VsMJX6+EeLYY
y+BnYr9MwuJO/V+oLF0a3Wx1YHxLCl9svpKFN+UfNxkQCoya1ZzNTo6ttk51QscR8O6HeRAKvher
oYCdzwxecoTsFx7RxH/kNu7FvDuJBX03vaham/CBbVFBjCRnraUcw4I8bilLzVWNH/V1QAdGrnpS
cNvcpCOfxMf/xCeGW3MiSn2mnh/AEFpp8Hm4F8iz/ZKSKGcEgXQdXMkmoc8KoOFwvNl2S4+BRRzB
pdEgeo/AzVr8UkIkUfknUmpIdSE6WC6VABwaSW+9FtzyX5N1EXV64Nf6C5XmGl36aUN6DQc4pOnf
Y9pDhBJX7+gGQ0L2jcndNS9y6JBQoE4eZZxcrOKfx6R+b1iCGDB/BQClevQE/yOeaK6kLI4wpywp
5YF2Ee8Aw2sOi5PsMmKo6dr2+UTFk7wCf4tAUMJjRJAbLE7GmODkpHw6Q1u2kukY7HyRf1d+bZpB
Qr40cAPNSS+tTFY6QE/Hz789+7kYBqQjKDS54bJFx172zM9uUaGfVw33WMOEB4cx+jq0CC6ty3ss
sz13dfSTouz4Ros2UaICbk9vvk8GqIMbCYTbZpcINMDz1oLbTvGoZ8loy6uo4ukH6SYaS1e4AlYV
/Ic9gLxrh+iS4Gx8+r0BuB+oYDk632Nno7Aa27+wktL+sa9EwKSdSNwR8e7UoFeUhbe1uciRvEIZ
FbyQ0O2bjS3py1TFLucJVq/Wb3nohMvvtXGK9cli+IZG64Q1q2YhN9uRPzaktLUjLh5IJD7KMv/f
CWlE1Bc0694Vdvy5g8ty6qlqUIHf8FoY6AKL6upcgyv2Sa6YqqLqY19yTVOELFJUM95VkrAJ/2W+
rn1hZnYynffAQD7kMN6mIwmWT9Q90ICTKbh774ilVwT+Oj9H+PI8EfT2j13YabkAx+aBYe796QNz
oDN8Nj2uBm53lK8sYiqghMj6pDiNI7+dbOidxFQiqTjZjP1v1UU/jA1VpqL619ogDLDBuKvu68Ew
ZfoALLAbYWjyS3Bq7pyqUiL+3YxPvZvMl/ESSOKCbjqiPuq9nCLWOBsH4vCGpe7YuavNf12PXZWx
ueyIh1Er5gn5jK1c0s/N2rPHIR5MP4EUxdPgdOpesHKyRjGKY/lCduUO4iAG11aJ9ASxZTqfffDy
PSn9psxj37imR+tvkZ9Oa7Ew0RP03BfltQZgpDqpKiKmD8lsJUj319ErMjDU1a8cV0GL2JLETXzR
7m37J27g1O6JVKyNns1hqFtd2dZtg36Z87aAOVnec1tMZKBc3SslvH5KALuFT1PyXKFElpqR73ma
4n8FPep6p3zNySoteDg6bqEK6cFf8Vo1Hz5ipkURM70ZpbOC/PuJUUGIekXjHyzKBoPWh3yE3r4C
3RegSUTDLhx3MlKgpoXdA4HMqbWVM7FRTKNgZm/rye9gg1nGKQzQSTImukQb0jTVaC/2lDDdlUat
LI/3XVOt9H8IqJze+Y7ovBeI8Rap+8vBykVWLjWjL8sqRI4Tm2sfUUMErF7Y868N+IiqTpH94zIj
D2TRP5wv4xWCK4XlV6rrmcaljTVO4eKKehdxA8USS5Bap27a678oZjF6mmHakBJweO9TSMU7Pb1J
ib2tq0+x1cNMB98ZYa2MXy03mnfn4gRiGwC8tb5XO2JusT7ql+RNdMY0qDeTlP+fwQJqndz+QVRv
YsD2R76a2vx99rV0BncsEZ1h6ATyMdUT1bAEI7Uzx/7TvsTl3sscpdH1H/rfC1EK5Vv5BLY+SHT3
Cc8B7a9EjRF9CKuHr8HRH5z1kjtaiOAKKudfPNLeJZeV2dCPLXTHU78z2NbZ/WWBoI7cPdeWBKLA
IfpN/Uu5x9Kq6fYPYw1hepzid1eYsealErfjLnJj7hFnipSnVXUh4+4UjgCNNG9dm6BYsbUMZyoP
SA0ukCmBy1f0easVsKiuW3Ldq9fdbap6+h4L/5KWkhwIXU6W1aGMSAyDuvX3LQ8QIVVwavrYn8cQ
uTsCXIy3c2ED3t2HogPuDyiEQ5chV7BvNzo4Xtpk7/M9UZ8Ns4HqZU9rKJrb9MA1HeUsPSDvgvzu
L5m1ObMw3/idIFfjqzr424ZfZ7ve4Eho3fZLYQZwGDYl/rT1zSNsoFugQpUFLsG/Waa75aBE5p7j
xO/z/PTjhDqeOK27qZDtatR/4//+Yv3mnNoaBTZ2uuvxEdFl0+0d7T9pXbnO0IPEWH2YZkR8yf5q
uTgVk92t7vDxu9lAQBG9NE85IG1N3gFbE728pjeG4lVmKeIYzMi4FQHGAuWF/oavFteuVf+YR3hG
4YM5HaYDkbFmI8xaRoRPReFqSZlqP6lwXKGNVaB9/ea6g8vnLYmnDHp7tobONTXMu9Hd0ZU6wiIC
FWUY31u9N8wtl6nE12xS6VmD+O5KOqnFWGe7At3673NYORaZ67lP0YqNZMOpeGWH9kiwxAq888z9
Z1IPiEYQ6xH7kPlrZyg9OitCA5hkKZefKRY045Jgugcvt8hoVtTQ7SM8Mz/rOGSE6gINtvsZOKbm
kuqZvDjfq/y2t/DPXRPt6FXuXBM9w5oHq4z79mAjUnk8osxywgg7Xmf3puhp/Z3lria2OWrrD5QN
zvgZeYHtgm/NYyeeSsCWZEizy1i19/t7hINR+b5zRR3vDGzKWYkTpf1TQqRmssqOcE2FuC3Wh895
vt0LJZEkOJcrfpC2zQ6Tw9wLx26ra4jJFnTDg9Bv5oq6k3aFqHpv+tyXDnGVJhPMFoC11wllztha
zjKlSGZMyGCUc1G0rR/ZpZMicA2VhGawzSi6pk+xXPJx0IPzBUiB94CGqHsyDzQcmTw9b6ug5uxE
O02brCOh6D4cYbsrh1zs65N+k8d0cgwF8d9RXTp7GDC6eFRQUalNHe/0l2LPrwnQXRdhmQfFWoBu
BpJUEB97V07A93mI5g5bG95sTgX6Ia036Uq+bvYj/QoeVKGDxEa+dooGeS2vyIC7v+vPI4g/352w
huDhWsFWCEmRFAkeT43PXBx2z5fc49npVrtq58sDGBP024O4oL63sJwwofNokJZm9+fk9GbvsG28
eE1l4CnTULRgajeN7t5v/EFE+XMpejF3n9tJ4xd+pHfhKfzTxkS2GbmsZdVAoxlyaoy1us/dxHHj
YQH2iIcoDTAkh0wswfBD83hnRN9akDDRZlS/AEDEUyaj6uPe5jL6+XZN+hCklfBLFH8TTq0/MUVA
zVNAxlO1OQST1QJY8im54qzcoF07mLJpN1BrYyjFHGPSAzn1x4ph2JRQh5jMXXSAao4Lk6R63elQ
33EGeKbxrrE+IIj5fARHER2K2C8Vml8QOmZHKrS9rH4ZSnfp+90H9jS+YBZ4IPyesdLoHuQZCRhC
7PYJ8SUzinsXqwtC2Ytac2QczYOi1+X4wjhuMvXWmS99X5NxMarYFeawZMeTYWr4c0bNQO0ZCW7x
hacpXjReDXTWMYLP2uZhiqFRg8ZiDeeAiU2M/wxzNiEw5xe5xg3KGiA1wslVprlT/rl4InaLgxI0
2pE086hgeu6YDBlIOAIbm1yAxY5k7nI81DPSP0v8uNH4AMyxN9nUydPvIe+9tc1DWGQmhXRGdHsd
AT+F0kgdqQHmbzg6ob4+05A+eH7bRlpwqLPBPS9ix6ZfG2hKJ+3GkjuNw9LW4uPEOrxH9T+ThqEm
VxqACpwBwNi5RokQANqQY/JyNo4uJhBuVIlTNBxI144zAY14alKMpaXFSVywNEBdRjR84R2fbfBk
4k4oguygqj47JFGPv97KBDrToqYvC88D/he08Wfj92cma6vafADIsFzF32kKAO+gTWcsmlVUL0vE
6pD1qaN+rnXM0LBg1cuGhmdrIckMP9JfrI481R3eTSB3f9M5sgmfdzOlRpp0gwQ1GpnQw4vaOjNj
rFKhEyssptMm/JcnPIA7VYAcUwGegq430Ub5PU8TSayaKNSVRzOEkOA9okNccArI5GS1zFkU9qNe
2k5LrFEpXa35YkgcFweIrtWZHb9O/nFuwL5AOX5xkG7EL4znCXTAqOsv34lqQ3Te3yfEinvaoFjY
Wy3J3k7LWNY5WqiCJZZYT4VgSKH1LcykHeIWsmYsgjY8y9ahqgyAxjUP93Uwbg5g5g1NwIydk9bq
nS3ByFueVPr+UGZvGksW8h23rPwWF5/Ezgwx8h/ibGN8bcBKAZhkOVEshUbx8l6SdddeRSNGWjK0
o0Xgm5DXjtr+apFRey6oG3OXgdstC65jmQFyRFoMhf9p4yOOi/VtrurBmXl22PjQp5pngOxjh/DH
Ivvr58hoO+NFzGweD5smmX35+Oxn9+5/PZAPIpNuCA4g/Z4NvgbeMN+iaKc+Pte8k5RGUu2sjTIU
sZemq0C7HYBrgOu6HxUQQvSfqsXfLUT6wrPFZ3xHkP+iE/gCLrS/TBMk44hbf6aQl92azL75htBy
99TiwvogpgNdp3zrQrTpeVhYHyQ+h64FOwnPdrJR6w+xpzcaZnHjlulJmcifOoj4MQp23wwoghvL
GXkDt+dG4gQ4ofhf/tk78BvTTx6Y82tbWaLeNzFwGfBHiL5OaOE0/gXsSokAMIQ1vKYvCM/bBZkd
5PjEAPmmpSNNLhjo7H3C9FTb4jnmjkf3zijVLXjhrTr0EBjJ5yJpbnzh3BlGJ+tly2gi+91XnZ+x
H3nRzHzgxiuGk+CXfuoQoq3NhWOeolhUswXTQUZGemq5dQ0nmUhCVj2slcR+nHRGGsHPd569pHH4
t+44IBAb+xVC/9KBMdMkYCa1FqOyBNRyxmttNfGqA8ZPT9uLjlRpEf50wSZ9IbG/r2JaZha8p91T
caA3rfOcRA2k6h33+UoyA9gsG8ZHsLq6QPkUuOKQx6U9rYMO8ReUviHvMugyu6Y61omPY29F4xga
dIaq211TeJTgvOkRJhDH/DnuqDOCqPBVcIa63fprHxdg3xr8Zn/zZO5aF1CmXVtie/6aS+UsdWDw
mTFnV7J9k3pO308x30FlMpV4RXttbqU8LecJuZJY1ozw8e6hF1CW4x+uB6OFfnwXpXqmO1M5r4AM
Mp94wVB3FdgNcaBV50i4/MeIVV5TXmt3RCV+So3Z3/B2dXtC29ZNImudFsp0N7f+FRGKH/tEASPO
X0Zt2jNwcr9ejDgddz7uqWBqyMzY//dK29MFeV4TI8xUgPzCqL7vhQL2NzAAfCDYcwvE8geq0TFd
pqC88AhwIl+FqZhm5JghMcEfxtTOSfb+0WGPC8hBAwgM2y0FoLKi5dA24dZEB8aUUvsehAnMxQWc
iH49fHqBRelOd1tJyB1cfM9ogpf6Bya0bjagG4tbaGkNlcDx3GKwOS/abaY7cok83oiIJ/HigGRB
U5QYNxwHdDC/Awf/TFGr2NZ+1Kcbh9vwuRhi/Qm4zAUlEF1BnlU2kKQNZAxpqI2yheTYnxOrbBDB
06d/epjrWwaL0UrBCaRzzOhmnj2QDbNG7N84XskO3tACFJvLFENaZMEPTohg5XaAYLumQ5wSGtBd
xDhTVNhrutKsRTGq1+8APyNuhGDZFEEbBA91HP4Y/RsFYhQtKCT4kUICXSb2MwL1kJEq/kCo1q4C
vl+CBjQrOSo9lYb+BfKBDrP7eT0E1K8xcxEP2vYXhz4iAZL5B3/CS3ARv/qEQpGmMJImwny3Aynh
03CslGh7g3f+UZmzzVvFr7L229wW6yuFQpd6ndW/mag0OWx8/iFcLdj9Z2oqzije74xbXgc1fVkD
JZO5+cDOnAA5/Gk3xOUFU/Pcmcy7gbuqrbTrYmmggw18Jw1Rh+iPi/2O50uZtrzbluXiYMY8HEM0
uVhMxEYOu+FojBe8QfGsC91CFj/+5isG6c40HZiJ1jZbUtkSFpGkcX9chFHeDDQBzOhrNznrtOqj
jQXqcUu+S81z3hfXXrJNE6bVxYxWvgST6Z9lRyH/HnCeYFJdP6AVlgmRGwTy06C4fuzMIM6nsBQH
bxXVOcwShHPWpm+9ITBRO4ZQYxSA2KK4GYZ5qxjJeyL6h+s4Kf8vK7kCaSdr9jNcnX6xMXPB1Jaw
/b0jn6Jjj6Ap3vQ2N+qj2EhebaUp9jedEX8m63aBzuxd7lzYHfJ+pDbIlpXBMK6gAQxS5SfzI2Xt
YS/sKKwIGL8OEKyrdQ7yFFnVhR3NZe6gvNWA4n6sIFsmZOov12tkJ/3cJckoiN1rQq0QkT8yRDkh
SCFgtL62EkXPISLWHb0WCQp3u0U8iP4mXak++B+aLpkI4jb2RJIajnjaPy+ZF/JmrvjMUomUtXuq
j5gfHd7OjVtINDjxE+SO7oy79/CBJn639/m6+LgvI4vxI0ZwvjBf+ZvEAOh6uFokmMyRmAJBJ5Fc
o/JP0VP4v4qGajms2WyiYaIswvIeq+qy2chi4xnr7OschaD5xFKnGK/7faThSuTkPfEXT3gWYaE7
n1hfvLXOhSmzjXqtA3knvhQgaHD9sDQ2VNxXN7pCYwWYO7lJIksh/udvKAJ4TWfe/jrp49HGBomG
Q/LBP1BsS1QATs8y55MmI3fHhj/bi/oNj0BRO2lnk2UvuJgmjcCKISmqq+oyyqSpkQ4uaWeyD4rm
EnCM+ZmeDphKQiqTJ5RhiHEykjP+xhqZcx7ZWK7lyyxoIMZzwnY/5c1q4iRIiwWzFKMZIyTijuBU
URw20A/mCR7iew0QR0gxIefQCkfQlipJY0HXrgvto0XhBUWh4YWaN4a0eM9qTKZEUuu7qybAMaIm
uXDeCMXdA7SHoZhjROkm0rqA245XETI6Yj64hwni2MIbQu996GUD8CGWAdRpkBmPtoSaF7Bqq1pF
GbDdPbySrb42sr2qrVZ1mYIZlsbYjfUMwPw+J5wZx3cp69GWkzC2NgC57Scn/AvE0jiZ75ntAAx6
voSMI2jkw6Z2gg52q7TU+3eyUulvwtk7AHbzcQTbi3RVsOJQkid1DgkErwMsO23LIs8PAPnHAPha
ovj3MQgPdk42+FBpqaWqA8hMVqtcq1Z5wS4ZQt/PPp+fyt4/CEZ6u2ukyKdRcnAhHX+d/3+mUOA4
JHEAWNbg0njonp9MGKV9bis1G/jNgdg4QHhmhzWcHVqNnMLAoVZ5zuyENJkYahiptiyOv1eFYpo6
iUPOpwWy8fxzqCJ/mzRc659G08v/hAft6N+ne1qPxodE2RBZkd2ISUvOO+Ex5wGSNFx6rI+aIrR9
qXYYhug/zaRXrpj+6ARKVzpr7NbiUh+76ZVxhBnq3oP+0QhR8I+RCudzs/QJzt3waEKglqCrfqh4
StBDeifMa7uYwArW9bZ9MgnOP3LW4mKw6BwoD9NE9zK+/OAzRpnVkYD0IVOsXzvx6PsUadkYARrj
Epfqcm7K4Qe6vPQM68cosGrPeQB8E1QLK4vXo/ktLJvX0gZbeSp/JrPkBz1bnayj4OxvrcdK4ieU
HW+u4eVA4loZACVsA3QvqvCXKPzpnR1/tDDl2FgaZmfxfYSUArtKSVxej5koHNsilcQ7a4LYrcq5
0QcduywV4uKwpiaT69zu9OXKcLW7qKD9tBnZXTqmJ6aO3xNxSRAMcSIpUiUtRzImIgHVJUAZufQT
YDtLZ5icWy+JMDNlq79SbSzQXvl8z8RmjYpVEiCkglXl1GpCsts2soWlOBjS7V00JsMqBbukTojc
AdIoWrEx/NAzVFM2CKEi5IYFpiPOekR2zWKqtqte7qv9z6BMGJE1bCHLe0EVYF9aJNl40fuUC1zM
WCEhuj6pK8fwCPSa/X9tpbYV8d3pZDu5Yjd+031LqkcBxwBA7Q0BkEeQCh+d1cXJIcYBbuqvptdu
5nlL9hJMlBPfesy3ZizSvL4ZJToB2VfJKwHFrTMkKnhmqJLYZMsxP5N5AgRLyiY+1j79QKEJTES4
iQDr1TJtakFa3lnX5xnNsoB0Jro9v2xAtXhfUWjf21KUt54wfSm/eaVwOGnnSfq7QnMkVbzd5KeX
0p2i6mHZIKkgwbehVsRhlZXRoB1pmWdBq4O9bgFXs0GF6sVK2QE/KMUV3lcolUP33yWTS9MYkUUZ
+OToqRq/t2itAiDJLzBS4yawz7czZ2dwy8O/HGMnSYOPD3VbzZ7cXxFKMaQJEWa8qv2jgg+zLe9u
VvUd+5LYAkx49iqkwrTyARcxMuw8vAdQiNVMfGMHYi2xOUV4gVPXxxHozVC8ulgusz5NcKGQCQ0X
S76grNHGNBVT5Hm5zad0IQXmjWcSOIU6qqmX7pDqaqzKXSyXJY9kD9fayIEpfrkcXUsClcBLj0wJ
k4uVnLW24skOhpXEMDRjTCrSfzoIjd+5TnF6hQ52uLrHcMU1JbhJFN5Whj/tx4cN415Pg6WsO2hB
IITA++NvcBI8gYpP6chOprfYzZeQrw3vR+L4kd1mnvK4igjtF6c9qHkKxLRFIdlRLbNPtA2s7DV+
hEl6BsjTyIYwZK176ebhTPCaVE8DvBXtTHMRqHOS7BeSJAXoZSpc2UYCMaFFgv+B9ALE4vXbEV/B
hUm+bp7T0tW6hB7HtgimvCyg6QFG8aT1y3qm+x2giejISUZ9Ztq2SfDbYe/qzozBlrjecJgT09Kd
5UdwyNXHw7Yg+t6LnDUIgBlcRLGxT4CP0FdeMMNMY/ZrLk1ik0fKSd0StNQZYWOU5gvqaQ+nkB58
e8UGBS6l6faVo28yP3rhduVnRg0onk1QsB15/ImbPfk71TN69jY6UKsEQnMpXMv38vevq4Y87xwv
AT8ErJSo74hpLfJqAUh/wnC8pbd9HOUuJoyogUa/EOWb7TF2THrCkMgN3xRpvrAwqjEsKxH66HiG
23+K5gTFGfKN9aSNKQUmpy/xe/ybPpNslFLXKhHh58dHLLmF0pAN+quPIcFCpRmdiW8hM8ds9y54
+lP3MwczeQGkIHvipWUObhvJlB+8XekWIYE23uYXNHpIZa6q7jFDncVtL1L3EyAzJoQqK+nuixhM
nWxCJzTeAn1zNKyjA/LontIZEI0Q5U7fZCBTqxQqLFbCxKnxlCWn1gCkXGYhsDrADCACwvWrOESg
Cj5pUf+U3XF/P8NPVqMiAlahUbQe8X+5VKCN/+p2bbI5NpYEfZVrRsi4hlefZNq380pg8yP0xkJY
YlXkob4haVlr5uc9CCFemvs2v5+7h0J6YZXOCukjjyt2J8MyBoY6iN4mTcfjMC1qcCguzM5Ij08j
TxV+ASg/o/+nhAAqD/wurxb4AB9r/33/D3IoOcDPPhYggKgutNwoX+jUVQgW01BLdxYJ1zEMU+8i
pUnOSRp1zwm7SAlc2/ShMjPVl3E0kWn3YeLVG+7cL4q6U1Wbqz26kmLQZQaz0uZ+NB34TJUG1zE4
HjkKEtguxpmErz70XdwNtRDXmrbpM7IWs6+fRQCCragfytduSfrMINeMlCS2BNboDoomfemiVoSw
ZTgm6/gbH0P8XFuLpR79CzgRb3GNtuoUpegoRt+NUbLTE/aiPp2bw460rUewL6RSd6q57OJrxgHV
1d+Wu0plHzNV9UhpkwWam6HoP8NvWvKlxHcUw1VZTmjsvQGV4hht69djbvFN1+Xtt5rIMtYo6DIu
gcm/Y4YarFUw0PZL+XWZdEIFJa2dWcSqcmylGTodxzgVMdyHNLKDeO3ChH0iViqJAhCRKJnfbnjp
fW4fXFB0aRkbsg3NDq/Sl0O66bBPTXEXwejLxCYsfDuJiZe65hE2desrPyioZjsr9n77/svERQp+
NCPV2zNnJsVtUZvxXWSdn8rAd7YqxWV0lvdVwKz27+YrnUWDnyoNw64EeSxND33pFWW3FRQvHtk/
3llSkT8AD/43cYvViyI4dMLBIVtW4h1+0yKR9Fko2d46rS2icrJdTjonTTlWcnlFQjealqMDiN28
o8XgvJeum5OBfZ4OI9HOP3rp1oQacwMtsA87DRS0kurup89pIBRJ03lyaz+ZJeLu0c2byPUyR9F2
gAR0Y0lz9StZK+YNkJI2u6/YonvnGmJnufOqQ84397SPP3e6JNDpRzrYprHICzSYxhnjNTU9kiOj
As1HHlB/cF/DIYRzQTmjU0A5AwTY3tnIs7R7UajiYZrEyicM1lWXyPaKSSmSATZkgaQ/95qOwO68
4LwsVIxlsBGOLp78apaqmcXZj357LX1kYjIH+ge4G3dN4cJnjOTR98yI+G/G8qqgLySQ4HgM+NE2
xxwBk0oRRhD3yYo18YMy+CP9X/VaFAL9GGnICBxS5uWa8+Zy/4y1NQ5EaeC2XnqY2BBBbsbKAnvc
56X8Ppe7mhbRA3gzgDEkxNFg0R9+xxAuEpxlDaONweEaAW25Jolq8xyJV1k0xvE0UIRa2qWY6wKv
LLGFDwjG2jMPLY65GGdjw67vD50d224MVqEC4ZhDGv0PpudWP+MXKEIEpou+bF1kTcsZuOCLiXEF
FXtKnVF29dUIQ4GZ3gijCDychuwBNEw+KMyXhYeODcoVwFmNylnPT8oHg9A83H/Ab8Otz/Iav40/
ttpbAd9AxYiLpyolrdh11nbA1nJQl9oIgQP7u270Zcph6itP6IANZjcD4D8kAY5uF8VX55V2STMz
CIQoDv9vr4su5mXDENkHBdYF38p97Nl4+bPCsJGWX3HFPweJUI3ky8b8LnQeikbTnqZm7c9QUZdV
kB+kSaTOCu+HKjBgnA74DfDRWVIM5+V96L7mZ/1kzxhD35qPEmtL2EL85LNzuj0Fuh7xRDtplJFT
J4HHgOzuAPfWjTf2jJnUPrewWWZtQsrey8r4pwRJNEqfuq0xjZRj/YhgbXv3fccQhSc8TvgV5EIY
XQaUgppSlyHXur9ypclVZCIZ0VerZSV8ikPLKiGKAcRvnKcLAxBn60DTLS6s6ffFq6GGPZZUJIQR
yohi7MEObI3VxmC+9T+wD50NAspyHWM6UjzPVZt3Tbbbmr4pFDNL4l5UEF1hnTZ+v4U2G6fAA3e3
AHRokUaOJ3wNAkrNRg/LbgoF/0xy3NMeoJe9McMbnj0WyURxy2aHDjOk4R5KoREDQg2LHLIQKDhn
HKhJzuII8XbNVPI2SOu9Ow/NBxcwf4Q3y9O/OxO8qYQFZG70EPGa5jgppGSxlg9DVl7+iElRPDwJ
7b3T0SLzyRcJQAg9I76GoaGUL3lvDVoqCG6goNj5GUF2trKDMBJ/d69cYUhF2dvEq9R984oZRdQY
XUqW7SBSNY0khC6CXgNdAgfFjo/Nb1vfQZeafC4YyrDCnAIl4ahxC/kqTUTpjaF333ywLVMFdL87
AQquUeEBelb4pVhe6wrs9f5WogkiTOfVVJFMUJM875e7MCdafpRy4bgnyy29Q6Pv56xOcLjjuAo9
AZEf8OcM4TgehrBhBm5LliDlMv2xoS2TPYiBKWlg2DDFxuOUsDjYzG7GQHZIFU9pbKAPzyOTSktY
oqtAs5CYtjA4OOILyy8nIzKS+EGF2NsNcr15XwOUPcxRoMC/eyiC41cSu2nOHVm3sU57AmTBxCbd
IE+ev8WFTAgruYGiCav7yq474rgOEqI8AD9edVJsWCrrrY4ROQ/Neky77kRSlu5NegcOHo1w7Pci
t7sS5xFrXmpIxU96GAjUdxfTY7pew/SEq2C6AMyeK+nmGqYg0Y41vk+Ya2ysPqKyhYMA0McCfS7D
lcd+1c4f5CVsHPy1LzO2YAMkwcQfpKYBDJaPQ2BsPFldw09noeGlIGRrtjTBmut2MhyXvQpsxvZ0
lmvQtNZHHKYL0wMt92lXR45x8IwVcfw1qUUpm/IFJkY/HCR7Vc9qLkZq1917mrm3vSsha6jJ8xXG
+JBeEaKo0TAxNM1IcuYIqEJsHkQzsv2M/atLIzSVJHZrR3aWuZ5wQOjHq67I8OU/rul1O+eAeE3v
sC+7QyDHT5vSVhYvh6W2Z9P0MOuXlCV1i+vGCb0Oo6hwM9h8r5Q3s0P95ierwI/Fl57bYTQXERxk
+frSCaJ8P2tuR33miL1VS3xic9e5FnZEpV1wWy9NCUCVjDtjX+YKZc1T11gnVPuOr9TZtPCQZCU7
xEuQrS8eLMZGpyusWGeOn+hWyo++MKWgl0eVjfwkoZ5dbw1+Uo9r60w53CCyfOuioj9Y1wkZuI0e
Bzjifnd+Ebt9si2dD62Jpy0QVfEpAOsDuAb8qjb2k0h1FyhX45h0236Q2Oaw+PI6uLGDiFen/U+1
/yv3geirGG+Mkyg+xOZpAtMacoSjlrUJs5v7bYfrvWosRLLo8uu9KmLLNA5sE7Oh8eklibEkWZRX
XZb24IzraY5k6Uiaof8wFOzhs9cCAkjbATPZ0kNHR4iDHohDNb+PHOUhz3e6elPzlyPAZVehqif+
kyqwmNAXRdd7+MPLLyKwFVU8xuuougqtQztjkt02AFmj6hfhVGBhMyna0Vw7fBiy6LYfmZHMI1KX
E9exp3+sLAiC6BCoPtZSfoZbPTEfa7QtQxuHVBOLPIfqApRsJloXLX6Tjv3jfu4J/ydw8XxVcG4C
gV0K5mBjOnzPEuFihK1tmw4shG8IoXyhi8uCx29ozAPay6otBa9lwzZeaP9ISM8tMph2sOT29o5c
dXEiMMFuJl0jZJa+gfHpKCuoeBG0EqvvYr574AxXpE4WLVa4M5F0v7vmaBg10NCQb9BKm1nJ0zdc
RGq3+WbtLwlHbgaoZimMWrKfrMaYQaR+ZEKcF/FRv45f9/V8BmoCfJo96pZ2v+nK/RumRRHrGGPJ
4aBIJXcgKeAm89iNDo/N+fws7qOwClIH5bwrCnXnmeepomSirRv8tKLX9N/AB+BqiNhXzGhmzbAv
OOktbFgzUfvdQahtt7NGh8NGXZW7hWd+bf9GEuPFopMYBK1g54DH0XnZp7uyuxxuWTYmUZIyDdko
YY6lRRGz53+xOPGVBWA6EtYJ96Ldo2ytqNzkRwU3UV3uP7PX6dxrgsNhREV3zV11cUOP+K8iH00t
4LF4J/YnA3e8MOC/tJvIWGAokbwSohWXT7Po3HaeHt8QHwa1Ua9sQ7IT/9js7OdfBsunF2ROeBxA
DLaGmve1xBwY44sAPjztiOpCmoe0s1AzOsfmyX8ZCP2oQfb5fO3cYOq3/4lAUur5nhiKMhriJTmP
Do7nOlHeNyDcDV56IGWdvmoXlnAFUEGIwkRuHXxzELX0Bkz8sEuHnROsIdHtbCmBCW7PoR/RcZxT
wtYrlRbApXptAlp+iDIIG1qseY8bT31DXWpvAYxFQthGK/mMFSHY8JHLr+TKVp1HQzpwLNyz3TPy
wfgC2v7is/5spzO9EbiYxn4WHkStwbxyIrGN9dncjWzADKmTrk+SFsswIFwD9QXudRjWP+8tolH1
yqzHj7AKOcBIH2Wf0qAJfaIwLO2ZhFAHia9WN/+T+Mm6AG88rHYrjnYSpXryZDrXEUfS2rh29MzJ
qUu79sJgMFkODt0M5hNv01MB/n/3W5u7GScJgePeKGz3ZnsWIKC9xcU0Gj6r+ihS/7kt/uhKKHe/
dsuJPo/14od6zmwXM8tI/cGy5BDvVrmSQX23pqp7150V0AdX5gojRN9TRAhCybekmPnqT/++/akj
p33mL3XVtWz7C3w+sEgSUZQC0MREvy84l9EHH2VEf0gmhNaTqReUZi5gyd8wR5DIDOdC6UUVoXWD
ZUJkVk3Mnc01NJt8gI21Gp31B/1LDpeJoeNzrfKSE7Eq+a4H1HEhlMZoVFjubkM7IpPxHjdLiVOT
jigD9550aTvPiRbKIRdj4d19iPWGM3ck0eTutiD9eLaWhk7bbUGyzVMEIt5TawFKIWZMPTewFlq6
CmMKAURXh0raHm8G6SuTyB42xIy2j5hAHuEbfR+ZNGWbG6iRbJLve9q3uQ+bUm2vwJo/pmdwGxb/
xhqvh+kmQ2nm2yz6hz/qnbQi1ZSfuSimg05lRUsnDfXrepEr9353CU8w9qVozTSbWZhZI5ksy1kY
F8dHHuvStvOhdUbkAHWBKpqffkaQFYEzL4pM4VoK0hjgIC6HmFFIIP1T15MBWP2swE22Pap/KdFE
5c3VQ6JO3jYCIdhXrP7qqUM2/gM5CKPkZWHJblgb1BKzJKzqxU6dDyrgbISlnhk8BQO24pw3HVYk
WqtNoAfz16nd5B2O7wfHDwkpqIxlt0r7xLIyFBRAoC6nA+6zdj/gyQC66XT+YYKCmi1kvnyZIeP0
kM1q/lVVhpHVQrxHf+noXzXrG0lyCFnS2FqjPCbrLt2PFLBv0uGPESeKP+Wql1YxPRGggrI6xCmS
KKqDR3Pv0FoeXM906Gc/AypJlGwJc1lnMIZY/uWdnrLSp3JDLwfgDq96MtCz/foRWxeATQb2hnfw
eAMxSsY2rExzxsgt0HrZ+pkayF+OqMxczmCeeLvTOPFv4SMvtxtqe/lTkxln8vco/Lr8dv7ywn57
3JMAKUgoEXG/HuyFaWMn/u7gBC9pA3EcBJ8RCgFGj5J496wbxP75Jtuyu0Lm0RQY+nfz+65VVDzB
lWDLM0ocVjoUvqqjcl1hyueJp7j29oBUMJlwZQNcymN261bYKfM22JruQ8JNFJIF8AL3vDNvePJ8
WhULyNDLqk/+8Ri/wbB8/irdFotCA9BaUEoqUc39G7RCu9mt/b34Yf210oltPKU3UwFJNiYvnGv6
dlA3pXO2CEMkx3471khPzxrKehacJjj6Q8L0JmvUL6d+iexYniSSUV2OF5CSHs71Ybux/qMB/+3s
ifmdH3IBXUci/CnAortbmnkN3/+mDq7s3euUbWRke4CKsAFucZKzx+08HjTKnS5D37VNCO1RPsfE
3/jXqOeGEvYZZ+sVOmUxGr4WF5NhIp0CGjSEqIeI77NS1e2vHjKE5PBFKq1ja7nko42+MyMfuQpW
AwFlRAhU4Mc8c5Dobxh9kUPhRQGy944uTcFDo8k+giRNRFWA5RZcHalYGSyVh7Yyv3cRzzCl93BK
ebcCAPDPwoK8xmQItjvktrAi4RLY6VD8FmliAWbwWqEp67BZwK1+03WIvXv1/LKTd6gPg1VtilyL
AIbTRiX0MP2MRK9krLGYAC/ff8g8mvILCOMypcOywr2tgwK6K75slmsxrgUXXvBn7lPbcw/0k8UX
+rDZD9AlRCQagI+6cTqWAJslglUNv/tO0TU9jsE/Iv59Eza4OdH5AR5naIAtymZmKso6+kpotxYg
CrR9SLJVXKX1wClZEZRPG1XlUSY/txblJvyfdotjvDNxtLXmpbwAm0dMIR/hL3qQBZ21g0fQ6lVR
V3mDQuPawEy9OCnN7oF/j+cOud7Cv13dz6+DmH1e4gZqbtNs/D18ddjXsVusu/wS1vHZIk45tyDA
u84wTJsTSvjKgTCXRnFsJzBoxW94h8Xut5lJQtLXz5WWnHWyUmB3It7TT/vWuclwB7GBytLUG5aX
2cTVEx8U0/9SXrhtYYGZkl2+T8ldSvkqvGrmN6QmMYh+1/paZq/vyo6Xl4XBZZ2jSNJqqQDNnitd
8uwwU++lIgwAkGz21dQfQXeDvZtuE96ZHDQ8a1ai817+n2Yg2fZj427A+Ab2fEfnh47W9804klLF
4lLVRo0tdNaKVTVsGbj5rFpoMI+AzJ1cxv3Ra2/Fpi7zJhDISA6ky4yhgvQYZ8oOACKQFqLmI0Ui
CXOuuzh4wjL8xgBMMsK1kvFd1uueYsOpJocebHQ50hpvVdKEeTYdUVVSpEQffNX/HfVwC7lX610D
zZ0vs+/IswDQQvzXSEnRlVfzD3hduY/ozB1xh94vbKbRv3/JtMouK33qoyHPM+0W5YqkgITa6Uy1
Har27JV7FATMbff9dh+750RLL/GFsAvAOdxi+ns9PDO2o10huvCCRKkK1HoWkYLj8oc30Cy93lkk
Ln0bZLkiHVnDvwTlQio/zWtBB59klpOJMIxmwP6tqNIn2B+QisYJNZKE5bfiO12pn59tuIaGSCjt
2IkYOXPvBJe7LXGiwYlhhUstp+iAzIaj81v03RCPkOcDpEAAoAnRB18AuavAaLLlQW7KbkqoJSiv
Ji4g0OP9VZPPnhf7oyi4K9pGrXQ57nYeerMMcbtwdEPQxlDs+XMlvJ5i76PSeVSMarHQSDqA/CKk
PBLksneEcih8PyI1NvlWjixU7f1CgNTVEMud2lGPTcjsDg/DJQQh7NSWcoygV78zPnrr/EYeohZs
S03eAMQTt/4uJoEXZ39V1CUermcD0atkjpC8xBnSIFEITUZ3cT0jakEzrOHYM8duMoLZNiLM5Ezz
gdT+Y5rpPG5jZfFnnXpvPV26emlLqCJSfzNO/b++b7tmnkWOKyd+rTWPugAvspHCoteqYTk/adtW
3kJfDVob5QXXWRoSlhA/I+8fRIJa13cexTZxtRB71rdpFVtdm/ajCpV0gRdb9vc6jdROjd9GTRqH
c85Rd8NorruIVMmq7+szMLdCKyGrvM/M6rAmR/voXGMhWnNFBK6sHeEibztv2GE8NkFfeY5GWdV3
ujxBHUvYvUESgqb9nC6hT0NpM+Ph1FA/++clT/zsk0/uFjQVMeAScG27O/cbIj7+Mt3aL1HSCgIP
Jm7H9LuaUDUrO63+KiL8aj1X/BFyCG1n18aelpATtV9Q9VSDzLxiiz+QvBEPRkq7IBmSY2q9hRj2
nbPbxkM6pWVtKjoHvD04W61xW6JLdvy/zq94cpbdGWFpC9Cmgna3YbFllWtc56k9J5DpT39vHTdm
nmH4GpE6vK84oJGvExXQiiR5FS23tpsx//hqVdhXa7zoM7p0rd0jxRza5egpsyXMhugq2GQhK2jP
4jRaLnGt1fThUVExbit7+GNDdIFWyJt6JvBJizpNi2dNCO60v1OOGiXPGT4CuXLpZRaipoyFyk/I
bQ3BS0sTQdtaSZc9mwIGfSB6QC7/rcBxZDAYgpP5gQEXC/sp2pBY42vlxn0zxuSVOk6lZ2BxTrq8
fTjic5fQDXAcBHCIaaAfvuVGkI+7/U9+lBt5VRuzICl4vELXdl/VtHflB1FD4oB4BonLuUGVa414
nDplLkAiIXm0T+EeWRmjPTvSrDyCvwl265XpmWmKAdKCBsrBKE4Yvm7lhiHNWcXl4Hze4R9Xlcc2
wZ4QbMLUSYhzzdPUJF9n40+69Q1GXtpiIdIhejc8CgE2RSp2lR5IUNbQ6Zb5cgmRhjnjt1zsVmNM
q5VorFkw9nx2V1WK4YE5T667tr2HhJ54/rQml2cfy53HHEVTKcIl5VvrAZsYLv8sjL6kGLDm4+Yc
kuDBuY9C0Zk44fjliYqEn4IjOAxy9INlBHAsgVT+KLq7WmsQHtHufEzmum568m0IKKYhwtrxQxSL
OzJK78fVb0xmL/suhLJlB1V8URV/2wVhCicPyThvX1RCqODHheL1oFoYnv7CQZQckSLVfA1skQYL
RoPAGDLRXjXUxVAgTG/YMjCZVwHprn8nNCv7V8jrAA0wBwRLkihSCzaj9qSvXSzPflKYFy4ve0uZ
m478xJ0lyZWuUZniRg6HdPF1Nwj3pAkVDGYwoLMz7cVoSRRfOy1Sz8ywt5YKJt1NRgcCA0kgyHY1
swtZlohIytN8ehesyYLvdhQhJoghwUw/Q+iP2NSQz9fqiKLrKBmAzDI6P6BgqMI8JnfmegXXY/9d
9OdU5vl5pH8sIwxj4OXP1WphUx07TkL9bWwJuJwhVPcsmsGWP6j1gi6j+tZP7GA6EyMyAG2f6CO9
yM4HZDc9gDftKCaQp2jodGYhIa/cwSie4u6ROcddIN/8Gqq7+yhNE3PsmXjChNm8nwGt3QUg6Xnj
eURHjVDVSoXmsQVvAkqG35XfJz/xQQ7ldTXLKWuy7/Li1TLs0xkZjYEOXwwJ0Hn4nk+GQEDtHS1m
rWYoSePjbjvGpPigw6cZWKKIM+dVrHayNGDgaI4vEuJjlB1JzerHSGsb+ZtkeolsZRqu68ipiyb3
OIc58SWXtVntU5aKDft8oB5M4/zusLvrCZkAICW5pJ4Jd5IXpXvXzw1bqMeLvyyLoZ6Z5nycdS5i
bIanXOjfun7wC07lhmWJPRai2K8QNc0qg+l+KjCwxY8jhTnwWvp8HMIYAkdRBEE5RV47okmJ15f5
S0YaGumztxUV5fLPvTE21vF7apiosbjFIABywsAuXjhrtrYQDs7p7af8qBMc0iq0eOhpcZY2nCew
JJrR5uVh8mieuaQcK/CYI6F9BFAVi689TG9npwcFnYzJl12fip6b/FdY9RAb5wTONoy6477ZERal
EinrS6WOLsHm+Rw6FTwGrzTevglz8jMb30b0ZZBvsqe9t2/0kcbrg6i94CzfG3CsUiiHdYpbupEk
mFD0Yjacmcjx58urZXyvn9/xCxBuxOCp70wjgxdoghQTr8PBdIzADOaa1kOIwwGTW94GffuR6DA9
cUL5/E37C2D0TocS9Ob1U/1lLD7QpYST6pavOWaidiw/0I5YHpyRXT7K/0QOuwiNWe9nnQQTEmuJ
lDknszb6w7XRIMPPf5aBuz7ldnbV40yPAHJIkeYqSaLlKTAHoHCBC+BXzGk/JjvLpsJgISRJcKXb
knG6Kz+FLLUz6nYy2l//HkLlrGgleSGjDeCQ6QNpuRXKGSL3PZBtwL0AJvx28BNZ0TK7T1Qts3RU
3yTqg/9Rhb2YWDoMppBcbyOB1LK2FSidxX2E/yulzbU0tqxcBQqpekcaMD5zu1JDS/7b12F5EWqH
YtrTRniE93j/OJFjuhiQjWU8ZHJa5ox7sUF00lWSzsvkIpkg8y1Ik7oz/hQxmqSXlzcqw9eVwfXD
k7Lq9YsxygRbUrziexhSR6hsnSNF8fJCZvckkUnsKwaO19P9ZfQmMfNxbKBP9rRHJ72/KCTTPxUW
iOUCOMC9WCZ+8CvwGoNOHYEqpNDD/UE8ysdt8ohU1Rpe77Dp/9/5bODPorF8L9yzFU8lFtcb0rvX
fJ8y4PUYiKkb9kAWlY69nG8c/8F7MQ26xNJuFiqm8i3JUwwQtIaheix5jDfznwzvlN9HRxWVCHch
cfMi1uquMaSa3HSETiPyaNnuJEWfkqF9pa8Iqhy6lnPER3770G4Akjg9MEPbTA+Jf0NowVZMVJNm
FeHrF0JmBAFbQ1lCvVMQKxW6wiXFQwgjg2zTgoeh3ejiXwxMWob6yyHYrAHfmZj0maFzu1rejG2d
QfLlJBWUsf9RWeOMAS3/MnFcy5oMZkiOlvfmakjRoj96fY3sIPuyPtIV2GGNrjq+A/06WOnvCKuG
YdYu8HwyQPSh0+bNRvxfIF+4DpyzLRJBeIADVvMdlGNBU6Cdb6E9jpYSlW3jR5oF8YMvRDwDJ00E
d8NITLXGOwnZOCKf73DG4osJUPeT6SO3o1n7be3pZEsjwxy4F08s5usa6n8aB/ySBETJs1z6jlj3
lOyEVSTeojuiyu1xWPYyxFS/79d2xsZCQVSWQPYUZ0Po4K93nWqx26c4aUlXIIoSkxNRCzuW8/Z8
LqR0bG/LJP5wzT1cNFcOB/wBMU2bdl3Xrg5iPndqvWVfidn+/HRhMveK9bwTE3/s/MACD+waTTTk
biDxNWtKsOkoOusPSlUrXeSFmmacr1fpE7O104AzGAMC3UmxbAlPbFe9mIWwV/SrB7t9hRqWiBHV
1hRhspeFQFSzbc91Bu61HCmk37H0LA2PZuJce6KrETNBHsvU8sVfYrESonPXQDNSVIDY13qrxooa
QovfPyNg4nEdvfBUFcNrXGmUojvHkdrwDu+RSeG8fH/DAtT+M2teww3Le3szNEjjbepuX1oZgr5m
M7bAAX+PAc9Tap140a7WUT9Cy3vD60O5y8mB5bz2/knZs9BH6wrhxM2DXjKGO1ULIWrtDhozi8OV
aed43td+GLTL8hKiLmboi6b+qV3blaczyUbfrWu4MpSQingf62V7EHAN3c6ArmTNdlOEMMKUY4ru
7Yjo/i2TRSrDulZhWk7HjQ8aTDpnbqgf6vj+hu3tRqNbLE3Us8CBFKEr9BWMP20sayuk1cXhqUp5
HVBbeFdEzKn+SxsM/VNTl2xk4Bl4dnNlUjA+ihXE4n5mm6AzCwZ5GT/cQCFhqArHfDnDqMqFlaV7
XswmPHARHqjRbn3nV75BdwKoCXJfaIuy88rDctbU0SrRaRg2e5HQqKLN4EKxfx1oo1WVAmfFk0WR
rkKpU4iLjZwNVQRVMAmsSMQnLPYI9Ou4h7VjKz/2E3DQMmaTjo4nTXUCUeF0wGN8eJJG/Kk8Mxj+
cJMbsiMp3J5vJ7SV/MKdiLYp5w/aPGVGKoUUEio7EYQZxvx9g4Np8L5Po4dLn8E+V6RQidVFD2to
bo56uZG8RUro0ZXww+RK7OTfc99b0/w/N1A4SD5UVeMwEBxA7dgg+U8sU6BaF+V988f2Jqjczohm
Xu5wgTI+tHqvWZBA2hm/p6e4oL19Kdd83hby59TSqub6x3C6QstWsFUdtj1E+FnT1WjabOHg91bL
SECNLq8PpxSFUkw3llpJmhRACbSkR2cQpCoMO5OjxNibP6V9Wwp3+H4J4oIdVHAxWfu206qQlElv
cf5i6k4ZX+RjSK50C8Jh82LgR6sFHSUITw8k3MSgMt1QPde0iLdxOI565TjK+lI7SlLHwHkkeX+B
UWSMj/7/kiAuE1KZ4dgV2ZZ9F7ZgOWF23n6MUMugvw0FK/gNGClEtOhI1TkN1n9EME71to3vZVDD
KIU9RHjScVhnYjpAhibYhgI+Or62i9W8sS116STwdn3Rwy3SYjqSwcwIQWhGE0xbVqGMtdHvT//9
tToaJ+T+0yxwhK5wOlgKkFgZ0pMlE3kME2dj1XtD4Iow0qyDstX4vKH6G9GitpsfxiCiSIv1zX4+
W4dnNhUTRGMiRg8odxBzkjgsP2hyuIgBqNrPTRQ6eanmu3wD0VkMiBgPu7Dva6/XF0/6SUETTRfc
3TP6EFwju6USiNfw/78gLfNsaKfq9k8B06eYEQNwWgW7r4PTkP/23rXfxodLocIcsLyDWLvwbE3S
2vNv0rHLMb14kqL0KDAi6/aVaANjFPQ5KwIGDmHBiVdNTNynRFZMuZEWqOqmRfEZPE8QeusxsxzQ
K04yMISVoFwjlUqD22Wy1j9/9OmALwrSeeuTcIuGyzwRSOm8vMZ/le8tg/t2B51qMr4zogHjf0VH
SrFM1+Cl6KHrgsU5X/wjX/bW1zH8wwJFeRYOfkrj7RRcNurDdQgR60405mHRvcKR5apGRa3ZaO15
zk0ZjMkCjY8lzAi3/Paa9+utW1izU16YHCaGAKqZWDu+1xZcsI4Yja3ZBumjKhJ8YjWNkVHREFa+
a5l+EPW/tevy85DoT+Y8mNJ7ZWbN82Yb571iB8Pm33K2IcxDH+KW+kF79KvzlxJ5yf0j25csN9Tj
4xjKyjuBctKvVq+JL+Cg9uA7/rFA/ceyS0g9YZ0/IvUK7qx7hCB4kbxM8blPr5M82dFKRBX0SB5g
zWMfvsO3OzpQP7pSgG4WzUzuwg9CqyYN+ylG1SMhFzRlTrwSkEw28SP9bBemykVCn1MNi/jS+Rn3
SOLzfN/hLyc116numATZbj1hQZU172NdJAYNEUbsstoCuvNyOO8CD1fCyDeuZgI9jjszKRVOlp8E
iDEpqxiSVxUiQErZP9W6ytqwgqv9mznb2aZ0alJ+3MBRIgtRcaejtQTcl06isFgsXUe2aM/BOjEh
HbpXSqVPjvcOVzQYwwnys5YIpQ1ijFTQemsRlQjtdSST5bGEUQRDkRMmAPfKTx1N7k+YKspg6Ql7
sL3Bs3gsiOAfjkJ5vTG8yogMfsn/Lmii1lidt1njgiXPWtA9yMIxZ1szz+7wZVqeRdpEk5ojPHVU
KvArf9hcDjmQlOHfDSCpJO0O+sqD7NlqST7cPOZzGTQCDplTeyfoWs5l1TvMUBIUcmCVbyOw2UR0
QCjlFXx4nrvokNDypj+kgvuFjzg26S4H3zBjS0pq/3svBU5r1QHJC588FhY0+a0q+o7X9vG4X82P
RnQz2UAecz8F8hcbBDXuylQgHVspZVxBqPpxjTBKxZStztbaLFwrx2GTFf91+VuzdvcAOR3GSVam
+j5W3B5aH+edPgBdDbJBLfVJ7xeJ7nABeccUGAfA3U3U0ABIweSyjYPDXC9X7Ve5O5AggT9/aamS
7ht7ukSstOgh4pjlnDHkHjRwXOpenEzVFLeRoSzaOMxq0AdF0Fq0Xh2wDIW7/PPhz4qo1slJvB1l
ODIRaSqIBKva+GNawaLeRStfAise9rV8X28z17HmjjxnFmuS/ouFzKKjgZ0QK0qb/nBzcJGJdeaT
BeY6tQaOs0n5DjvBf4A3iFDOsxlFSJd3Ajc8zGnUWpwDxCzCa+WSg/vrdDfXvBeiFAaTTKqkT3qd
ENWR3toQApX8svT4bxploPB2sqRM5nQthAe3eUdakBf9zusyumc1Nh+bilUCu9dAz0082/oBzx8C
OguaoOksRawyA9YX+mwOIQtaY/pwhJLGb8LYv5bDiSAP7X6DHgczKvd+U2gDfCKBrhgJ+G9844ve
aGJclEFzlZafgcWHQpNuc131pvdtO/f9EB7xzCGbeVZPfZVX2MRsQ0S3/j4XSkSgVmxV9N939xpL
jscMpqDh0DbEIRaK4+qUkT6oSNac15UwiOsbovJ9M7aWhsjNQW9A8mRJEceRFS4PV7O95i6Xx0JH
aIU+0QsPp/4KfFWhtMlLfnFkfzK1/+qcOx8Qm/3k/VXCdhZagnSKooFSXvS/D86Sp8L4aBjZVxHd
ux5d64sScRrqwtK7ytAwpUo8qM400vs40YO2ODdPvla/HIefmCBQkHMEb8EOc9Oi6XhHkBbVrpnp
9p9k/YgxDSeo09cfdgE/7ZQWu1F1rdsKNvmyS3BdKFhAHSqHhCGFHdrBo9ZFVgTPyTkArAKi9MjA
YD4hokvUSImmjQRMngoYIELrIRQUJ9KUZ98htuD0/av27wE6gKxVdwhdwzGeEw5t4qjn3cgi9yOl
aiAzVKThOsJo1tde6+z8Qaiu21dw7b6FZPjABkMrtoz6aazXeQQAf5Xy+ubbToWU3Og2PHZ07o5r
E9CfUvWakL4ze+BGF7G2eXOpPTyKFPMdUBPnbXxjSlBF2qRm3Bzc00h+Lm2RxXursoMQuPblBJCg
UvxBX8Psj5ZFLfxkKi+58oJGeV6gEtxlCxpwfM8N+cKOUfXQrZYn/eeodwHMaCcWNYGIUhdFJto3
VxexMVxxRlKp2KBLVA2z0OtR5Dwfbrn3mySAUbexG6PZk3KRumBG7c2zKiLTrRxolOT8nkOC/HZa
yUbwFGT3Ry1AWWOX+SiW4czKMSLo+qCnp2vSDnqmHkDEtF8RD00dlZ6T6jNNd+7smWPcE1I8EYIL
mmwsyRE/5MPJCT1SglzcZLEwIkqSF+QpLNHhxK4XWMevlXlnhTDh8uB96w+fcDK2UDxYxT3D4IWh
U+8VY9y8IjDsiq7eizjDS5GjLClckiiD2eAht6p8KRt2z8F2iCBQn5ah+E/eRA7fQUhEfVnYNM4P
7ZYs5aK//SUVoZbMG4q3rXWD4Apiq7AcyMFfBL6jW2gBqGxKm2comF9PzCFjuwgFV1a1kjA7Yhq+
H/WO2Kxp5ls3WHnRVAq7byRnC4aAVlV+SsWgnyGrFOgyB4sabcUS/DdsDdqwFpnRh6+4yaLpgl7Z
fXMiMSi6QJZRtfnMbvLPtRsfnKodXeo6YcN9WyA1xmxrr9L/MsM3Emq9IlcGQxKV+vo/EJdQnA95
Dea8gZyahb7vQZKR2vBXQ9RiD661nQSrKwZZpxwilyrDAOVHXiWT9xOIkI/xNJj9zu8azZCqe3uR
zHZDbB9B7SlUfNC6Cyz62DPnS/AcOEvYepZPW5lj4lKFMRWwXAHvIqPTB/kFMCWwaCseqY41P6fK
5LFUIRN+3IuztEazpEkDyJA0vkGDWI57thAK6ZCkLbP8PGvR1AlWGn2i9memP9CMV+TaLvlX/e4h
/xiTby+/j9PJwzRaOsk87oQpXHJwkKOeN6vM38yYoluEPpnYoFiW06CP0gRtyRkFZDVnSlQvifV1
JVk30TxKeHJVs86eIOZCihv1o/hhg+MwQJO6mks2Lj6zd94AS/MNNqPym9LOUvLXoue3mmbki8OI
ro7AUnu3T+Iuq009fDaOVfQRkDwXuRgmNXy2hROxZDBctkGgFkSE32MoDhaTuBNpRkivyVgraIc3
srXMgZKfK6wkvVVuHDzgSmPQou0tKXmkI+pLuj8fGIJrtbi7gozdrJ7odEpoh/xoW533qLxVzulH
4hs815dfw1sKcr7buZE2LumO0pefCBcAq6oHKuOjCrhBOzVyFOM1wj5rZp2GJWWyJFsKMe45aHBQ
jJhJdcKt2j9i2mSes2Y1Z44/A4v6GjzL+wtV+qILI3WKSuGM6PWSwa93h/GgB9+PYt9k9JXa8elM
lXb4qA9a5tuvz6WNTxdgt4672G9C/LQ2T/IgR8tUJ5ze5SrIQtzV3TFYxZMa/TrtF65XrtpW//5l
xx6cncoc1+tENjPR43STc9++iYMZ/Wja2Lrg+ljJQdpy4Cl3791PkBDogOjMAQkpyDTxQAi8t6PR
7w/2fWstdXPUOj3z/0RzrcejuXT2j1tmN9bjj8AlFYjKRbg56moopgOcsodFynMOlityr7zQ1xHt
NucK5+JOq3QO0C4dVpwH/pjdL0zumGeNsE4avb+h0MPeGw9PRiOxY+ncw8EEe5YXeSm9HjRbKyHQ
Ql2vJyMtY/lH2qShGl1FIsQ4cvkZHHal3C/QTLEr0vi7fgb4jkvBy87EJc2c0kuzY6Naq8UEah+E
YtdQdIJIQBhf72GFYd3TmU5QCanFYxCibbMthOZXJNtBn4WaTXWxc6c3+mtFng5thqyzV79KgG4C
A3xx4aax8bPlkOSjjzaV5fiKcXYnJ2uFuLfojwmmjkH0qlB3uOBPHgXkNM6xa8Z56+3oNu4wog6T
GBI0O/+Q4VfCDHU2m6hX9UfwwLkRrwW1bSXgKM5ni6n3efpOxygcTsQRr8FsRa1IgjNF33f/n0YZ
tWhzR6Bfk4bfxmrNpCCOWNis+xxE5Xz50ZQE0W1tJqFLLR5nHo4P+1jc6ufsrqkDDLv5OB2xMexQ
Af5BcB5zSHWltgXpnTQygdsclLJSvMzlswDD2fWi0U/N0LV6o1Br1HCC1QaQrJHmZO3T6BK6NqkE
7/n/2aJnDPuGmCBZf61w7WLO7R/3/onEu27DDshII6LyFZ21XuMcW4R+MxTVmQW6Fc/rzfshzci9
/pC00oGyJhimM0imdXUFVRFBmgYgj5HNXbdT8NnvHAFMPyKtEA4nKFtVIwM4M9R0j0S2wdTqlOTK
gVRVQP8tsAc5gpLA3yXvpxmMlPGNrU0zGpocSAe0wDFiPq8GAyq+HCo0maUVnEhjpreH60//1lrg
XSx60Wd8dgYr7BYIYd+bWQyZg3WFXjI/CFvptwnKQQZ73qCU5SsA4DUWeZUmxVOy5js9duwZWTGB
Oqi5nRN35r7mf12NcbrCxiidqtLfIzXDyOAJoLBMP/Z+aha2qMDXIanB/5N/8GvzgJIRi3LI7UBQ
Movtjqj0J3ggBAi0Cs/VkP64hNfMyAmeuOsrb95Aev3BfArImzfdG5B+koOWSLRQvFYi9DsLuP8b
LtoVSviugpVqmB8NalADURRbdlGa89oHDYLInWc9atYZkDonj/Cy75p3JkudMsBdp3Lj43tgtTOA
n0Coo5EXnD8fN8YarQtQGb+m9xHtyvVJFRDLarEiIkX19++cS8cVGXuu6LXphaXa8iWJH6AMpQYv
JUjDJZXUTtOUR5vTJnOLUVtpJlaJnIb14B2XkGXD7v2STEmvXNijWWqk0ayLwsrxB2DIqaBVa/xk
vMoBuQSUhRSe8tvbd5A4h87y+gqWkk8b8FjALi6+JqmjDWSJlweqGCgOhmo1iZ8picedoEfBXGyB
3v+eCl5iQM8IP9VZpYzGcUl0shJneTB61h8LT8NBzXXuDJmz0hJl8LO0SB044lvWLU6FWEaScj16
WODmY84lwTBT4jwWNYyEG645RAq68IztLrW32sQlsA1RuyWD7RzhBNTOfTdm2QQ9gknfIGup6Ssk
N712aSLqWlbnpsoTYEvD7dLdG3SonhHFFn1QybLTam+/GxKX6FJ6aZHUP/v2ruhWNhFrjfh5GQKt
1RItESzyYduGyQBgWZ0c/g7/5yiNhXbiki5EyC1Tm27rSlKFxyk9yFm8AqiOyhBMcF9/6iIcFOPk
C6QiqYg1XcH5KBaM8fvyWGmzWRzw4IextsBt7CRmzBA9TH+hsx6rD2MCLPo+Vl0gIZd75gPFeD+W
JfHLiHGZ40C5muSMn8IaxAkiy6FPyXrrTAKsKZViovI4PG+h6DztTPKVGKhjPrmnG1q/QCYI+ll1
mA06iefegAEVtX207GMsNzwGDFfs2uPyAhtHscOETmksgz1UYbW/26MoZx0x1OqgLXxSjU1gDPYx
nksemUkYKSMSezktNkXf2cxFBOhQzGBs9r3+ZIhUnOop7yB5KDc3h34OzeRqYJv38AOMRSKlsDFF
dmFPWUT+cqi9JFKnA4o/GC10vFI8uipbmG9jgu1HNwN+WUJFArhne3ke1rI6ce5W6lQT07adgim8
7C/L5HVHtJSd4soQNOpxtqiqhPLPp/4b8r4FMn4j/EBnKbJUoraB00fp+rs8Y2lj1FINqvCgiVxh
syaQBWmSrNutD2QIEPl6/3KOZA683J0jHQGwJJLweTpq4A3k8gQeDoRxEDbdfBc4T70pQ3QQouUr
2IdpOdBIAdDOO5LzdaUXNM6JDPcN6YnkgBPU6YxEqU5YTV3nUTxZP7eRZ+uF0VEvNGIwsc6Ji/a6
OzrX4Rfg8s8BNQpw4wEu4u/JUrAp056v0MCLmOxyRfM0vxYgSQ4VVehY6X35fwk4mbIEua4ScyGC
NRk0Qm0Nx3TP5eJ+QWv22IQrDegyUoGMb+9f6fH4+mAEhjcqNqjJ6xxFILA+czCFt6IzQWJpv8Q5
Zo2pnFN7kQz2wSWJ6ZTm50QYtQUm+d9S2vloYDOlXjdIqQvD+M3Sx+NGHAtTxeCY9f2Ix1u8oVhB
pu3bdIuyz25Afv6FnA0x+g32QSARw/Fl00QcWlOL1gwYapw+5enarzJG4aelz80B1Xrh1hNFSdBm
+/jqNsdUeFs9oksxleLeEpXRM8Pj1Q/5OjII1irdf0ELCOPC8RW6MrUy38azj95ZQ2bUYyun1/fq
6d2Np1njsGLkfQYjO9+APQEfSeNP4X1hFkAyYOM+TZmjkEkfBme1aumqABGcXCQH0KA+ECSwwUWb
VVH1hjhwrkGKxPBI7PpDs8vu6PKFNZ98Zctw/dTZMAt/6DFYvwRTIofKvGOwzZdrbPFxRSXgkmup
2l0mxec4bK2tlcmDe+bCUJ6HxNQ/AKfEsQH9W0LK1ZOnIFAxmrSe/YTvJ4jlrCNjog5mLPkCmsrs
CwqWd6c0bcbQlVddQdan86DFLVrnJpG02mTxJ3cFnT1uu8VeuBMRdgKUQXkOUGUsYQ2N4PIf1/ps
ckK66Tc34KSImb6Vp5reZDp0SyV4pmqDOg7oJji+5SJjrmXeOPZYs5xbMYH0LZM0ZUJFnpz3At8W
vqSuIht4yMY4VrQa8NVYqdtAZUuEYrpxnTTogYEL7OS4+bR67/JOzlDXWUuktlMqN0Ui6kP7dl9u
4KmxsBdqLg9WUAnb68h+3p5e4b0taE+W9VAIPp+nR2K4CW/prPLBdUXRwA6QE8c9CqDnQpBdypWE
xK2sjgxeWxxT7kCw0XTZqe7aQHLAAyUV3LOtujstpDE7wWoFqdMAkevWyfrpqrhodVob8vui5S7H
rLQtNq3M8ZMwiixupkOL5T/QdnR2pdgUIgCXShuMlrkeqHdP3eLw2D/7sF5/aqVoSTFsexBRWCni
1DLW1aCpsnXnIqvMwZgAWEUk9pVlo1ykP6MEklFCPec9Uflgr6vz1msXLvVNrHS53m0wshx0j0qR
eQn1yaB/2BnO/QBUz9jXnFfJCaAD1hB0D6uGe/3kaUg42uZDi8OA/X1dfOP+rmhxsnx01EBBAReY
b9kXcN2aUh+DuYrzSNOyRxQ6JQ36CORLIrn4/6rikVq2EM8UnipoboRTf0mQ7hPBKnBOHJbUA97n
+a1RWdEB/GKG+9TrL896Mq9oNTwfe+CwPH7jAPvj3S4nkZOQBwyFvjyZzCTg3RCZuyP1nwKbzzWg
1C1Jjn2dCXRUhgd2je09Su32jnj3+vK4Xbkjp0ckAbsbFLY0f4/OxujED7nPqJCDu0Bu6OiRBElO
G02++lskcXD01YK8AAVhuLzUDPVoAl0Qp/cdde4QTGafWzOP0gaUUQ8blrCkAGX7odQKFL7StAzZ
6ehdhW2WxR9S2LHQixBnKh8mUbhHnKlE5y8wKlXhpIxspem8wzIhlIxzyRymmHoS1X8Xs9rmZKUG
T1lXTQX8qESGXYgsuisnsvdllfVR524z9b5OYJzPcK37zZ1diSvRvXxCPtMgWs3ySbPVVRYgUn3Z
NzjLDYt9k5gicalC68JRCDdgIpbie/3UuKLK/xOSyLq3ov13WnUqiSrIC8LFFAr/qIbm7yAl5mmZ
ZWfqUX9VG+M19cCLoSEM+ed7ByJB2mbxS/YAcdPhTvtuECeVcqoD+A2YEHfQ9C860RIS8/BhwlUz
Q7LWGqxURwq7SCN3OaFtLBXF3kZr2XCmJGSgK2KAEjPOa3MiNqjCzthGzCqNbo9oa9t/+Jp/6d5e
o9zD8qTAhGFQD6JxlZ69G10wIbNiFQ5Miegkkj+Qdcbx9qm1m8a3oSm2WVKt1kY5FWSKw7sAeQCh
Jy6eNN2Hkg6WfZ5vVgQ4Q/OmezTmS9iOsDm2VrOWPcqmUVsNJgZFjliMFrx5SnCYWlNBm5n9WJ6P
yf2B2gxndqKEmLBQsGBnRPiQpO9qxT80rjKdhuG1LydnwH/kaKmRa0HndFWBrRlAzT/AHkQi7s0T
VXfhiLEmzqvYqRkmxS1LPsP0+ZkytZS8vvXDyCg1cOIEf91M552hdkctvDGxKusNc2IoTjvodgHM
ciOIn5Qk6dzpgTXKsAj2NzPLfxJx/8nPBxlO+Lv1lC23dN0yJZg120JREMsoewVDQJ4MUUBkVxLO
EucLIdWvPYc2g9V+RU95RKvcAIC0IAfWoY8fywMYtMLcroXlBc32+CfZtgXqVgvTAenk9sbca/ab
F6bAeOQ4KJiEXSbQRPJsjRcXCz/H6LP7gnsbL6FnGaJWQE2WTDO3UK4b+GuWZtLomd9oexbsgvC0
wp9IqbnSKLWWCFU0w5MsmDL6+zvDSweldu5t8CcxRWeuY6T/mggo6pLpX+1sFsFYdMB0lLEqL1oK
Qo5MngabeTjxlE3Q7a74d5CN9QBvEvOXakE6LbcUBhOJsjr8wpIzCc/UgjwOZkUKgtelUyp3riqw
+RuW+fvPd8GGi6RfAW3lZ5g4neaX750hzqkMKMeKXodLe45ixRKpvX8M12EUPiOgx4GwF2G6lkru
qqy2JKCsXQlyhvA56DMgDmf5kvfo3ksQNKhfJug0Sz+Icmcef9xDNsNmF6X9YIX3SUQc8JsRj4tp
2by0BL97TZ6HcZ91JErsTTMIlTU3GzOR2sxOkmMa+GfHtKL+/C7jJOAwlk4AybQDirk8b/9zy3l+
McVBEri+ddtIG462S0AumAjJ6/+vd566XN8tTQYIj3ZMUGeTPG02cy73ZJBO7+KicoX6FVIHytin
AwIaVNaw3T8/T6kWEIN1zH9BnK3DXVPgrtPm1fLueouQLflFVFsc8bv3+/fF8UkuEZOJ7Yl98u+4
7vx5nnExXvRD0GbQyM/QPU3hR8Xip22tesbUeSIt2ffXBpXzacKDG53z0T+ZZyXzvbBJMCDSzjJE
NUYQ0mRxguIqkZmXrFPKF8KOJckcFBbClraiW5IoOYjefkPwW6/rrXhX8tPrThAHthKFXYqqv26V
re29kdWvAV4QDzBekwR4WBb/AApAUsFD5cZ6ybsH+78OEOaICKLmWw70dVrNkP8v+qfj+wgorjdX
e5O3emMkPrFEjgWUDXxGa9VlvVdaOJA0l8OPYucSL5x8V+95bvwOemtq4KAIYquERfUT4sisSmQq
2lSoAcNxh5LW5wMe72HuXJhJvlonlz2DCZhfQPUYvqEzTf7x9cWQAwgysx65BrHRgmEsghlEvuRY
3+DFDetTralP/mVr+Yv5SqTNGexKtrPifx71cBgv9hxKAQiN+0W9bVQl/zK6ZBc6DTX/pVACi/S+
qb2WgQ8GJeyDwVA248uz03mhRk2F0stFy4XuKoVuLnvtQZ5uuCJpqa0l1B7KW8Hn6v6Zc9InPiXA
iw9m/KLprM+b3XfUCHorY5MjFlXd6x0+eF5nt+Kt4gfVmlBXEf1W+jrrqgguV3duKh/6Ve4Dn9Ii
lYMs5eduq9LG3z5gSktOgRNUztj7T27cJvj5DX/8UNxh1RUs6o30BGsuc8c/y9lpXq8zyjGw42Ue
dukO4CXItqjY5QkV6cfnYyI3Ib6i83pbfVnOb8WAXHZc4zMvWvf+mddnJ6ca2i0JxTQv7E4rwukr
jC8KNOHBCzwnwQrHkA3MS4bCf5VQu0rniBA3Mz5uI75e92aYSybfQyxX8NcpINy02NTJSD6WfZE0
KjKgurZQAYLUfu1rTW2FGyfLvPIlwEZs99DzMLLThcQKPlr9Bcten2LL78gNeanfMO2ScrKDqBBa
ZaUxLpe0Hp++crIyXs7YZ88zcswaqaMvaM7fbKJcMUwec4ioSAMaK8vXciIaY6nvWwQCeHxsjubM
rcAxB/l1pKOXzvJ8s21O3UrCUkMdOaS0aTWMG8pR3Rt5bL5Bua5yzK8fWBAsqSnNm2zFGZaC48rL
kxlmhBr0T5/lDc7fKdagn2GAKzImKIkv0fiweplyjoHC0iXSsUxbthAKkcLbV2SK5r+HR2WrXqYK
fxs1T835Xc054ZOO4vZ0YiuLspx2HY787x9hbUQH4nAPzKs3dNWSqySv4Ief0I6O9NrSUpn3dq4E
y99VzuKN3vz6AUFai/UuRLvluMZF43wlxuOXAmB+CZdVph7p3wBiEfKhHgScsBOO5f05MVGY6E3z
4Xbwk11oLiNwAQdG00poJRKKP/jHhkVZhqO646BE0J0zSoQGDd5KioxbY5ANREe68BMFl55LxhZV
Sf1z05XG0h0MdM/USxYGPLxdgezFMrcZCfQ7GrczxM4PtKS79ELF/UH/3bAolAt3ZpFTSc0qd0Gw
5RVAnK9rVaDjnuou8Xvo8mrq6JMBJJZCLPzh8Bz9p7vPdF7cuw8x17CRQxnwUR6jMbe8V/dganbp
JWXAZHevtwZZsqWAmQ0fNzZl4QBpD2KVWQ9hznb1dePIo5Sko9ln3jik2nou+kU996Rl5MPKYEXx
n6ht1nBWDOnu/U4K8AH71VA+bX1Q6a0vLV3s+JTwFd+2oxq0NWj1fEIecnx/bc2GuD9gLcCzlro1
Ejzd8YiB6rU/o0ka9P/meMGpPIVGp+dCsEMkASjxJxz96ZntsKLObt7URqyTHM2p0To6yOl8vOFW
MODwTv2dQlXnNCD5P3gtUQz3y6FxBEycasmo/rTYUQrRqiqsdXVcLYhMZ8Z8dPt8CHMF0iJs7uMG
P39tXgYeTO5TB7tl1ee6vciMpQmD4JIhoNXm/sBS95bEl5UWT4Tc4H99ukuzZ+3CpOcqu0l9UEdA
jizPdu6eNR35/evP47x9HAptZptAErhp5mtUjFaUNTRvi1Ro2uWczm9cDPdLly2ArvXtH275Tqr2
5SKnR9Q00sJ4pQLZZLdzLNxFqLMGLyRUnEUEKVog16MY/P5psKnCoqmHiLJJrzey670gZZxVbqOP
+u9HSgGIwdxXSQNll6/PUw9Yf27xkAmZjp2rB6ySJHkcb5H0fkNjU28Otuf3BNj+Ml8Fp+GBNZWY
KEYMUhtsYs/rDblJpxOPqxzP8feOBmcOII/iGmfSsia5sKWyY//38caLRZ04FeT7vYkBJ2boT0B6
06DUQt1Jc2AHkNc37BEy4a6spTm7VVGlWedsyq07bH0o0RV+NcHOGqiwje/15oazpMYBI0dm84zV
DAgAkFoBklfkJrOkRHUPcHP9smDAYizht88EfftdONLDrhZ74YiYsGzQ0X2TQ+cLdI4zAfKwNUXY
f75TgX4Excb3f5Z8Anxdli5FAeW6kDY3XhqFzJD9gRqe7E5ikw7ykzt5iNhNS5nAkIh+rKfY5vwk
N0tM3uBtz499wrTuVO1Q7+blD5r+3dMy6Jn1WJi5g6JQ3dWghqP/aoO3OSPs9cTPsei6oxLU7KJd
DgkCb10Yl0Q19dVm9oejyqWtRdD4EdlSBdkBWEnkcwxBCegP449mALl51gEHrpSeRyurlwon4B2j
VX0owfcji3shZqwseHSx2Xiq8ysE6s1cfBoGFCPBqz9ceFeaIldJl0nva4pPUIYCYgMutMhKBfyh
FSG9MH82Zn67tdiE9UgWodgqjcGkqn3FK9tDI30WKEX66T7exKTdp0I1NEVs9c0aMiE1APp5YH6m
a4oKVMFaT60iogNd/In/Nz0ZZ3xbQ/mbzD9NAI3fILvfGs2lE4Ol4ob7rzRW+36m+b2QrysN2LHI
5vreOF+bH474nRfKjxTPFIEDlCBDfGSiAs+ATIVrbRRjMZlYxS2tujGXf35tvD6OJwxv/FRDCjfQ
GrVDOb+RsA/zrtC/NI65c1xBKfglXJCRvtALboii28Oq1i+10Y1k1DqGnUDkpZ5iviiEO0atKQKK
lz0u8YRRlRBvQ6FA7MpXZZ666O0FthK3lNxR5AafMT7TgYM/cmE/pOpiUVWM5Dz+InalgKoVE85V
m8Si73AzVU+whIv43j9r284b57lxIjqfr16liOZXlWPXWGppdVS4jVEM7P9VNpzgHui74zd39kcJ
/wXrb+S84DeMw4vQhgKQPadzc8YtV+lhB85MjZeRYPUozqpcAWhdXcuQdU26PqcNeJk8F4QGpXiI
tPOtQqw+OHU25TWzAcOaWQKcrqFUF/axEt/9PrNEycKp7wngNUifoZ0DYiEI98XknPTwvHCMgoDj
3MPyO7zPPuK+za6Dhv9sTD2h9AJOSaZghygDwKlbrjccuCNg/yDvmetYSs10C20gzMF4K/XOc4CW
0ju7BUEbQskc62XVEXB1G3oRoQMfjdAroenETzny7Y2gwbX/jPSDIBxeJhrfc360yup+i1sw6mP4
6yaeYnCy7rrd5/daeqycJZBNaMZPU6g4L7AlIM52vkNlB6moDQtW9qNBP0rkC5RZyidMyelR3WFP
NNyvD7WKSz1CgqDkmTMRlHcEPVa29QVLTjk7Y6g5jiEL73qNJYMLrrV32NNeSnx/oPh1ZNnnNBNV
6p6Ueh3IjPBRBgE76/bRs2bcch5sgUrKxRAMoFzxE5pNbhIZLOYVYXlfJB0LKL9QjcNcbSI9lanp
qLAwzkolVKKgx6sPfxZjTLJqfrhTCXZL7yoW2+NOBquYdyJuqOsM6AkJdP7aTGGG5BlSaQhv9vvE
foL9N04q2noH4BkloJGlWxGF0Xlh9nZcfJREOTGGUdAnUDvrR+WQ1u48WlR59xppF6CjaDAe951A
GaI8gu23IFV2ySzPX3i9axLb2poz1uI9INsGjmOOoljx9nrGDS3cZOOdrqJO6qs4yudK0ZvpI8cH
5KQy6F4wcBuVcKY5wCAirl4mJNdPfpGQ7B9pgXAx3ptqR12z/O9Cy62x47x/yU77veto48rqzNBb
UDVpoWyHfg8Tan1qr8WwTsNdCO0IJM0cJBa1YshLDx7GqESg0Awp1fIMtfr2F4NfCo1R3VpZknQY
jsbErrwzekbhHQuwyVVdNnUj8zkxR3k5iKsJKBPtNZ9izGUF24F3mz4aJnXGUv0uUv5KMS4BCBE8
hKNXxUq64gwVNY0R13BKyIO8pJ/RYKYYuiorR1cMwCj8L1Kt4MHjAfnf/S+XcRwAOY6DQxycYOci
onEOskV8WX+tdvIeG7e1RlZJ5IDkRB+hAvrJiknRjVGz6MptYJam53ZOmeKNN9mXzqtJdgrcWzmw
sPptZyqbFonodonusOoi+cDV9ZbF4oBY4Ecx0fFgmWl0b1Qkcjnkcgs5BaZjna18WCzibcKiNpM3
cZ6WmViwNmz2qVDQC5lhMMY5ZPtVi4SYJc1DuHNL8uR/4rNaK0+/YQQK2pg2miJkEGuwC6SBXnBx
gTGRsWhXcw95bVTxkjufhbIxo4CJRvMZV+oSYCafvBgmo2KOOcKNOPz+NNsTwAzCovTdAii9sDsf
iL5WHkXV4CuOYWREPKy0aYu/d+P/wjf0JZ1cxuaresPEs9/YbDXmDKMNEO9v3GAe12YwPZLQ//KP
GfUYseGjPi1KuP8qmb9ig65WA6ak1RdG5m66MjIJT7YVt3+bo+PJ59LbjRKlKJOEkrRvc7i90kN2
V3vjfxLeTRvymIhHjeagb9JZFasr5sfVejIoUaxkLAxOxSUJ/QB/NQynZ6Fkvjlj1tW5A+ACovtR
jHp890J7muY1B0ZIPnMKt4ETcjfq8glsOit1OlxxHWY+MyOt7ruPPG0AVCy4Z7VnqjA9jS5mdu8o
mo/vEOMY00vCzjNdJbNhEouORcYiqHLH8u4K5K00k8/sWMdeLxml+4nD2epLQxH0VWUVvqTWtUBh
wT1UPpAB6E9Jh3yS5C86P/z1frGZovin9CMFGT0vtA7VJhBz3xLiA6kCE6IY+333oyuG8I3TLCNm
rmjSlfbdPwFz3oq6pF+dSHHoA3jyc8kwsMzNT+NyAzphvAPjg0lasJQhI3spje7ZmPiNdH3n+Y7R
Ql6xxetzPhC2f1FpAul7Gtd1YgtOrC8GY41zDSueXiq0CU91Q6GWS/uIMAPec2O22vYcDuxH5z8O
uDmYt5D3/CeJVAs/5k6apWmQGMob+CnYSiubmpuiiQch8gqegZQsUyXDgP33ZlNxwFGCCOu2FuMN
uziYSTiNP1tlUf1QJufIb5VlK2ya+0piNoJIO7+BA6HzBn/ZQiJhM1cDCYseRWQ6z+0jGWtrzSm9
63SmuoY+TjSv2Ljvc0OC3w+h/Q1M93aNE3cKbHhXVZcI+5YGmLbHPUuIWVPRWXBKVU8XiiV4ihnY
tdJ7smhiRYRLx9Hxz2pMhhE1ujASLhy/4BQbganIVs4kE1DNCXqJjlwxN/uaffktaotapIRILvrj
ZW5O/wDVGcRcyCxxADJiTBA0Zl4oVGPobwa2uKlg4oEoViNB+YeJ4la98m3RBe2TgG4SdF8+yIPX
KLopA0T56dGzTgU+nb8MC4rCtX7CZkuaA0fhTKVm5+jizIxXeuB7IRep6chKdG8VhgYd/n60EpTu
3+VFwaqn38UQJhVDDi1VELgcZyjHFz0cwB2QjxtU9JwzftfwVPEK5DJ8TghSFOX6hJD2Rp9sEslU
FieDvtmvdR+fyBmirZRQrEIn56tOtp/soY7eMYZhZV3sXyZDBVL+S5biZpQDYKA5SXpoBjWAL5ZO
fCMHjSqzB5RGmwi7s+DzC+a0hMN8BCEU601M1Yf3xWWOf5NGvTT3QssYrIRYxFvrvd+ENYzVjPF1
8w0TNtYJkRSKK9P8DJ0kKi7cguJ5B3b19mDUxQli1PEH3yny74plpKRPQmnhLAp+HGkGba1kdM89
9aIQS5+VPXSz3cThjsqEnSUdpvlKlead8ZayUfdOJ0QtViMZfwByRRrNt7DQooKx9Em74RPfj9Iw
6aHzXjvQDVgBBFZDoaJBdgMpnL4ksSBkgw9+egsncwIZG37eqdjIXXVoZva4d2lHqs9LucHswad0
49AX2+Xf/LJ4GB9rwwQ/VbDINnGaHg1pplt33we5riBXhSMkhB/EIzlOzFeGvVM6OYthXF3NLwAX
RWBFbGBrXnrdw8+5fL3QTfgXSDQwapnl1xi9NQUDM6xntL6zn1l/AaDS2or7sVjroiyksnTHUZg1
4aNZ77od6NXYKd9g/5Uw0kwDxczSDjxgt+AKYwk4TzrvxgYhgGYOt1mASoQjMOaa35HmiCdKVtaP
oXTQSCa/DK0INy5bXfLafJk2s6NKIAHo/pekfojLdvzixpNjpBwGIAtqWR/Mw/U03OQ4m/Ymdq4W
nTU6bmW7leB6HocyeANCA0NCjuloyiT4/+ecAK4XxV87J4oczn/gYrgEnCLNlDCG3ho31A9tBPhw
9M1DiN/8Z7qfxyCJATRgLteTCezkpCf9esA/9KLA3fsMM2sWfefZpKTVRGGdUtuYnhYifp0DDtdA
eUw32alCLja7J+rrUGHTgJ40EJWiK4AMTk53E7kG+tnMb1JkRk1RAFde2wprlfR3W+8jDcouChQJ
/G4nsP7nZZNYVEdxcOMG92Y35D4SWXu9QtTxrfrl5eq2IJN5vNFyzfyxFUjC96nx3Cjv3nDoskSZ
stFJt3/88oW6ueTq2x/T8EBDMwi8cHZAx39wGZTSeZ01nRJfpSfRZ9viYSBqwCOT738z0QzUEvU0
w6l40Lm5yXCWPc6Gc32yy26QzZzro+V+JpxRFFDA7iCd3f3B8meZd8x5M5yFSwm8PtVH+0Fq9ZXG
pVlmnBlUtC2wD2EQJ8yn7gW2JjMYhPrYhJOi21b74VpAtDgi6EXVTd9SOeAweQI8s9pE9dyMg9y6
yH6oKndzlrTRl8PUHliS4UmVUvKqKGKlnvtytnzryMkoboxoIWc6dQFw0ho6b4tl3x1oGXJs6OBi
WZ/R4AuCTJRkXBUYepucp3aIRj3EPZK0KbUE5KnCaUWs4th6syFuj8F//JKmvI2ofSFc5mHp0E1w
eK09GzqLLVANjUwGipw78tNiHFyXKMRzFzbrbFmUARlFWXrUBKmS3sw3VAfzJRUc3/XSlQL+u6OL
6AOwE3XExFvDLnLMUb65No4yjJw1nAqaSWDlt0xHZv3yrZEqVOgHyDOLH6Ne+I34qLtYVT8bl/E8
ZHwKmhIBjE7aTmQZyGHcKBDGxi9O2O02MD4HnnDsJzbQznTVWHHQqQxFyIhWQkDU6TUT7giSb8WR
4q51KoCpdb/x7HyRxzcIvyHhcIAgwFxoQvGaunvmo8TuuXuFr+eQD2zCxuVGcGiHgzNN5w/l1pVF
l5OqEnvZtz3ZIlqHLMlPkRdFo0zHVD/n9lVN2LcWsMCqkeZ18qK3UWCMlxDh0XnAsb79J/U03S3G
6xUoymxAjvCIWGiMFu7A/0dJGoZPEil9paPzak31eZUg1oukv1lCxNus9O94Z6sITYmefm2Wj0Sz
xvOBSvVNDnZFtXoRvvV73JdpoaPelWcfi2wofwugqctspEgPOc2w/dB/Ekjj+znmYSPr42cMqnaR
jKOzK56pZ+jhOe9+ToK2hKlGkRDVDkGbExk6imyx2NCDySrYUIXVlkJM2px2kASnojFTZqDX3ps0
za6qhpwekkxaQF4/4yPdi+eIDF1TG/NHH8zB2v4Ybiau9oZvEkTmBhoLKJ/SeairQhrEj7Fq5/Oj
oSTy4+ixBPMYCiY0GSJf3ARIq9ZP2S3pckQwSP9Cgt3qtQfj/uaUjDKglHA01jIWKKWPqVzPULap
MxLNAPsqZ8fIpFOr7aMPxxIFwan74PJ26Yh3ETCHmKY0C9lqRw7MJHfsZ1nQ7qlao1xDrioekvyx
+XFusvLKvvgRoZwsDdaiIk7vJ0whcJRsJ/BZu7BC/J4SQoKPN6CJMj5smxWQWPPlGhGSqeQtGAgf
K1Ire0M422fCTB8mpOIQMpUoiWBFDbFLeD2aYyU7UUODukwOlZZaYvgCdYTSgAEBd4HvbijQDutt
+b+uGs0o2IUMdnO0Cd3MOjYAHwY9d0uFGGWejXaTpzyKEeeF9w7yIbVJvIS6t/zo9EZ5NLEJfr3S
tDrAs3aPpFxLfoHvLktSdwwMih2LO6ewrfe37Y6nyWgeqdQdsN87tklNyJQ+u6fd4EfRD1TJMH8j
kE7X4sm/4EacJM3V3N3Me3OhUjvlYgCh12775fD2NHnlKzdzLgH4sdQvFAHhaqQfsIDnYJjeOxby
bckPJUTBWKQmssyaJjUyWot4PhjaH/2vaoNXUGUIgMSCu7UydV4Chm7uq3sFl4ALKxGpL7wgZGrr
VoMmLcBB6i6cP/PmbHBD72KV5roqfCXmWa6WqBubwto7gX1O61UuSBGjOKksF6u9qlNrKZZk2y39
6lJ9tyWcRshuddWa/EuhIsKhL/IITL3+TeyNqw90wWlaQqMmFLynniSAG9QbeMkSjiO/MYelOytb
jtqBcb/rFbbS9gmrukmmPuAtpjAEhpoM/Z8TsDMw6mFr9n3Gfgvp5jku2S01hbO119+fPGj9lOWl
rrd2iblMw1xnD7XsmdhaDLdgw0439MkQK5nwLK9vvTZ+TZ8hGQvTNy8a9DE1rheqZhsQfzs8cuGA
J2BYk1v4G55pcAph/4JmNAe4pF2I2SFknklqvnkWsys1X3mqvj7gpeXYtkHu4ZY4xV/62poT4SSD
19m2n1MY3HmpEoTIYanTR7s/ZedLFQrQX3uPtWgS5oyMG42i+BtfheXkj5CusdSr0stwlUV8u/pn
KyoP6ak0gqiK6yCAVBvLCqBiUCaGgJfP2ggvW2mbhIdmuznPDW/+r8JNlsL+uX0TZ9HFORVdBgEU
i4A3IRlOUmbnGBwhTrzd7RId/i2b7J1Lta/CnhmjUuNrow5Pr+VuDh/+lUHo7Tm2Qk6SWAda7z7E
9sntWjVwhxGbJvuBECEnOxAxP+405YLiYIZ6+lApbZkDC+bjawRt4K/4Eyxj7EOwmxb70q8ilDDV
dPDR96JCWMFOzdyxn5mnPYH4gClFY0ZAXTlFQHERdljNftiqOrnG54QiWV3HTjHY/zP9Qi6D/jF2
6a2PWwElM2oTT6XJliM/CER9IL5+XP6kOvnVdpeF4RMglGvl285KebGhTS0UL6Gx0PhTb71uXJVy
7MD1Ob+4W869dW/SdMfEpvqBQ7G7BlmHIYOtQV6ljZ7vON6qcePDTznKQFTIiqIVhkuH90zrNfzX
ZKIZbzM43wpuqtlHoy1brHYA2rzVuiSBhDatbxjFwwzzxAhrjCEJ6b2nu5JG9VuHH7EwQ9d/cFcq
C94EerNndlZAN3nT0ckek9yLfpWPccTvbZFkG+bxoVOTPRnDERTXXj8n8UdSE0IqC4EE+4XmWx5T
K8f1Ss8ZO66f9CI5fjiV/jiA2kfAxs4BKTGnsSiiP9PV4+3EMqsfozocNbcEux98EC7Q9k3YiivK
1JTbw9SqUG6j61j/OGzawpXjqWP6Q4euRBj9NZQMJ3rqCQlBSzjQKoeGsmS14AA+VN3pq4mnAAVA
QStoBF2N9VRNYxhNZcskcXrZ7ZPmNh94/L4XUZ+TbQZxJydepwykp2JzLXa85aFy0Y534oSgdZs9
4jB7B/kBUIXVS8+BnnWA80tx9/AfnfpKpYCNQI9HMN9Try0ZxExROCsrgmH73THGCNr/u172TYwL
GUXHnbdOseEbD7WV/aAPS6nb1Y14s0Cqhj2aFSFu6WqedXY+u9fx6t/+2RsnhlQzlXVCiHOwWrUm
9Ty3akMBGEgxkCCWtBuDYhCQGluymkjdHzCGXa7E7+GUGJHHqYpMh6MxBKBb2fN/8LUjHBmEYK1R
yCiJHo65MFZaZvkrxKRorZvpdfNiBTlSZMUuK7VUMUlEraw54bx1b69Q6IQddXj9XyiSNDL6U6C+
GCCpHn39/OzGg06o/BY0ovBXDk3w1HzmPZHWHO/wTnvoVm4Lr0HvNp2yGrAn+K/YccJ+fMFIP5LJ
OsEchWEkSakTnSkp58VMATv1IuVj7C5DynP9J9oLrg+XOHJkmHdwVVmtkvKuQw2fWuBbPWJ7pD0Q
prmo/dvcPKZi0dnPIoUzHVz4CHI2/cLkAdFlBKGjCtFJT0rZcrEykYnxSZynXkdUjz1b3dPKu2Q/
9AsakZOV+MVcQMMlxchnXmtH52A8ukNto0nU0sYse+yi4143Lqh6lOFUf721sIDSOhXLHrihBpdl
o8WxrrEJ03pvWm5j5VPcriDAcxRV1VFnyr3K4pcLXLNCuqMpNOEyONkg1SiE34XrlJ2rMRlFoL8B
9QjdF+o9h/FNMc8A89mv+Xgv8UvUpLMpQdGXiER+IX+z3S+GFZ+ZtIcVQyxwv8cFUhMElVBHZNk9
G9OXNTHp0aTs6LoQGd4oLg7f4fevKPnwHcEF4NenVftI2gQt8Nx1FoyHKQHeZuOSlFUI4gmCYdn6
M4OatSwKUKNzOTMYjmrE+dvhQUNuYMbCGo4upoLl3URrspPyaKiyTCTAFByvONEXi4IsrxN07Z9M
bNJVTuKLnv1No4BOUnfhqbmwa59td6ivFgv05/uo/QQcmBf2D50/vCPkBjveILZddo3dUbvSjOHN
hNHuN7yZS67pBjxLXtrZfBcIAx3D5EPPs5YHhJKb41br5keh7sMh2xKJiyk/xVYgMx+aWAvaQv+f
DQwkn+D32zTyGHVFPnbSihvGEpQgUDbFatzaTHBkDlFR6lklNws8XD30t732K2mzKpe+qOseEw25
YPVGqCdDlkppLPEUsw6XXTYivVxg9swamGnzzmTQZ48KtReQ8yEmOX/cDSJJP/lB8ks9cL2noN1h
JLpC8vRoILYdwVB95+5XpoDB0Xpkd/nYez+9CMq00q3+ErBRX+O2quLFPy2tB7XbX2dIGqFZW2kM
PHaSwETbKZPKG+8UolzF2UIZOWDWJqTL6otqxQrJS0maPmhl4mNj8B8SztuXMIKvp9Ii3G3qkIBV
ZasD7mvEkG3IRTykanxVH1h2qIPEd/QMnnk12bO5+PjxMuIRssLbmDBoiEnWdLvwNUE4jwfyXs6i
vpCyo3Z3//RT/gvjXSWJzxJVYIxGQQvN+NuvvYQQfh5oj4t4jLlo8ZXl6Ofr+MtARiKNnzk1AbUC
BWUrDkeguLsKsDFgaq9EzqzK0cysRYstnCUHup2sXb+Oxi45yzw6+Ivk4IbWv33rTcmdVsEU+OvQ
+uLzgE1rv+V6f62Gw7rFmYwNw23qz7/4fPNG5ZRAJlJMpNkVFfgcywspztdNApedcZrPgSM0LTHY
q2UPGrCob5uPRtO5J44Fm5M8VUB0KbauVhfAwSbqbgn56W1mOtSXajv/q1zcgcQuhuw/85bFIG/G
UKZet1ersSkuhpUfQPH7VjJe81Ua4gAp8Ytb5CcSbeXuws1v6jJXTK/1zy8GLUzEcuBVszfBuobD
r4oj0Ono+wHOw3v38gBtswTCcQVqdY2IqZ+x7ScZPN4Ok5YNNXdzmOB/0xknyzRE5d1GUejqlcHf
nl1lAjycxxWOYpA8deZ4xptUbZIMK0brQXDoPqOdOq1tMh9KYthY7FGw88qvbqAjE+dO/Xndk38K
5CkZKHsCirjjiuAgsJLNXXjPqZ/31dThdleJCTDlRLb6+5Gt4acKSKcoUXbWQi6NGvR+RTvIzNji
NW7Uif2tujW47jfgrp6XxQw7icKILqModKeNLX8UyjgNXI95GKtsBIiciYQxIl3S5RsetSb28VNq
Qdo1ITDujvFJgLsttWWaRdq2VviN2FLZYjOGB24mobc8GPXhx1DoVtKyKFq8EnN1OdvV0s19OM8h
x9gzYnygpR69FYPo5o4GBAF+8n3OPdliJBZY9o4Zd1ON7KOnOww79BKuKZht3vNaQTFjeYNZOBit
GNUzUk4Gyrv+AVxba5lzz1JfoFMOxG/Gsy60kQA6x5uLAov25g7ZDCLZaeByLhjdc2gLgP1E1BLg
ijq9T94gVcvZdX4t8VFhUrEcjasoLAhJnV1c8Fnt2/d+x1gs9XeacnRv3U1kjOO9RdZNuEg6jWM0
uwURx9BJ3lljEzbsg7cciYK9PSaNni+iCU/etFEyDBatCmxpGHIPBLWNNRSVhndv91WfHk3f2MFE
3K/h4oz1bG1rJWG+xPsd8GtBYHTSRbzKGjuXexpOgqZDVym6xbOh+TMXMqT4EgSFXBNHz87QR3ME
Do+hjaxj9wa7iNo9eqvSef8PmAh6eoyuBjuTV6S8rXJNpt/aFYZyhhYyI0VwVeajWo+vutUS7GD3
l7YcBeLmHESYSPlY6d5gZ0hfyPnlGcybTf0c1K0NEilXBmnLAeKdIJA0ab8MFDB6QRxvZCeT6i14
7mDErRDYDHwYYDq0qqCzB+4or/KwIF4Y2sj1yPenNpHplROBY1Vt/piNDEXPqYXXinQ2thSldBJZ
UEP/oFg3chuCzfkIWRD5WreHoetvnJhpKP/KuH0wXPE/H0affoplbrP6Bgm8hlFU+46Vj3e7EpZ6
D3pbUNZmnR2MwQpMm4nczV26jN9sY1tPnTyyMPP+/yPotCOcm+EZFr04EEyaMXCwCBedRf95cMx/
e7Psy0GxIGZINByBsxeSd4Z6qzWRcCHYjOuBtnYdeGD/WB26sMzg7rvJGY0NhTiARjqFyh0/y5Ci
ER66Iscvh39NbXYxfd2pmUKK7s0STSMNVPmIjnS9zYLA1Xm6OcedCp0TONCGnYnfEsjVWWDtsWU1
lxaFCQVer2cBQQIO/T/lUGC7GfCvZ2AwrUaZsHzdvHXoZYAbALYcfggNnblKjonRbwpPYweXI9yn
dfNxAS1zm8axByaUARS3sfI6q4wLtRD9xmBWG+5wVvyGGin4emKpsuAVpDQqEBqyJGFEWJQ3Sp56
2AKh9MyHd4vbjt8VOGn2DRvMXQswqPqOxKbAhzTcCUNadK+6nLZogtJXQMHO4FIIOc79UvGazx5H
3h1462XXjdnGB1sO7uqsr2oVqeerAhJvLqhLGCW+Bib/NhMLJ7IY9QP2V+fdOf8jOIeTM7IGRmSK
pP8ewpnBwu+zIjm1+D3CS869vXW5VYdO0raOAPJR05HvRYcBynDBQpTZ5yYDSdnWMr4wW8w199sO
aHzAuPBUTae5SdynWDjuWlZ+xIxhIM129tuh/DCARHWxWZhyxgoTVW3HPO6heR8wKWyP2TG/NlTD
b2bRZuLJe3Af7WyP9QSKf6PrJQ48rhNg5QIEPkziKVEwLxvGEvVj5WcKFvkZW69y15gha+6WP9gN
xzsf0MNMT03PHFNzto4OVy0iYdszhHLXO/aK2TVJ7s18FHiXhY696rTYoxFHCy3OUkRvuaGVSHGb
FuE6Lj73hMv/mR27SFTJn4ios2ydQRGcgivuDSxXWHMcknX03o87be7ojVuZV0b6yakLVkHeJEwz
jQHdZLD4e8CuJJSiFbUIk8SHr28LxsexJygZKOoDY/vDRdYkz/+yA89kAMt9oauY7togNLhhdysW
Z0sD6C1hgJ1yYwCFFet4o/rMfShxl3SZBG5I3SvNoocbDruGRFh8ANHRRX1XwBMzdoQn2BVvNJLg
VvGaKmEUm86YXtGN8g5gmIICQq6iAXkaC7D25sHuJep3WegQn1/dsLetS9meLI7YfIW591HNjn92
cpmlKDnGzJzVG8N2ZnU/qKuj2YzUn/N+ZRHaQF1hiCuBTY++bBgK1rPRVCTvec569mzaCnCbstkh
qqTzyyeZltpIIa405yuiMh9DKOmCXYvoVt7maEBt1Wz+lr23feWq8nDbwNHZ2HoOiFpSguAhu8O7
Ucw6K1Snqyp/6qaXgws0jhoTbmwTohizZIyjZexBLfLYK1/e2TRsxSQ0+M7boxWGQJsaco5gVbjv
YkljlHhKkgR7MgN7iK9lf7JCes+P/0O65J5IZKG2HiqmteE/7de9YUlPXzIakg8g9larMvbQNgN4
XDs0w9iE7PczUWRC+B7nTSJj2kr1KkT7vP9bbOb5r7oZl7/e8xoxAHtOjva4EsOz25/qRFcOqjRA
UPCb3q3yku1HRdXeOltbpF/74vb35F/eTJ7CEbabJtUbbPNSGOgQyIgvjGm3Jtwic37x+bOD5BW1
jSzfUygYLqv3yfjuWQ0vLcGXPD9RORilMN9ApbRFGS5RsrF0ZpABXVSOCcolheubsbzWGffNN7e7
/CPPX0CThwcs8xtCfxepTBvj4PErJkx9WygmqVMI1/7S+bbXiFRbNOOXxEewwqNtsTuIWnJkPylO
aveJT9DqYOqZsgOiFprL2E3AUmOQbAoXyA4fzhUS/7A1eU2c5FZd9zg0yFyjVstiEQ67D/sDJ1na
0go3klUo2Tt1BQQj3a56KkOvFdX/xi6IM9Bnunu/0Y/p4RgfhmYqvDTAZ7OXEenCfO9JwATe8Fe3
DJAMUCSTcS67k7PZrVpnBsbbKm3TvyfyeBkmnYwV+rNtP71Cl8ZOtfZPslC9L0W5EqHyJc5xdzc7
8yu3KqAXnZPgbwfqChXs/ySQ7IfC7eTnZxGl09cJ/r5tdObPxEjCFZreEbGOl0fGwjJfSjRFHcwY
qciQHGYA6Yw3OQ8uJqaDBCAuv7CLj170mC/raZUaHXSxM4zZ6Bh+TKTYWw7FT+MJIoVZ9z+p6wN+
FP3by/8dn8LlYELH2QFxsjpuQFWFw1ykt9QSN2LRhsqtan9OoPHhJRPqhpwKXgqSzb94PQBCqURi
IsSjcJfRJ7WGA6I6zVn0NwUgmIEkN9sxrPc8ZP/q4OXo18P4RH1jSkqE2CVjehF9TCp0nUw1jSUJ
l+3ruHdFo1U+A83DMshE2ItwiOslgYRGu8OUNOMCFrfX28oI5XzM5jGDwOdy7lTLt+JrCxTh7x6Y
QtwdmG/EFNIW9X3lpW7WHKfOoKlt30Jup0DLIxDGIZ9ljTWXpjBMPjzVCbAZrSEaRsi6z5+iH2pR
35GDqp6Qurc2gRu25qSywteR8tc4hPwZ1lzXxQWfnyHFdMBEBn+0dEaA747U6w/5K4nKv/4YeZpj
gHuAGfg6kP6gHEuSURhpKxl+PumC0VaQ4PU4xQKEpP3S3AOJTDM1RdyldIVHnTnooILe8zXwHeS1
JhDeVW37BWNLpjdck4mrw/loncyRlz/sFPUddu28bASfz+qHLaBva6xevvDXmOyvddF0PYLdWje0
dTXV1gz04oWMkbDV75HOuAe8QMGy8QSYmtE8pLaTIC0WjWWmNfdv8HPi8KXbnEngPCEMka6x8bF9
WRHgozoSEEn5MB6Ldv5o5F3yDvXs6RrW5tsNLK0X0DqXaS0d08dPJG2+WG46RAkxHxvSMrDq8AEE
Ir4aqkmsY6GkNbg60LxU+PF5ILDxgbxE1LyqVKmSMUGuFVbfrCIwbGUsMlnwJ7UlF19YWDqFXAol
dSQq2ugtGHmCgG/+Vljcv+zIoKoRJFf3g7iuYnomhXBlLSSezqyCtg65EKvNQIPxVzkkgZCWdF8j
TWK0jw4cwKUZhYu+jkwHSgfHFa6GlgxySeZkacTGHAyYtPw/vgfDbxCaJ6JXJLtRX4O9lExWk2th
8HmTemYI11rpQxKC3WWAuON3jZUmjUEQN2j2cAZQ3eN43mm7WORWx3YFtt+LFn6bFtdu7vrBjOKs
OBcvKJCBq42URUsHO0WRyaotDzCXzkTJwnAKIJ9F2Oy6x8tgK7EFh4lCrVAPknQQlxMIUCWaKl05
QnshVwUgL28pbE7VdszpIwGQ7p80Scp5AAHqbdA8ZKtIUosQ3wejEANvNcyusGxYVYUUpx0Vxiax
QC/TqGyM2Nyr+oMz9MzvoC0eUMggOA6n+9VzU9SMmQlH64ae93rBF1xSK6AXf1P3KlUmwCkzIwGS
gfptmVWwrCxralTNvkBds5XLcPqqHkvhM0bvUgv3LNvGsgn3bciy7gYKN3SC48pS5JheZXE9dUmz
OrG78V53ZhEzgfB19OTpQ7OFIPs52rJSfsL8BV1QF1Al4BcQ6flUQLpVL58H1jHNG8qWSKLza0eo
1+UycJ0jJvJhUHvQ52pWgIOceQqMvI3Jnt0CNrBmFqxa/kQBq1pJIsEw8w0270Le+8vW4rlmj+cO
FGlYsHSAA2wmwztUsWrwj8WGMPSWNgPoHjcDU16G1nsM8oiSs17psggQnPsBskh4g/seJUTMjMhh
6MATeRNBtuW0DdSRMUorGn7Gx2eYcZHxuMn3L485Zkib16Otp3bUNSKETw07OmRNKrrorfUMtJig
THu1crkeEAtAa+TjDymapQfHgiAFggBe0lZWejOf+IE7Spbok6ECnMdj1+0REJYWIW5UKYanZ2g3
nmTfPP89dV2jy041YGjBQ7bfsI+umFtj1TgBhNqWSmOPc0WCuS3j2C/JawEmIOh+/Lc0bFr4goiK
etMgOXsC30GJBRVkfbyAqJ9gXosU/CELZh/JU/nNmh5e1rD4v3Uv4yLaW38RjxgmyuTZENL4yE+m
4/DKQ1JISp28LogbqiKNYMu04qsOP2orGvep100QwwJ9dlNzpOZTFAvQRJCAUqrjwIIkd1kecdyl
fe3NjIwIgobknrT09Kddo6Kavj116KywceKn+20XmC97n58ieSd48Ng44tgqdlgzCn+eobMF96ad
Bf2dayUEwrzaixQeYakAGgMQbwYXq4dY9BdCHFIwZuyjUGKtQVFHH7HfVRyWmevW5KiNVBgdtYQD
aX89CN7H1f7Ae/08XUT9+HaMLGH0j9rMAsMPbfC1x1RfwGiMC/oBSqxycFY0w4LGh8+YFvlASvcA
oOSQ6RI44VXo4HhVZSLw/7t3EaCWnRHJBvyOlx6/ZFLfM15gkoAWgf9aKkUOI6uRqmqr+pyuv//l
hfsTdF4ND9d3UCt4wlGRiLfTxitc1TmmpOjkcq2iWMNtEUEq7qAGvoQ0Z2DsUFFwnQOmDM3iMkB0
ByHB/rBnkDGBwwqOXluJOzf4klOL+dJ+sGhohewjk1AZC/IhMm63DkFz4Jtr5h9b8KVVmzL6Lc4i
FJ3qEvRwiVRKFpgnrPQ9xGEgiHVaj/PwE1LcPWE3i7JR7FzncoiVFjWs5dagbGul8kqPh1TcpPdW
j7NYVhqJ2lAnnglsnrI7cIP2d27clrd6fnjtVXp5gp8IKf9XN9x8xFH5zaf6OwtbMN9XtH2uzSm/
S4eoQSQaqtUXsDxGrjuEbsHw/LS9CXOLZQXEw3lNUvVO71N99U3k7JT4zUIdxU85KIjVQdefZHK6
Jr3w3QC3ODYScZWA80kA0GJK7zR991VWsErdwZicqwAfwDPevhNLAPoTckGJDr0O/s8H1xQPXf6c
6XfrFRZcVuOPZltMOQZ9tjEaps47jASJq488uZdZofjErtYcER9Cl/zVmIMYGider5TyByBklzQ4
NF3IMY8Yzx8hfqpaB2d+OJ9Q1y/qWuyNGIKO/pi9PV08P1xtwj+UVn//gm4HjarxRBsWM0oGYdx7
/P+PXH/yrgG4h4Cez7VUhHTtUL1q12HSDNcgmQVpEcuCu3BdrCKfklQYeek1CBeV+QvKF1ZSB6k/
2jGUPS3YK5+TKyW/8bzvwh0EYW3dbsfN7QHkZoQvfg4XeqliVddy5ZyhI6Cu02W8Z0N6YK+i5XmL
p+MK+9ZgPpmWqGBReEvlvyB81WHABiIAnrD1eplsfL6ugXUY/6HA3SE0PZM16cjjR2J1nrd4RHMV
3kRIWlSxpRveRScHQ/XZvEyoWeexQQBHV8uT/m8P2bbF0Or40/wgx8//baC5vm1heyhngSlVmaPn
jidjprG3AfXr9UIwAXz14rGyYN3Ujea4cEi01EAYJxBPQwhSsLUQucS3lwO+VFvV1bTprfMIZ4Wn
IHp7jmt5dCu2qwn+cKGTgM7U/x77OjpUkCQR+ufc+RFMDpIt9+YwoDrCsq4WfgEuPjWShBFdkLnK
3/zr977SBbJy6UPxN2QJ0yvNVkkg562ZrSfCYsI6vmFFst5/mPGkKuL+hOTUdNPqhkQrZaUHNUpd
P49gpKA9vzuUJSArHshcT66MGo7Ke+ueTxn1riys0sEUUR/5xqxNvAtJwwkB9d9HVz/WtIFUJhcm
wxLrHp0FsuLipMD+mC2xuOygfnBUG/oTM5P9Z6VpIfc65ZdlQgj/fmr1RvgWh0WMJ2QQx8/VkSOE
5INf2kchea2AfcDoXp7InraaTLbLZjSwxum2fAUl1VMQfaIxhaZ+pbqif0QAZbLY8keH4rwmSkCP
sdI1BAITGZtNq9cdC/fnmSUU0aoBKa7Asie+uNwkV+gaKw90tzfTem4j3BwPqZcsgocW05CgoER3
TafkwewpSq4Tgnp3qXBymdYymL8thokq4quvMcvI12etVSYIpbclzYMlv3CrHfz7LPANgIUldZaX
Vxu0wf4NycmTQYzkXfYyT1nre9tsBocVJGw21OskkeeyD58OP75o6xuWBZYS8KFAxNVXfZervtDx
zgHipd+Tn/ALHm2UlgcV4RALYJkD/pKmE4A0KynUSe4GlfNsWidUjOBeplBM+3ErJOsS59SLIgMO
3PHXNl0wOmPtPUfGN/Rrp2dLWqFBsf8HUva5ut559QtjeaXNnR+5MR9eq7SmTPemCJXrLCxVT84n
zl9sRg46gB9Bp3l9XtSCEBY//GzFGWbWxJohsmrsD60eq9VcnyrgLMBd3fOLnYpamY5U1A4K95vG
sycZkpRLbqWpxq0M2AOMM2v/wLRSkWc8RxXYq7G45werG9APBNOxI8qdMzozwM3OieP/snR4ev/6
EtgfBKBK8RJKOg+UrryjmtJj7AeBSwT+o3H8kHllPGhXfHeBPv+3U/JldOvHYeejsxOPokZmS35z
Y+rWFWexrOcJu2P195xX7KAhbUXozpMC71nxi00IHlI593/7AcxxzRtaG654Sv+4krBqatvdCZOJ
VfJUj5eULTY2+lx10/v06WZ9yQ2AXNJWTE3WBWyCXq7JzFp19thrdeDVa18Dh3ewLMF/1O4AuT1T
4vQI4y6IC6Yg2GiwjkkSgIjAfxGz5+pKndFl/6w2FNU6bfdH1XNvdQqsObUWR4kKiueQ90Ah+8Yf
pn+QZ7wr9PWROrYY87klE+v+0RJAHR6TFWB4jpvCkfgGTBL8To4Mt06el0TDKJl9Ymw/7mvxtMMa
Zck/U8Gt3gjP4LgT1J37JQp2atV2HkWrD7oRbw54yMwPe/BcPN0IcyBwHK739/xu5lPzGmwNqbH0
Ln/n45c4iyA1hKOZxoe4du2hR528Auor+9oLZfYk4G7GW56Bu/1tZfFXSCi5CC4M8lAj4GMiRJnU
cXCW9EB9gWYhm65GQ60T1u7wL5czA+9jYdqMtjTQ99nISoAsNPyCBxuTx2gSn4sMSWI5Qtk1/GIU
hjq8RWReX5ExHxiyvKOOeqD5YATdWNTpHwKEQnwaj04c9a3nvGP5o8hdAfX5FicfTGFwsjtBfIuY
8hRlAGsmScTCDUkUtuooaLCAfQlp37etKENA3lRfsH6hdRf9DzcG1uWTetCbrNd8eeRV722IzGKD
NiN+3ZB6X+C0OkhI7t+/sVUZdufe5Ypn0h9eooBV1siwPIFF4t0+ACcBje0qrsv5/RqMD+92a5CF
T07ZDfVoVXZ/nITvQp2rXyr7NcBMh4dOlRrP2/K2dgkjo9U530kN+M1GJ5bpQF4HJbV1NqBG2aj7
sklJi1HNsjUG7MKuXqwcf00TDLu7acs85WjKuTe/JytNQlUPzxqCQPXPzYGpAMrG7bNf5gsJsFBC
zDCCiFK24sYHS/aPkwdklt7O7dSyz+dqrbH5kcNweM8GW8GhyqkJKrtlKYKnfEScUWpT4Ol6MYBN
Gm+3ep7pJOlXIaG+UuvWGROql3UGyxiko0cknMYGoFPbFVb6eZ9T9p2vwI3hBU7nm9IogeSHrath
ocrK6bWM+wy+wM3HVXdB7KC2luZoE4C5+acxvuwjYr6FozcfXLDd+wA57SsGtSYJKzMju3HRzk7n
jga3w45F4pFV0tcjo+5gYIB4kRvyZeJj4Q0O2Dzeh+ys39/zvBs2X7RzhhTJNNTECNDA/Veo9D3p
uIGG21hOE4P1H5TbNoJ0Y/U5C2QfDUOfYF0fMvFl6kZraNtyNGWelk7t74cHzyOXM7yYwGSczBxB
zJbLNdyOCVw+2ewRacl7+L1iqHCgiDITZrx77Q+V1lVHGPCfZUUud7NHyToG1XQywzFL7V0nMNGX
yEg1Kq0Rl2gYooB41r/RrC6h4Y6cQ8FEtbznNykLSDEvxUEW3OOuXbgaMJS3wL1hd4AS0ywisr5I
uO+JFqO1JMNNPVQXW6P5ofcUr7ustT0Pe+pnO40McZqWHxRHwlJ6UILXlu9657gPH9n+mHleTPOZ
6HZZF8f8JzWnbC//HnL8wGa6dPG41mBcKxkwxz2Wmu1SOGTiLs2lJfKKoGK9o720Oo2rLDMQACh2
F2OiBIT3h7eY8HNPJTEfvCnCcAjhzUSgbyrHxs9OI9hj/qa19KXZ0C50A2VBVeuxX0IexdqXc6aV
dvzpFz3Be1P3fNXatqtEGLM+9B7VlTrNx6uO4Ki2NsV/NjcSVz9QuMaip6ODCaT2gseGhiwTt061
68P8KGzD9J0DhLTtsgFs3CD4PhbFxJI/c2ZC8ha2+HLldMeRwsjF4L+XTC/5fcR+aZpdVKQq3X/G
mUZWbCUDh09iR9KS+2b1gceEFT/2EfHdxKxkZ5lmayM5PSxjXUnzuIBVeVbu9GCi2km+ZAMm1M5M
rEUYbX1cGL6nxVb6xhUpYlq+sgw8RFT4RTsz1x3JnEm1w9RSHCs80W8REtgYF3IxN6sHrgBKzU5v
/U6JMIsdaYAxcasepLc9rTw8NS6R3nZp61vIbK6lIGeZ59O7tI92cyIvEf9h1PBADoyeSTFjj8/M
9fE5iWM1s/ssP5e2Ysd32KGbp4pq9yIMRJYxcAn7Yf8uTJKHjr/nTUodtU8donR19ONbThWRZwiv
KSYY1KirJWeTaVC7x6NOupRdxF2jNFNK+wNdbYcSo6QJm8IyPugIdwxqA08mZTDTYEPFMejLA05C
YPPp62cYU2apNG4Gd3ulsiX7bBPsu2yIiDPltSlcRz1B04d3aJI/nTdra80BWvuMbqyXLtkVOVDy
6wvGBcedz5/tMnE3jZ0TpIMukgWDyjq2X82YjdsO2OWoU8mi/j1XZH0612ulJXBpxwEHLQRBG50U
yELz7EXgxMyoF9+NbJiFVYh47wAWWu28asvuN8uoBFU2G+D9BEyKDQucxOvOKpc3Knt7corkieQ5
wIYu/te7/xREhY/9IGYyQb9R0rLSJhuMBdGCU8+0ovbfyyvLMBpJdhHB6sKjBpzsr7F6LlhOsm3c
LtEglf1J8WvbQNdRIXkcJ8QQQuIa2K6U+iYjlcXsI4g5F9WbpiAV3WlTQWxNU0v7JCQr4IF42ALJ
z4kmNqx5vIsZDnCMSFfEgJdI1KFs1P7JTqFZoN8Mn8tcPjnRrxV0ExlbRycY5FUJBYSdofr4WdnJ
E/x9KnOxO0hzJLDq+NB3NAIGwWWFtNdUikcOpubYlPSA56AZf+/UNJ7YLyX02PqZtbGu4pr01Dfs
cynK7v9l30mjKUnWGslZFXcZV8k0hw7q9/YzCapCNTSvUU6+1XLNsTvEopPj1Pk46wr8n7/N/rYX
vZeFzKSZf8vbaGtN5HrLnZEyiyiZw/Bt5NSN0PD7sJE7QpFb0mhOMRkzUyRRQl4ZIkxWoHStiJOv
xrAga058bvg1kuY8uiApIQEZo11ioibZbKt1TtkE5Hf4/ZqyQYCXeH8rEdwFsmuGkAYHfuQGMGQp
tbvHmT5nRr1XLBR1rtcdERPiq09HxD4dfFvdgqek+WBiuk/LbBHjVirWJSEOa8fBH/jXDmxxl7HT
9X9IdebbL4jq5qgf4hAMiuzorce5CybsvRg/9rw8yFQSClar0iVysdIzdsKWUfMMfhTjiUbPN6je
BooRvnvOh7fB7oL6hKUIV49tM73oL0FLuFUNPiNF7+wyETH8JgnERN4g1JdhkIGq/WqcAo8YMOC8
a/Y4FOHya1IIp0x014yYuieVwx7Ttm0V+Da8cvDG/6+t1N1lrexOMZi8RFQnOUfbByRtIBM/hKh0
PVmw2HDjVTRJsWaixvu4KKFyFoim44BZKEymClHS7apyJPMjI9hsS8zH66DhNSQ1dnOLypexIpkp
MDA7JwsNHh6ADsYQi4i84Z1EOJHFD+hnM4MYlSnvBIc+bG20eFzqI0mdDe32r11dVHTa9XxsaNoH
x2wwEC2cuZkqUkWHqwZ6itGQxdnRwziTsVrXU5yoZiBMHR8fRarPTwVvLtC2lQ/WZldcuAufdmGH
JVHPKxOsnyNlaV4xBiZZ3wM4RyMDY7hfOtDXaLi12RAg0ILWZknALQiTPXJ20rGuBJEFhB+C1e69
/2GC4hXCEUjIALvCY7zG9phNamtotn0GwIuQ7ME3ywu5RB5axnEoTmb3k4uhyW79fjrYTzrYwyYj
fJfMfcIQtvlLvtsVoGF3dHdIdudeKb8+gYB59dr6UWJRDZp2mePAJnEQrVbto3dX07gyPAOOrvvP
e5o7Xht75IYhU+lqXDtTxmK8uuwqnO6b8k5AxZy6clU7jHnLHTCi946ClSBOoDta9kO9NWtA8NGD
nI4DHwHnGP+ukJRh04FdCs2Czzh21VrDMdi9r79AvXBm1rucNiILhVNFanlRpA4R70oF7aOnurR7
BNp8lPei1uEVhdGTdGGvBI6ewW5P0B/aMrAyLx4IPVYMoVPAun5ZcBHLMw/QyNI7iD788NAU0Cit
b9qganaCQCdc9w2c1iAZmP58KFt7RUrMg1LMB9IcbRFkbvWxC/j9e3/0l8xFw2NSIc6qgTHa0Qtt
ppBNFtAhOfDyH17S303ol7j7SycFjg+BlWWLIOeYroC09h/k88QW+xP0JXYH9zqiKIeN/khZTYvT
4cBY+AsPb7wzOx8YrNhi6qsGnARfwAI/QlQnv0UmX8Nuq6RxW8siwK9gnorcyqq7/Bz2l2l6YLzX
AXbP/olFxx5B9pccBqQqGtlSHl8A3yDnpRa2HqacUpE2ED0lq9vmNKJbyW6aP3Sc3xUB3U7QfWnP
CWFVIpS/o6+KWnFqaE9CjoBEQFDnYqmDh3yaMzCc7ZDHgqpDpCqH0hgXambJbAlxvRZ2FtHMvEo/
Mgwd2f4PyFnOu42He3FGSsPJGee+ROidh4wx/iN87vkPrZMuLROmqMXVy4zlkVxtJoJUPiIj2z1y
Qw6trO88ItJ0oMx8SZjQgVkufVVWJW/8biymmu0PL3oK/0R3EaeVYboJ9COujVlZZrU8Cy7A/vFi
Y04H1gfOsNqrzurkEV5l/QtOo5cJwsi2kzwK1qjXWr9B8jFmUdlB+pvYy0VrIzdmIK/b/dWB6qp+
ua8Z4uDGK+p2uK1FyXSrUndHFuqtUnx+SMWHZunIDYwQO/bKwkWfjmjAGvoqHGgn5OL/N6/QBFP9
FnA3WwHWnhky3QjfSEvkNk6BgzNIqiqGU3REXLvZen7phEOExqD5gS6vJXlqcyfZ8ZugThEyw7c2
gv96kxF1n2lqSyDI64f41ennY9bIDrlclFup+tvV3gdSHoGl2bFvTZSMNINulDL+j1pUpw8uKVIu
cSWx5f1hDvTe6ZA+VyFz1s6Tsgb5ZQLTINa3cHgW3EgrN2HCQ72XP3ApQuE0JKPtcKHis+fhYl+O
ZX4GoXrA/QwNDrmHlwN8RRoPqp+1CByhh3adHtevp9rhXbdxJVs2yv+EbEV18Y8mwDfm0Z+T0+eb
Mt5vJ4Act7u5cMm27LFpx6Auz8GYuKntvo4x3Wmytb4RbLrOsghCUtIDHC5sD9QMhgiMY93dx2Bc
pVfrGcxZfw9Jx/TRn/UXgfAqwz4BQ6hgMmzysmPYBIkHRZ4AefZtOduy9iPT+Xb0HmgrHuE/tWE4
5es7t6Va9J7e0MD6j+ZYEbxY0eeUYnQN7gVf2RYpY9ZERdQZitysTW13t9Ptu/4ABOO8VQlVy0Fa
L/ArA5ccIb+FS2IShltF1V9GFf+ilgLQhPAMCV7QFvmJjEifCXcBF52SLZHqpccRLrY5BE8ivyiW
UhbTTLbuvFbo8C/dVRwh3l0/Ui16KwgnBMLZ1F0xD6bVMKsXD9JyYEGzTrtczN7LVWIIcXK2zS8v
1xpW7tl5hnjfMpXscjm7+HtDgx+1VTDYCCC+3gd3P0HmKOHqGAtzs36JEhQXCFAektuPPY2nR1ud
UORQ8FNpFcq8hePNtP2hU6r040Bush2WacKeHnIgiDbK6TEMyZGfByU8JcJGp0F0D4PVf1RNStUE
XiKkdPOEzq5R9m6+jQdTY1IckuwDtOw7K19KzJ/UxrOSWN/ORRqPJouAqa9M9UFk89P/b8Hyb968
q2QZq0hGzQQImpUtaMCulLFv5T7sYRRz7Y53S/02wLrhsAYmSm41rgxwgZD8FBYXFkt5Mg1Jrk0l
LjHtmyXAzx6lu5uLlcvJnvvI4w/pXSjVJVidNAIJ0/KjALU+vr0yYLc5ocptaeZHPkEBjuJFv/LM
a93WMxQEbsk8dCP/Hu4A5TsBCsDFma5Ap++YQXcFgu9rZBqg//zYzlbCCypb6jWPo8uoRHtbTAe8
0E+hr1jiKPBh35YSZgRyZoMfyLpR/3REbd8wc4yaIdazygzoQMXR1oE2nPxAqrRyUwLv77cZhjP/
hSnU8E/CeY2CHAPoUhUnrIRm70PUhMJxIg1jzCGqj9OGrR3Fcc58yS4wbpxu7fa7tfuyYCopwj2g
IcG2S5A2FN54gi0aAuR1lxQzCH2eW2B8tAblh2xCd9Hd5YZf6jbE3fTxUZzKJ5sK5VgubA0/YJ6R
3FNhHPwewZ045OY65pLd/tFkeKNBZLFPtDm1IaI3dHiYVdYI15aTlHsa53oWuL1xQz+Nm0rAPWje
byEv9OZBEdXcfhjnscJIblIBlNJI+xGhrgGxFTzxvElgWDV/mW4zUufPztdrqHaItuO617XFBjKl
wMBscAir5YDA1ZIBJoxlBfs73prG/hQa+dHXf4jax6o1SmOEgLzp9PQVsN4GlOA9x5wRCzTFZhYM
k/uj8ZocNVliOSJZxRjAxKtbSjueJUTdsoR2qSfSJp/9HfQnW6VNNXzC9xf9tURkBXCuXqweqa9A
cQ6IY6qQrMZBvTtMypld70YHq2/5bx9i13rZ1cWm/OnWmpV1hy13gTyn/ANJmFw8034GlzXilH+D
mE5ht1Btbw4649rr0kkNMrr2q2MfGDTJPSXHPwHzVXc0utUHzHxEIimuPB4enskHfc7HlI06he9i
ObJSIiUCKn+qpCVVtTW5a3so2olb/EaQ6OmzQgqjUPLKstG8/7BGeRR3j5nDy1xxfSqVO4AJDu6P
hlJE+nRsmlYztNxUbuFl6HDdIgP/t5fnmkTKNZ5Z37ITrsWt5JJ6i8rj0WxMUodeyq+KRW73/0t2
vf7+yXjj3l9Va+0cpVDBriBFiwTkU7VyMaS+UFK5pkcfryrDtVykWfSt1B1BUjLVaI7ReUQk8l6q
XZr7T1JQYCh34zh6l9lGOyj4pnAnNOjyFEeIhSbh39ACVFa3c8/LAD2tTPPTmXCiGtiokzWFvt1M
7nXo564gGEH0yxDcHTjZMaYFuzstFkgbkkX5N3k6dI5SA8ljt2/9akh3fwEkkBx3U3BddvSHbbwm
G8YK5tvzSDG0loAGZ5tu4ts2VuxpxAMfWNgCGgvSmXGaH8fJJ/XUyHZmdguLRRTGgmv0LsLKuIjR
4zx+tD4rDROyth2KP9SOujuUI8GtpndXTCD4MhODNNlXR8RgDcAhRHcGavAWN1tOjEfY8L9m8SBM
MMKRvKDO/l2nUG2pZG8uHeRX/vy2lAND+wP8KrFP6sX7m5YBjHZ+nWwcsXLkOYjmGyPStfoqX0Sy
Oh9Fe+o9KANbI2y2qeUZr23+ZFT5YRL+sIB93IcMI6vBhiN2n3aajY5jv7Zsoiq8YDWXq2VYyx/W
TB8HFhhzGhD4vYghPwq9zEmzTI9g3MfRz7t8JSDkQB5nUrpMIykPyuQh0+D5UfNS2/gbvJVGJngY
bHAEUsgoETCaRlnHUgJiEGU8Uv0e96OTNJtPGakDCbnnHlyYR0teF9eZjmk72cqhFBDiRIuqefpY
mfDB7vRKbvIOMEIYF264EBMDfj8bPAlv0/VsXxGZTUnb2ZizAbdj+naa89hGNOMGYDvL3Luvkdyz
und8B8yKgt4Ll/drLB8B8VYlwICOM3xGabA2M0emiB4ryWJqIj1FQBMGoqrP5ChsQ8NapcJ0kTJC
iGM40Tsni72Na0/MxxRTJmN/I5K88x0ywHcl5Ak+AL+2Q45SZauvX3CHa7Su/s/qLCuJqx0Xxvf9
Nnuo/Pp8LSMcknIhggBsx9JyK9FumIhtFO+ogHHEwEect/c14R5pzChoUZPH/pGGWYYnqit6O2lI
6FWeyVQcrBYiyS1r1Km33UGQ/FQxrW4z3xMNTnxO5Zm/ni7NnDVDDH7SQsyYUrt2HyR3Q8fGwP0o
MPzK8G+wzMe6+kQfSvxgMTUdjQXAg/OwVn6Gwu/6RQvwa5pAfB9IDGSJs14bD9QIW5qt8bErvygy
gypH8/5eplkcCyq5z+5dezVkQIwXvT6P+amHtg+4tWkxQIL0n0yZUDq4jo7lWq8dNml7f2zeaaQS
BTiYytNltw1J/wzo9FjGCo2UC9PF14YryUAM2S/Zb6N5sO7h26p7zcsrL6U4B4/tWXMSw9Gik7Sj
0mTxo7Csf8Al9pIW/GIFs49dThXUK1p1HXbLQjmaaIeiPBxbvlU45a0AowTAZt3JeZHUknbY+cC2
0e6OwxCQuGc2T1S+2b4/Au7hNiRQwk3YTyGzhXeUJ7c5P+/xBC8FMGSGSfAlQVUqNB5o7IojjU4X
9XA/XaaTBh086O69JC7GkU6c48hIzx/bALeqD5Wjvm/RMwhSfHQzj6Znb9QMKbTym6c+8c2h/QtF
XjJJVC7HJuG6wdoEKIkKV66imSWPt5mvJoDTdoZOjUOmbNL/u3DQ1HxVrvyGZIEhjh6hTYg8owC9
Htj5gi2kv8xZ5yrd0eyU/co2q5nU/OUf1l5rq3owUprWem3knbWoDFtmGdMX8Eo0cvDe4wG43TiA
Zo15ME7I7sa8hT5+d63GM/mEQv/boFy2hk1lZZd7Wy6Au/kfYVS8rPw1AVhkzFlA3nCSi1Cz03Zs
l0Xq2eAVhEfZ4YLincki/hN0L7bXJI83XZk7YtaD22OurdHboZmPfIhvHcnrbQ261SFergNM7DkJ
C05N1FoW2B87DH400tNiyMKHj1jIRGHw+vB5z9pcUGc0gkwQo6xq7BTB7/FTs4WeXPgLyVOEylc6
A+Njdp5rdbTcbbl4LB7AsYeQdDAVIgwgtH83Q1UylEd0aG6hoHhOu26HfdgBpiQCPxK67rHkyJYh
H5UQDEeQTezfPIPCtMClJQXS+q23zfmDaPbXwbjr5SeTXCA+439YLTUVnVFH3840IAwf9rTs9Ehj
cqSqtzESL2hpHnDIGI+TaIssKUmyOUC52IB6eglBd6wzWg6VOTSvhZ8sbI6HgYbccm+2PBTdY+1l
be1SRPcWELtVg+71kCGXrnUNKDq74Oc88qmvdbViYqHIaPewEeUdppmMY6aPicDflU/p2LC0LvqY
+oVM8HvVwT5UePk1gUx/g78QRGCL3EfwANtEwK6Nu1IG2xuNayB4loFt0IkgXDFxDmTMm6mKNpAl
d2EssK3UPGz3LvuIJZVIC7MISbXVy+YRhW6pQx8Z9ITuU6AwhKCxcgxUhhs+nbXNeYFJXyUFq/5X
w082fCCmPZNr7z625GFz6yWmXib0M0zeea/vMlrXBM5x0Ca4RNjP6C5C1s7ld0bPqlw7Fk78yeky
kTbodcSZ0ILJvYQxclFwuu4cQPnJtNNakPi1RkBsws7tYI1+zAGpGpyGhZwX/ioMyn8LkdwuLYeF
HVrrkQ+ZnoxHV38Tn3KJ/18G1dW/3jjA+q8qwJTFWKFME98yvxlWGWs0kq2fTWqdDSnvbt/OP8Bq
6JWFUgXu5xxiGc+QXjWU7/WhEi1Ro7RvTqYziiGmNKD8rH2lbt2+EmBU4pw1t+ZUQns6pNTvJGw2
fa42gG2HrtyEtmJJsC6m8SQzWWy695n6jWiJOaqZZMbI6dwpk+7a08bGu8tQzoEI2SWXffPzbOjK
VPBRlKIdxAhDsiOvOsWixzipRPJ0XrQ6BnGiqziEHQKg1DhjtICatp2VTnv6zIZvMuPV8AQBcvxV
5quK8AJR70clOhqdX4RfsrdPGsxp5+uXVVjzkaOo3lKEwXymqKz5SRuXnXrov/GhkERngJqo635d
0JDxx9ihCJrznShYiPlrvLlDPHGJEImLEDFT/bhsW6t6Ge7qYHU57/e88rUJ23WieLLXFktm/UhI
JwMJ8+iIPDBDR2pBfymavWvxQvc76gc0zEVFifTPofkTqysFUn3p7S0r5o18LKjP4i3laSZs4RSO
IraWh3CM66SmVev+v02iDlVJwevIvoWsfv3ezdjzePLtLD36zsPs108yXZI4Q2Zf5Xq91lE/M5iv
VAwt1UUaUOqGE6kck5QO7padtg4PRD1KoMlsAPBRlk52dD4l883y1mB6I1iWkGRSIeVPi1x4fIFJ
oVhtBaHr0e9ZfQNcREFN8CUq39mxPEv6VSAyXr29zhyjwvRSi86M50+ohzrD1Rm9gVSveF1vc7VN
XmIwzzSUe+L4uv9ih9wbNMHJtVsVloNe5TxnAlQsE6QCG8MDHDQLPpACGqxcn9TY8UKGdGqfervt
PTRatZKpxp546aHXVbtlvTCoBgaomPbaFfN4a25CFk+hJyvrHwNF6IBzf2OBbbagwCTopF6OJENU
JJxNn5vhjRQG4xKmMfusTYW3zVI7Ukm/ji2jz3fFOKwfyD2wUyPxS2kgvo4pPfxIN8DnXQu22rjB
0Rqr+RUWrCadfP7xCOCPMUsm1cX/02AO+AXqH5zL6Xx2UlFgvomsyc3rvllP/4i6qmW1mfOLL83X
EBmv008qa9cBQRbpumu/ByeiOou4Fl5TCCF9Ra2gWkYUd+hoMWqSa/oPgk+g/x1lr/ISJQdYaGe9
WQIboMbZKUFMw2B3KCBNT06L7GHCiLdeMqpW/aS372/Ccf9EnAvzm4LbxGG4usZ59kzgTeD0VIic
6OvbQA8ws3XrLBRmGthDUDGadXiaOAFbwl8PVr73cZwiCXslwsvFiZ/THVG8Mxq+vynkQ/Vsa+gg
nCDvAjKm1iQ1NxXSGgCJ1223p3KE0EE2vO5Mu/q1bKw2AexUs8ELauvfByW5hoM/Rl+W0irI7uta
7p9Sk5rf/aHxKITet/d0WIU3bQr30AJN4pv7DdaVaY4N4IA8nPhzIv0CAoEUMd94DjS0mbNQB36D
6eegbxff0JNM0dUYtMM1S14VHxVHZ4pQk/2NcWB7yYt25S1qzZGGimRcX+bT398lQZBhtIJIgaiT
tBH6vs2FjU0O4T+3mexlO67wJCsopTJG29lu3+xjXQZ+2jQuXnaWu8W1TDjiOq8vKlFae+RxUlS/
kKUxrxkmTfHrwRFChvNL6iKmUGOqxctJhy0mTa8KzvLkcJXjTZV9MAtVX3Vk1S4tbQv3uYUy4TAb
D27vmlG8j9FOBm0SzaSFdA8U4xwT3vwUFLUkNqdZyCLEozkuv6kLDgA7gZKYOsUkOOZpTFLt4mEU
HDpoH887iiQ8n/u/NhwFgm3e7N7KI4MkGv4WkXjilW5xEBLU/MlpuDKJuTlEE842aOGZx2VPMSyu
zSr7T0nxrmlxRki/EebL95cAkI5MhJtvKI8itjWpClwJgRv6dfE6qYtSt6Kcqtwg2ge+YoWb3Z6E
cCmQDVW7tf8kzAuh3Rfb9bTLDPShUg9MD0Wc9ToNWK4ZZoTlo3KWu6bh7pMWR0lrnF4Jm0IOFM8C
WKXQpfPKME5RYDSZmILYXCbtSLRMYhvQRUDqTXEI1F7sX7hCA0mz7mOxfJBT4leeXN56tvlZhX0I
wT1x5VfdKny3RsLMkKNwxnskDwj0rf/jGmHlWCe7ZdA1wDB0QqY46ORxF+ceckMXz8KG7TaiLwMR
FpxIxKPPPoNYq7M8eI0lpsha0xtq3TSbtdc18OhFzOh6eKCgs4+P8CMwdx1DcUQwRuEZfaRr1cpc
mZTUqIl+DM3bpI/QMVtItL3E/UDKhQGHTcD8Z9oAWcRuOLC7/CQJnAer+vgKaYFpSOiXCobIraVt
MMS4m6zTuF1//bDepTyd/qpWfVaAoO78zx0jHezikB94J0Pd+mH4AsS1vRkhHUgfnBaw8CAVVF0v
iLNPO2wnO1Q08txYGGGqEFqT9qeEjF1jt8vDe8D1E70ihFe4/dZumKyhiDqnlmpS4tKHs6uahCRb
FqTr4ei1SAyCuWPwxlgrD6sWmpA4ByBSw7IWuGnK8CpoYYk8UASvlu/3RQkfJX+A/fnwOAk2KWCm
wQ7zzfQ/J/R38c4JQwoIMs2JaJEJOWbqnx3FcRp0bksdaPuLunAdjGY/xjQSy+4TxxiGhfLG7oH2
ycIdtRNiTXTsqz968gD7J6gAcE871PCsEIuu1fRHAdamqMEI8nYh83Fz4n9ffXN4g8/4+fJ+WR/x
IecBPPQP+XFntNGv8ypbPzmYmuH5DcA1mqC1hmv+g+3LMqMqTmHmS0jjL6nkCRzQR3XHuCHu2vIM
yrHjECXLMr51gUvbyhh5YgoL7pgWXuV+Z1u7bGSX1Fl6/lenILBlyduUiOOF2321IXV14V6uT7QQ
qLYJjTIeG7N6DAHcEBls0w1qjHgFgHVhjGzk2iv129krUYNjl4nf07iuvhI3JYQKx1wJoz+zI98/
KszHPL1vPvuoL3rpQq4GuGijWy5hHX9ydnErGB/nr/BF1iI9hUsxA5vPn518ujVVVlNCEhfFDFyp
5xB4eRfSX7vwq17bd4SMtXzaBO+bCDR0bmdURX7Jm3dT9rKsf44HXLr//Iz0PGiVachJcABArTpW
QONPJn5XbsWO/VDg4D/62j7FKV32+PgMEv/qQwscM+fZRbISfKye/Zp2+MmR4fipOvcJFpOwmqTu
80eGxroJjY13JpOWJyM9kp7HMcbBHJBVj7pY7baXf5ep4Xdl5fejysW+9eNdkPaz+COH8J9Mgr+2
uUXqG0mjx2r0lOMW/tBekhs9nw1loNt43H1P18kob67QUky7ZNN/vJ3zEv1GA6z67z/F1PcF3X0l
dnaWPkp+Nimmig8OhWkENdQgw/k9In8Lk+EpmAxVZVAlwmiZlysHF3Dzv0cU9ne1wxrl3SeRhx6i
u1KAHWYsTPMDre9m8vVNyuUoNi44tXGfAd+CoIJp6UoEMiRUbx0LVE90gHMCOVV5CEEpGsbsYHOP
J93AxO67yEY4IYSBHc+N9wdxuuDUYHZYWb7hDPt7/BEgY9Gy8td1Jeop3XLyEInIrzrKXsHGXEiv
OreHFNsK6BiPV4CSu6W1bSlv7RX4LFYYsty0CYkTe7mzDE+QO9GoYKP9Xp+j4oZ0ljXz5NMu69lD
yRckplw2ZrxVivMCq5In7PmzyapXnShR7Vt0Ctirwy/ODV+WQu7EtGbXWZyMHfBjyAZ59jhn7/w2
8vCbxNtgbL9lqUzKFfxKejPWvCIjQbimYXH0BG5MMifdG8h9rJdLdGbJDkBJHRQ9D2eTSrrwmfjK
mFVYYSMo1TgMaVkUh5hD1K+H7+MgV5m/g4MhJKIkRkjB+vJtwy4aPpChZef6vLCzaArAoJp8oubm
aKT6uHgBwfYNXTPeevh0uFAE2V1zROpy425F2wdXaLfA3lSKiiZvU1u8/Bx5Tzb3JE/J9s/09RKe
vFFRDNF8BCJ2YKrCnH0/ygb/x2VXndg/X5vI62zMpSAe8TSRUD2Dz+mutvnkvzczxKGeLbl9VHNr
jP6uEHm9WqB/omta4INk3je9EKUDssrKXK6orqOtySavOeOTkcpacG9Mr9RtIeyZvCBA9ltqBP5A
2K5JEnTGtHLP4F7TekuZboIGmb9sg37Q+4I+8U4h3CtvkD8gNJUJMS1Eg+0XxFZAWHgL8U/8SpYl
mWU0uYSP8FVGqrPKDLj8LuSBW+HPYLxJfw5IftR3zarFFV63spcid9gIwG/olo16UCQuz0HCU2nR
epQ2iU4oyget7hVwQwVyA4oMXw+YQqRXyNJ4sHmto//CAQtajr35r2NcO3lGPT9VclwiMNIzp45r
smGXMm8+HSeVy69xwNxG6SMlRs1+Q+RevkL2feo/GPt9RdiMhrCU0rKhOZEg/dIrJQ/GQldUKyrX
be01FlAyDK4QOA0wYex9cCqnUKKE1i7iXNe780Nk/NZ3mmLOCt07CsxeZRdT1F9LCmwrzuh3YKw8
czQHKtrMLitk+GAZkb+64TgQJix5LG+p7v9nLkAGJhkF8C+IrTLYkKzgyCFs28vJSzJrQ7G+UarK
w8nzXQ2PlAcaJCTQzw7iAd3IvZfMpJp6BzLvqmyWD16wBC9QtckKSzK1dpBI0YtjwbPdQRBK08qN
g4Xz9o+2sIudXueJHBjv8XN4My5yGUswrPz3WhHHBVqN83QprYIeiub2H9mKkdaMxNMo8UAd6cBB
37/i+WwnCtUjpaWHe03i3Mydkt2hHV8E6IOxbukTaTIw5v9MtXqICz+m/lVLLd1GMX0VonZ1Ytx9
6MdL8V/szG8zq3eTW4pknbwLljDWjaqWHpNG7+sLNw0N4mr7yfMWJ2xM0FXW7nWg+Y3dxTCDCsiH
DpcgCAe+14b2dT3XrnB7Q1Ylq7TBXhi9M6YcJrm6YkxN/mRIua9MtCpYr2Igu1u4eS6fvSpUVdh9
uUBVssRvr26i1IZtJPx58DcCVuc3b9GauL4/zRY8gSWvGcsR25H3hzzMtOontzzYiUXxYuEjtA8T
iLx9wwAX5RVpU+26vEkldHqPdpmKsUkiQ9KqBUo1QgRtkR2LBPJu7K3LPo21f/TS6+mBYzIkvJwX
8wt6jxNCa9Sw0cG9aHKkVk6WQRGzatscT506PfD7Hk21LMNGhFocqHs0EvQDA2laF4Pjg13nuNG9
P2AWQMWw8BDtFJS4LbeQhsEwuDNQecERiDYp5LzdqXHvSEsvgIERw0xiDNffLS/E7VYs5rvLZZcn
5zJtToqjbg5tUNeFjPZVyG+IcrNuuLFBfy90yZQjVA38rHLUmVMUEjfVi7VdWC3+S9ntC3hmVCS/
dADcrVpVjUD5om7VYjtf8UgR0XVUb9/G9BtKKm8ApKvyrZkb0eRs+Zu6NUL05texSdz/Drz/Z1/9
+BgcgusFbko4jNXB8UL6YKMn7q6WwddT+fpm8k/ll4y0imVtbs/VW9w1u0ywE+/YldV0dWvS1+pl
yUoiElVb+gY7lQ38NlvdAScYtY1MQd5o2p9QRmJBMPhqprDNmSW6gAozF7n640MVbBFGvGw0lXHx
UdpKxcEnhvZ1uNjHrndOVUVykx4tIOPQ2fFl0wHKs53Bq9HbeIgfCyHo695MJvAPmWJVUXh6/h9N
mub5V9ee7b9+NAxd+ewlZ0xZK9PzyPuHyClc5JVejte1qhusRP1zxfDXE7ZELvlJTFRE7wLQBa89
QtKg4lk6p/jnEkoroUBA4WH01k+b4/oovmjEeQT4O0pvMlsWPkuwwb5iyyrWo5e6MOQAaaHlBdFC
31aCraiOJPP5mpjRhcMfIHQ+v03+XJ0nxYjQPbA00sswnZjM3StUkkBnnLPQHk7sfYE3E5JCWrR3
Xs9ZdDN9tzO2xeqFpWFlARD3fIzJHP7MTFI43OJHAWmXiPPlMVwl5ephPf2dsNAYpmzWxlOYfVV1
+pRIQjOJNpLDm5I6le8oW6x9EykfjPOZLKj9GYgKbtVUA8EJ5JfRFz35DX1Ln1hpsyQHDyZgu691
g354Y8mv0hRDmfreilJofSVjZlLMoVUT/nQp9w4UCb24oMfm7HiUdP4DxtyNxUsfRUE025jKLEe7
wyfK58Pf5UFJ+OGpDQSPYe5D0hBmi3KM3wJM/yu65/NheP9KDqhsvRDLIxBmHxROgmBUB1kiRgef
wd1KG3jEJMr6cDCUu/2fGhORtpiWb1Mi9nrJKuyhLCOcjeHh33+wgfmjwzQmrKVBuAVSWsw8+bKT
BMssdHHFjmoudg8mZNXTzFPK9zViRkchQw8aW0JTyWuC9W6P0UBjOEt3oC6lLHMPOyvraqLhT7KY
wTdxAhUiO4cjjW8c0yOMUknk6YksMoVukZpMr6rnJGSu+knpK7g752dOjjpKlzFexa0rkHRIKmb5
vaBdfkIqHce3Yh4Yuzrbgrahhjo9j6MOKifDPa3z2oFjWMpIZCwb8B9pS6oFqy8z15HeyN1sS9Qd
ydtGSqxRTO4ClxOZX9CR0mmZJM4qdrhRqtpGYZf7OSDa03TwoqmJgQYg8SiQawDTgo1DJ8K8dnqP
kD4xFa8jN+kS7MhaSqqh7DZ0FLtur8m9XJ6ZPNe0H4yA96Frq0J6iUxPOB3fwA/Pf2K4w+qAaDAH
gzmMKrWQ+zYWmuEKFjGg6SSQ73v0+z2FFB26znu8R44EalNhXbKKQqV4gNOjOmfzFGjtkJSxL+tG
Ffj7FoSBB0O0pckE3PpsQh2Rn7dqsLZzouFz0W89WOnAHzGanWNenvaSUaSnoKOBWsR39TUcYzSf
Hxz+VAdtOD9Y4m/nfryZL6gx7fw4lkY23eBj3Y8eggUf02mtWHoQAOVwATFnpbdO7UmZiMMmZTL/
daQvnNSR/G33QwvLOTJhPA0uWr65nMaUEUopEqbPI+HpJMaYBGIaPBGXM57tPtmBZvCWiTfV0Oie
lixalmw8+oryXECEwz0QWBSKuTOi2a7OnRG43pMPzEaYECk2+RzDFRBXjUvStlvAtNi0ldenaXeL
eu0BY4OtsdCok7JpRf8YR9N8T3gccBJcWE0sJLyJOo9NXPjBRBNlejKSGixwi63cfcxAPkszoqiv
psUXfoSA76NiqK15HZcbwnvGCfaoScmF0fu42rX4CrGMQMvdWdHdPz8COB/Qp8im7v0JvFlNUP+a
lagTKDKa9biz05NwTLxwQz3fHBaDZtgLM5DjCPgpUY4zeGou8Jt+S/og0+9Ljq3VFBSYmt0au+Na
QLXVgqBAqikVjZiedxC0jzvwuRc47P6tL5l38XSsBO+z+Q/E2zcyh9YJ3IZnM25OgkyaJdVxrDpg
tHIgwd7UkLzMTM5mhuJWXFuY3z4aOEtyYB2YAsiJMZvv7f91jH8dDsVdrCpyPZrv1msyJub1OLCs
5Z0LEYXWCORMuTY48JTOUF4Nh8h4j8QHvGi1ZN1G0dMOZOgol+xuz2rl21Gdse956Rwz0Rwir7ZJ
id17rCabBmGfyp6RrnxNUmmJuNFuiT0Ik5xgFzGlUegU5LvJzFgGwODJcLEx1cYop83LbHvUwCju
VQVg0Xg+OurS9gbZ2K/I9ThzT7s64mCs57t+QWPOjKqWRGjMW88WHaXk5eqMnpHpIkQmO8i6S2G2
wh4rAAlStxM8KLseuJgPD+EwSkwtvx0/MWUfAQP6XN76HiRCs3AyQGp9mhwPpISmRhYne7bn8HiX
KiwmKeOkGqX26AIdOBIAIxi4VoS2ReY32TE6CzJBT1eH9hGFcZnD+CR1+AGseemNC5AUPxEgDoPC
HNh1cFfKrgxmM3tVvDs/0XjN1U1ldO4JwK8dpzuXsZ+5l/5lwTxzv/Fp602QJyikSrdZfLw+IXRA
0Kxk7eWR7AG0/k9uReBr0J08FFc7hmwGkEtBXhV04HRaTtZAD9d0Vss2QwkYi2lNBwRInLmDoBAK
Dwoif7eF/u27kYWHHyKy9vISHZvh3qLHxFXOLwYfVPLL1o7q/qADdipjjGEPlZW2LrfLSNifKiPg
C6quOl42DCKR/1V4jm3RVI6iDVN7Ap8+1jz/rUugw7O8+75FufrgP2w3YDJKRXzDRrYHvVEqHDys
86v7KnAp5qVt1G5Nij8BFR7P/l0YoZ18+AH81rrlhnPv7Wb9cOodtSL+7ORTpbp3NNVwPQMto/OD
7pgz2EO1qpGFirJiR3Obs+49emL6hP2ibQitVvQI7kKg/Zlrg/a5FJ2us1eAQkpHh0JPbt/5SHrn
QYjmOAOOndQx9zZHgohYY0eSBTuEMIRLuqfAHA7CJK+n+h1BwquCtDehrV2ZnZkaYCp9cp+0nO7y
FJNKVBuGXLGl/sSa/PhLVCknemC3ae1b/5eE2XGEhQIRhfrb/i9XqRXpNKLjp0NlSjMFsXqRjnpo
Xs8R3Mh6HSjqh4n8/J3UV1QjfXPCL97rKbea/5R7zuzhRJ0bU5QKGfb/Eo1zaKrQq/MFoLJ+21N+
2gdlKO01zfXraGLf2YtEPTILnQ3xk1MwmJFbcUHR8MrWrEcjfJ8YcyuUWzhiN8yPvtOF9uBDbbCF
SMDbx8p39uAus8HZlLH+CvKRcrLje6eAk5t5BlX5G4hSJYUFFCEQGpPV9JHQ2tedrHSkSoFZSPe3
44KJB3anYn6xSEB1YxQOiCn4/Fj3y6GRwbJhDMT2z10zHlH5DWlcqYRXGQ6naO2KQe+4ns7hIa2V
uU8m9TedoWhJhmY334BOUiOqdKwFJ0efFYFYS0yOT4BJMwXtnWIfs/84y5ibBpdp+5U8G1w2r3Dq
JeNQMsn/UhOvAVADPgJjaHhJlfXl/hH6LgV5KmcZD3D8VvFABssyZbi+a4rtxZGZbrUUp6TnN/Xc
4I+WbEqB/9DpyDE1tnS1Wp1CqF+LLFBrTZC/Cz0GUSPDFRMmHMoP3+KGBjskJ7Fsp2dA6yv0nlkB
+YVnr6fPw1RMqds+3z8eUyBpfLRZOKWGRzAltkxldZrAjISHtOeaKcUiY2q6FhTLiG9SK/0K7qaR
UK/qdvLX+RcP4daObYhcWILwv8ikn0uAWeZFo4awpUygDzzvdqJf70iaRrx6WNvv4EOQTYYxuuzh
Dur5oWRM1KyB7/evjOiid7Z9/8ad5/qpSeNYrDTbZMaq/DmSeT+C2SxSHz/cWcm/bYDIQAGTICVq
WoEc2D2ToYZBvEQOIWzVaOai14bnxXuOE/pen5aKuhK9CUTNK4fN4xx5rlMGK+a+6DdbxTqgpzRz
j8/S3mZ7PLHCwYokMkr5qj15oituawtk5cWQqH/W2+wbwmztmDn1Lz8yG4dfjrfe7u/iXsxXaXAN
pW/JqlPaOLyVbLiwENDe8VBOZjhGxaVoLJGrYYU89Az3YqGkENaQGY19rip9HYLUTIq87UvZrQ72
neOTKfrEYm3TkIUG4El3BpUYzYMfhKh2BYuWviDhYB8H9DygBLI9bn1htjgVgjIuUTWUB/z7a45U
ilcTRb5235WYviy/akDv/Ul0rGg/8ZV7tgKb6M3Kp97XR30p1ohImvekfAJFsw+0wK+lpv8i+mTV
5qq6UKWfWyaUr000qsKmuJ7SWnvKKFIy2AnSbYimDbkya9ZQoLCN7OkyHA/dgdQxpSy0cdIPOQTV
FORl8fOpkZVzgMoaDPUXnz6m2xxpMBhgvXKPyc/RccPL7E3MKv8LUQZO8avqw74npwLyqipsKluS
cVV3VGodRCMUIIcvk2kTVczrRJSGpfCUMv9unAAgRp2lPpoBtZnVZloSlXdHNHR2y7Cs39ZE9lPB
yz5RYcNYi5N3FzUQAWW9yT56y3v7pcJpjtram7+9gE1/JybDsw97lZuGy5Dn+jvaf4Nz+B+roMy6
8J+shmxjm1uQFqHueR7gO8zsuR/kUsNyo6JCU4A6CN02Hrm5PaPctLuEu2I9kRIW9tmqf0aRQRqy
NANpyYmf8IUO91vUerQAGkL3C0XrvS6WsWTwtmO9PqypPYU1Buy0ao+PqPWItFGD/6CjBiQ0YdQ7
B/GTsjc/uh2zg44FlHEvoe/ZsuQCneAENAwhBSNYZsCnAAdkHvaEv0VKeRfxzC0lvKA/b/axpXm2
Px4kS3Jzgm9MwWvUU+DcqWlYi/1arOOT6Dwokruur+tJnAUz6hO797thcy9R2WXnYWOgvtwuWdCW
grcdIXmz08NeRk1kh77cqG2q6kKRiPmaSz6H93MsOcYCnedZlTFDbvtLgTljpW4Vnz43oeWiz+BJ
K2nZm/7UMDROeKV4Koa/kL7YaMqlZeJl/4Ilmp7j4qkYwS0txGFn+PsAH3L1m+QOX+IWABPTCtau
vf3p7eqYt792joJMuvDrYsH886J+SCn/rvKL5Wx9ws3KQ2FdmW+fiZwcPpYsdolk1C398wmzoCeK
aXxxq7faZXuQ9366c6o5uEHYXfVqsJZ+xJed/BaWorA5u3HNFg+F3Gt045TF/f/Hlw70DYdxsFH+
uSmKGiPqadJ1yQw8PLTgLBCtYFuJT7L7zUJ29vBB6uIYBiABkzrrxSVqYzvAFRsi5FesL9BjthmR
67i0/nW3gg2vitCMATqzeoMQ0f1hMthPMNUy7hWfKRKyVyAMp5hNtK0PMx2FGeQ3yZDZf99RrFqW
l3Vy/rGOu4/EWBdAnnvb0rGq0chC3FT2RLOSKEPNwU3WwG8kvWFc9DH9+9U8el03937WWRW1emva
x8BEeDMS5dJI+LxxM3uBdmUzs6s3FoMgqejoeX3GQYHFD4vywCATcOm40wcV/pRR1HVW+PjaRHx/
X7HVO3NEdHUjaL+jKYNXYFxMWaRMzPWqDUXXw8Fu1pAy745HGOTBFjN7UCD28asqz+mxRAnP5hqs
q6Qfa5pfoUoZks8GBQp6zc29++ytD2mQrcX7E+D69csY3cEDAmYicSJy1Lw5gDBK/bU4tl/0TnA/
4P6QbYkC9lrqGF/wGf/7T83mfSQ+KLnGvcjFaRoQySNoYPUGWZ2kwHcSJaxGrGbG2l2wlv7FZuVh
bLfsnuMas+FU6mww8xuAAESwYCBA1AEeFkwR2CFYJkgcKwccJ4T1IjFCSQj4+/mGK5vf/1uPC4Zn
lRDc/m1KqK86f7J42bYxdBmDNcfbo38Iml9uaM5msyUhnAUlT42mWQtHlEXJeep6tCcI2/OpCVzu
XB6kD73PvkyxtBbE8+u0y2H94jsZ5p5O9sPHmdUX2zweJkTIgWgKX7qYhsU47ABIV6VX313UB3b7
e2ajAEswiaSSlVYxvkz6VPoth1/9h5aSJ6bRLHCf56doxSNPaSbXNROiSar9LkW+sO2cfhj+NwVx
aurzE+NbgBASgg4Id87pcabBrrmvC46y9CQsLualF0nZwsuoteodvHyhu42yQcTaaiNlnsDqf9VR
8Lj7p1ryeoNCMjcLG1ZWoCt3I/gUCUP6QL3x9vZzlq9w8S7vcOff2JtXft6kf8YGuoHB/pVlJBzK
vuZ208mSiKdvC8N1Ia24nM2xUnj1OCitpkFAumzJIF0zVLnGTlQloB5pRyyUg9ujawoA/vjQQXZn
sBx0W0JzxJ802+YQahc7Z50xJpvP1abCdNS2e4uJMdRklq4RXdFsMz7GD7bG/6wgx8YSxVj8UaUK
+od+pCdY/9aBhkTlJos/rpJOW9jvwIDiVMWfaIimh972YvMEQubwWIf9NoBgn3aL7q1afqxH2qDW
J3NIj1tXgfIT7uZFlv4+t0jfrM57QbFaFODIRP2AQPeg9g/0SxFW1NdCDWwILxT+tG3ImbKQofKT
wHRRO9iTQ9Ix7x0UrzphaHbRvwYzEVqSLHSj/32GOu8HqELhi5rOg3WDCk5Vy8c1DjXkhcyjX0LX
Sm8ePBZn/a9vjrQD6QVXSPm4DtEoKeFqLSiKZigTN65vbBq8wRxNlT53vZI5Q4R2wHRKblxZgAK+
vK9qY3dxfPdGtHiF+9fQ5UC79NW6o27CeDeihs0GJPziLFMAJ0qKIlDRlWS8MKvvcxgNMdcejrik
1PR9xrikaCXpMk2zPKukicUTyqY+/3EVFYfQH0GCA03bkO3aaB4ubnKlyoGYpVHHJdxwYl6F69N7
i/JK8LwKq3ryVkJb/8hxc6wYGOAfSHr4YLUjLhxo8eQh6WLxqNqncFN6gauLRCTsRvyG/aBDqm2N
X+0jhKjMY7/qt15Zpy9Qlq8X6iRu95CNh9AQmyMAbw/7JntbSZE3GS9+3FOH2zyGXDF28zZ3SJD4
3w46I+e3qeiPXgrsW2RuX/L0PFk88Hmn//d3em42IlUsPOhmuTJbBkkvmqXOpiIxlYQgf1DNBM3q
Ixv5JLDvcmrudCd6Sil3zuwAprf9HhCt+peMYC1jsRJZ+C1qbAYst5nBx+0K2wqflQZtuqGOAA4g
8RHLySaC/lwPpXOOKQPljahlYsggwZuVBpVHwFvOuyDzuGx2C9SHCA4AEAtKoECpCO9CHpgsrteK
iTJr8zQnIqPE0ODtQvAZeYGunfiEhqqCWQfsHKMP8puuhaq3g546qF+sMJ5ZVGdNkTU1kCu/aadX
QdN/FLukX0s7KBzwgd9H6qca74DqHag9Cl1qfhg26Pu65s6OgVRFtD/llGKaBqn0NzyR5JT/mJL+
IHagfFdN1p0EAJ13EdVRxAvYZWpLvKtD9w8nRkQZvTzscMkEfMDhJL+6DTpIvNkoGh3LTSvBwRz0
CK08OUA+bvwdPYRdYd6iws7oMWf5B5EexeqbHssS+e2FlBUAtAEcnmuMkoviMoFjC95bJBzAbC/F
/nD1qJb1TkZU7ct/K//DbqrmTpK/qRafCCzcKzQK+cFUswt4hIbED5cpD5eggAdFDD8ff0QQJ3Ev
DMXrYZL/4L06oMkp4QKG48sMFQCsYyz4A4jIy6szNcmOG2dvPG03gUYv6PTdP1nmrEfRJMIFMiQ9
UUII4Gbq2bREZi3axUU2h6GxMVZrKDNOTlwvraGCw+2AhibqBsdeqDkKsBd1nJCX/TT0ddxkvIPL
AiiDa7K1BPDSwA3rtwP+tkXswBfYOTKHSD2YJAcsEcMx+oXAJcLyKnV9mmVo2JFFcQELTh7qk6BG
yxHSVdWqY9has1PLckezh/u0tPmmkFsCLEuzTW9mWjYDi4rVhBm6BY6EhR5Q/t34W9sE10sC67fE
JKN/lUdGU2x09X15RdcA9ypJFj0HT8P9W2b3iUqnCTJTwjAIUghReDaWDJ+A0+THjN0iyM+Lboy8
QwxY+xWw8dBzh3UrDI1JfT3o9tBZo7+vQ0F6w3/PnxHN9uq1/ei/YvGp4NkpikQR1IyjAf9fisBb
ebW8QVr4m121AYhEBVdxQN5pMtYTbQlWgiKLYIWvxPlgjjUjZ6UQegzw965i4+l9e+hE8F1Op7w0
aEbn0wiy75URrMszXx9GYq7n0IV4nbvUp7GMQjxMDyRjs2l9EB6teL/a6LdnRWV6TucAHlCHFbWd
K/1LQ0iwnUUAyCRhE0NK6lDFXcOmgp5xo9gcdUvf2XOhiROOEfYeWnrVVwwyjLIHLZJvfythuor+
5+3Yi/L7HRgN/YFh4JdkjDRUD2gAMRWRQ7I4xGf05b+KE/Q4ddE7gP3zWiAP92yf/JrKgQmCOFrr
BZ9IxvcNPZxuNeYfSDHAl/O1egvB71cAjm86G4eki/JiklfGczf5x+GQJOA54tzohm/c8FjN5z2b
auw0RBqw4S5ruO4pFJYkDK3DQ89uj5cgkJAcFJRAP7Fv19aU1/Ysw6eBmkjG3i0AWLLsFNVG6ZSd
mFB3xEeLm8PCPNPBBJqjB+8IZl1H5F9jQ/23OdCE0eqg3H2eMlIMG1eSP1RGnRxfZyaPCWfpFLxj
t0sfe+2irgmBzpBXSsIZhzBU6NGKU4mWZS0VoamGWO4loBffK0gc87kDXgHlTdveBD4TpbW4tbog
hqtBTZMPdfgWkaiC7P2Ce9qjzOAYUrA31YAg/iGdRLvQLa3hgyjMD9V1CEY2/G6pNfd5Ocot7sXD
WWcV7+NtQFdytpLfFm86b+MfS5Z5X0qkmCNU7NPVRbxTJByuRRV5Nb9vr69L37yl55pjxJe2jPrc
yrOzckvGjyiiMpWrTaQxSWW2lvmZuGm0ot4+mvi+fzFeoMWg/7ptyYyJgozol/N6NcioeLZ26HYC
5jxabge3V/Nyvgwnl578OCaxHKcu8casttuhBi3z42eubZVs5vDUrmka52F4ueeZlWeD6xiHCBQl
3dt9DQlaPwpMlbvpoJAI14+hD8ZlmAXwQ5pd8r8FkjvYSHfD8ZS/E7oYYQlovvhCP8encFIlyuoA
5x3uirETfNYZOXeGSt4w61zLoWxUCrlZKhzJgMs8NJI0s4++FrQL07ufrd0gXFeugQHbTBh7bi7C
NU+OCEmjdjtGIlro+cVF5RcsiTKEr4lmk3kZ4vlrHIb+7XSnpls51PNkJUqrpBQhgQgqjAYTVmCp
dZ1xn2C+wgpheg80NHGwJRIT/MQ55IOtR9YLyVUuW7X2p5+DSa36Xy80BOpJmlvfLurXfaQwJRvW
aEMCol1yNHwlPY6evlwabLyuJ/18aCzvr5gklVmZ7Lf/HqPkgaY3gId06OqeQxqrDRliviywVR2O
QsRguadqFIK5jRrLMtmE/V/y8j8GYGNf9MXEcJTtoxOVVuhwPMHFtY2RqAEu3O8c22q0xePSFET/
52rI5e21Y3mfHSK9Ei93kpKQkoIUw2SG/3yYrmqzMs+LXvXlt7EL+EOvHxNj49Su5tqCc0n1w0if
hWGoNOFG4eqkt3HEHfRiB+m2FFqQipTGmCMxUKCznsIQqunBv6dCa0S0mvSOtKa5huQWGnWleQ89
1AlpA/hM056b0ydJEmyX7bm4RyOUzQsMGQR7GXJxzPxr5SPJagHAY6qgdWVWUXJK8XqBMoWxIoGW
k0Q1FxJzoUINoY0MUSVsrTKBVDots2h2U1+qWQd4MrG6u/AeXctX1ndzBdjxif3hRbahVv0dWXRW
j6uR+dj8Cz2Log6jLUshkAeqtoOz1NwYnuIzVdDvSl+iwBRoJUxJITe4FtnXjEgtJnsxS9HKRzPh
EUSIUaq9cee+JFtYvE7IXP82ylAvB4cfOuZvG1ekT7Exw+p8MnzpPw4/dM4r15ruKd4IcFQsO1+N
TPd0eIhhpwFLQpt/PB3CGd+SPFcPO8TS5avEq7k0AnR0nO8hI65o/kk0W+yKZLoq5AyYARYVz6ZA
lpl7uj93J2xyzI7G2bnhNuvV19qkGvu/901lG0gaKqdSVSK9nZa+HmLTmKT5YwFLm4J2TcCMApGS
G+EVRPaK2drQlQlvufabAMPf+GcyD0PfwBKAthLGC/FLxPBS/QEdU82wgcH99+mmga4FRPb+dbYw
G/ICvp+g+K4cL3z0Hi1f1C2DVKAdGkJUTDdc5rMAhhxlLtE+Kb3g7y6kCnQGCzkH4eCCuGet323v
IVRg5mviIxHHekwmi/TMYf6Fg025PaE5sXV2wHI416R4r8IwBj1x7ggxaOJToT0wwmTJcsPds5yD
M2i9joeP8kyhrxwXutm2HXBJhXPQGKnGPa2IfCoHHvD99noVWfXhTuFuNP5NXLZ4J4TM7Ql9jg4c
T3453kWDIOAdFxaPvYgbdTyYkm73rUUkcFb1Ag18QGywyAX7JQ2MLkVFSgGiFf/HAY0trhT/y0jg
sVmm/oAfIG85ZXQjhPcw5/nXxmPP85xi3DbNIIojqOn/OjOeBRq/TXpEfUnbCkC6HZ6kfX8/UPXn
JY7l0OBXYW+BqknO4ptX032qkuRPqui+Pbig1DM8rRPsEGTozxOvma3pZjc5+iPF3p+5dJW/BXI9
oVLwt6tAbmvDBp8F6yNk/zImUDmknakca+BiGJWKmcKZ6DulvSPiAYnJxDXJIbY7e+HfNtuTvhmx
ihn+F1k44Gzm+3NAj80bbrIeLlFpZQHZC/I/ynAtc/Lx2GoZmhBmdmyOfzL87rwUn7RCyxnta6f2
GApms8cSqSAwW+JCdUf0zrUwVWgH9Gq6ANy7KbY3eB0bwndj5sUjeKwgzwpSfQrARPAcROkuGb2S
fab9yBDuSpTwD6L4+68GqBGDMOHx3czLC9juO6QcSfgzMiRk6LENO0pEdVVjmeWmnrloglpWRvph
BeS6A6v8wpv3JQdRnnhpg/XSRylQw4EHPCSmcq67PyiL2z2WZCGUO0RT3nRPs8GvlD7xRZCJnmE2
hVPkhYvqrzQQGHK9dogdCV9d2D3zNTTxUQsyt42fe8y4X5Ypw4oTmQOPrLru+WNlpPlTuwJ3HX8V
4lG/SCAvk68zqJ16rk82mAoCP45FgMrVHXSWK0jag7b/bbiedb/3FZgkPCvRzmEYw6cfA+eNESOX
gTa10iSOHkzPM+GlUMo9cxlrRWd2l5MyzetksuqrE1cT/LK7Rvt+mIdS3PhSEpLNWQZJm3dBQbE/
DPImwK9eM4WDeBZvZWAEFXldYfthD5NihhRlTv0JAMwDXhDHxolPnwhPvPVql7u2CSo0esAttH0u
4ZFSHjJM+Ru0a6k10zjvPMGHY+3UAidhLPaDMEpUIsWXF/mx6n18RAbVA2U69fF+g7GZMi+I2wJZ
J6ZrE55zK1H/t0WPQNZgXZD/N6LCafPU3ZNlMtIdXBvm4eqHiKh0j/ReiNUOVAZCxrNGd+w2wN8b
Q1g3GpHn1rKnNM3cSbZEJZGqm1XZTdTT2SzPIJSPJiESMpBD49jaS/zhZz2J6RLrnTaVQVN5uZaM
v8MAXK7hSVwJS2e4oqiOE6xGXlmEsxw9LaHCBdlP7teBrvb7Zh8aOC0YKcVGrP3iOdV3lSK6yuD1
ZIKVOKCe99/YZjiKjOAzmqHVnSwpZFLbBOk2esOTbcPJCHlLzdLAinfMb3ZcGdPrDpLq2hDF0D4Y
FobA9fDe7fD6La+PI/jb1kkh+oHei4JFRCToALJdJHmZnQ5AEKbp1B3Slq96y0EVB3a/5bJBTKFh
y1sA4SHett0aNwKjs4GgZWsKyOSOTKTovfSKCPI2b4Zmh48hxO8Gg2i61KlupbGfUWCD6EZkEg8Y
My3+08FUeGH8L5vgjk5vqQR1kn+acdkDUIxL6YxrdbT/tZUw130NDWirtWCFqgPGk8CbFpfpEnhi
Mrafeka5wxFjgDj8fFt3Lt+eB5h6qiEhXw9/Pf0a9xxFSqEZo7tkRxrMVghZHJ6EN2+Ovz3Iia6X
aB8et2GcNIOeMYcHsB+hKEb3RdD8xQ13LVyCgmFD2gPj0dO5/6roOpdBZ7Qd/ej9RCxMJJGcM3Vu
X6GbXEZ2+bmhU+30Ib6afvL4oZYiUuQWypueQT7Pw1PDOXFkGopw5uV09RAmsz158223M0hkifjU
6jlrfcCcrRpLZV3snWeCOr4uHrgh0D9gweH2NwCMeF8iyG30Qc/7K6Nc30zmwEnX++8cz1Xaq6yC
5rpFz/2lH1mo7ZNIM6nkz+xE/htW47ejW0HFFzi1RxYo4MQA+tTh8rKz1S/GuzPE/2Oba3WZc3Kw
aL170R3LojvNvwVfsl9ppWnUmdhHw/6M4t7IYjOHge4pvWS8XW7NpekUkFugkQ6Wiko+6I2WYXjA
ha1ypS6cPWcdb6hx6l3EPm4cXzo+TrMBA0Bdry18aNbY7+ABctFdxPLDs3Nos1D8+Pt1DiUm6W+Z
5xpXYwxzmE6ZQ7hk5iZwrOnCUIveGp6bggIGuU7BHO4NJ0ifGOAsytRun26KP/aC3M0Nqy0NsuhY
J010csfjF5YxcrVs9H6rs9WEGrFcQ45Apxn69ZsoAeTpvpY7b1C6XTqRSuanjx6pbzlaEOou8YfP
FVJUtGw8EZowm8J96wsmQP71y4kDfyz5w4bc8obUl1jiXCavfzNISd2xjhVcEb24OFWUuYau8458
61ZL5lET3vt/dyXkqMCnk+WP5DKS+awqORNWETrr57oBfV+8+MnGXNuDBpKD7P98+DDwI23QOUnA
f/cfBiwahpbj0bwr2YU3n7dh2R9RRe4seoSJ7hlH8iPIX2GnbklQton6KIuKlaq0foHUi3Q5Yj3O
8HjlQTlnmvopkH84MLFaB68Ro39HB5YJXg1RTpkt2mpQB/W7P8Ild4Wyi0DNSn5ZO8fMXyLclrRX
r/uU8a0civOQAeUvt8if3WvQ7XrdyO3aj3V2BTiktJB1oRmy9zKLcohguCL2S7eADLsBss0raRg3
/bEKhJAIMbtHKtWJLLDbi/fUJBVYMWGYDOP/dI5tN9SQeDCDsOMACcRXj27aSqX5Sv8I398ZrMFA
gER9XltwrbMIdQQgytCiPqhIiBYUrFTi8c265uNMtgqJvBpQ01fvshbIBpTiL3AmReVlAsKcinrm
tP5B73huWDhkX5VvHz/NFHVcnLkQfb5A5baKDuK0sBD1Jj/NrutjulrehzDrnF4WlBh94vV1Z+XR
QRpYHxEVOsi9wNSZQcBGgYDzeaBAqFX/gC920H+zQkShljGPwyheSvqb1v8SR9AwO8mYCnEN0VKT
TLY3gPNw8R+LseDZ0G6bLba8NyTtRjeOfeAccBIy3rPkz7Bb1eHTBNwK3E0gTEWW0GerV5HouBH4
rcmC+GtIMGLPcDQnGEcFdzAWck6gRJrkNT4jisr18GQ6sMoliO+DuXABhm6AJ/xtwH5y2t7eiPzF
VwgaPRYRo4bxd8uRnsT0KnhJ0ZaohEuN1LBtaOBv8Wv1nlWl4K3AJYea7Ck7wrU8JlM/zKGLDGU8
L+5HVk3Nc1bGw86+hP2eFyC5LVKAcu5+OtfWW84zXiGqKqN7VFmg32nT5s86GS4jndcS9SSU0dG8
ERkKol2CcSziUe5HPnVPUFq7B6RhUwy5ctl17JpPMYNam9mU2q72WzsUtT79x+M9h1MwpbdNgU7m
jKd3mlPD29z4CefzPGp15mpdPDktUNUFTrxuxtpdjUbJ7XeD6XNtqoNDtJDt+Mw5kqBMthQEokio
6GVjhD81gTSQ1TjTDR2RZ5H/vGX5GblD5Fk+R4THg66QAIhkrprxlaAxjcb0RP1O3hQ+IisHsCvq
lW1S1xa7RfCBnz2CWApOegLEV1Qxfeg2AX68Pg2aiFaTkSS09RK1muqQ0+tb+UvIp9QajPb/fR6P
ppyfxPIi0dX3CKiSA7wbprtEbAjfOnHRnjAOdQeJZ4r1Lq1tvYX4+KFbjzyjZZwS3M3BttcOwgDE
U6l2pBYF9bk6WTW1siCR1SxdiQGaNYgHvZBncOBJvN80hDSDBJw2NNHtQ1Llx5Lzckm5iUHUjyMk
6H7Mfw390/JIVsQJLeCI8PFhFThA2U8VK6zdcWLdnGVovdVzsjnam/4PMmqatAxERQMD7qzAHYl8
6Sm7vJkkq6PFWPMxJo4c7NDqj2/90L8zm2oMZYQ4gQk1dgR9WiC+/+aMPJfseNSYPf6U8DuSztfU
ImDwNuabMgKBm0GeC8ux7qaKxgMe522b9XDTLnTRCC7NQSz55C2cTll6TEQSn64dJtcvxYPNBaIO
kQpT3y0R9o/SVHlYXwEtHMNziCSMez/0V73/alwoAmNebPjFNtCpWA06yk8XM1DeRFsGoLPWuT0g
oTsX66ZNWdBCS1yupq8FZD6sj5xJTn0cF/SA7f8DkaAbTJbAloBOP5A/EAilYrLqNRWUC9R3dNRe
vnlk55mpl2ecJEhweAFS9RFzb8Lvj8hPBebqiPlx+sX/j41N8a7iwVf9PgxLD+vMrjr2tk2zlQc/
jaZc+r37sxiW88nctqe+rUOp2H4svQRg48MYHMwOHtjg/NhoogUe2F8hshnscV1VMHFw7jx38mZ1
rnjp48H4K+gibFFNFLce6R1x17nd8s+xoHWsXc7O3fJ16hoHEMbe2beEKR4m+XqrlHXJ+97G2cp9
7whOO0YGM2qBIOs7gch36HPOUHMbL3WzICAmgCR4CG7TpjOaeFm8loMJXm7dEooM3PQ5p5Fs0ASH
32BQMdX3R2KNQIsmD1Er+YoZm9F6r9I/VR33UD5hJJsaBGD+mvN54DKVjKxAdveOLATgWYVq+uAy
Ba616N/vj42D02R9seq/TCc95zphuRRlPJhS8XhfVaDTMKP9UTzKPVBVYG70ba8lQ0eWWWtzbbg3
fbnyO+hQ/v3Xi5GFtQrvYtIgo42zmSIGDp3kVRZ49wlrD3WrttUbZss6gvtU2AQVGX/YHH08Vfum
Hu4yEU+hNgXaQ6979IPnNyGpnXLkWt7sQk/Y/Dw91OUCGkpzOZ3gNTxwPw7JpiUTGZ4OHv4ENN+B
+0YZULH5HZOUKf8KHyZkgssuUrhe3D0yg/sbnQVH9/eE1GY1qv0S0GiCMT3mHAsOoxO7ed8mhEXN
XayscF9DQ4Cve9QVV8yRl/ACTXuXmpksAgbBnkwCJF1GUgKsoVtA8omiWVbP5UIHw+RUKQS1hPP9
1tNvoo3Q/EFdxwkOporCbl1m32KmN8at5XqlwUmCEANt9MMVCx6bf8Glg4eqqM8NbNvBCLwHhjM/
mNJTa+DyH9RN0zsqnZEmUUIC7mreKj+Gj4+B4+BBUN9e9dDmpbFcbK+1n91WlaG3fFkeHE5qLXbS
UFHzxR85p0Oi/OLH0dibmnBeqmO1NFTVD8TdhEaBN15uRKipjq5BKzeDBr/8LU7RUnTsAaKu8iKT
055jIqiUSoYbav4XDEAz55oKyYJzOvpKoEA5zpSC55gWyLO0oIkychlSQI8qazP+kk0aTOKCQCLx
AsP8MV4NCpZ3v4bqUuf4Zg7OyZE7I/5EHGChwnf8OnQTJrK+ebwguDpNyKE/YEX5r9Tn5xM78eis
6mSX0NJ/d3sHjRxnA14G91OkWz8pgovDIFq6afd5eTBmeKRfKUau1jRml3gW9g4CfvoUyX2xIQIk
z407qXsvvvhbIEwQ7Kb+54Vpy0IyXRLBjIHDMs8XsI6bhTuN3kDoflQyIsP2l4rHpXsB9WCaEQL7
qw8cDcj0UXvq69lo+t8SDsjxE7tFSh6ywBJ89itEU8SkfyfT1y7laxyACJNmDxN5Mt1hXOXLvv+x
lmFF4Ei5M0n1Of3ur3IXvVhY0MPt2ReC5tbAB/T30Fj5Trh7Pcqri3TdI7K7CDaxt9F3sD88gVK4
WZ94ATFB6KWd0lYjteYteiNx+3k9et6vBbGdwrJEVs6kFA+tMJObTDHh6UIoPkHncP1rLEE5D8o1
DLACGcGz9NtbJITdH3dgj+5YEN4Sr/PKBA9Ul4jZidsnLw7q6nQaNw0z3qlvLhBT/UXl61a8l7XU
D/kJOewt83qVXmeqtlwEEaUphsliVL42xlCdUCKFdNpbKa90mMko6zHYsuJzapOAT/NimWFTorPU
cMEMQzfHyiFS2Owc+MFf5G0bjQ5t1d9OgfB6A8yj+F3/a3ql6ByP4d1BSvk+1zh13u9OP03VikVu
tm5I7vPGWuQHBm7fbfqoSY/pHCiAmEptZu4epW2lZNboAE2GG6q2aBeeMcLVK5MFpnjt/rLvH2n3
Ot2uBZOtsKoFBSGwWcl0lYcNKm/CcDoMhee5qy+yPNx0FwIV54BVKm/GQ6JxKcoypz3N4dWLyW8c
jXkbka/+j82ohOQR3iWj199U54Ag1MKcvH65VBKig5jpPIjpqjJ6EOKmiKWmZzfImHWdKGgI/aDS
rsNncYho0XmZV+Gnde0Y62biqvvTrdrbC1/v1P20xasuvklsFXneAf2+qP0d89S908F4Y3E0HqEW
ABidtjfz3PbUJ5dUXfqfezwv+ukTSuU+S3vWBJ1eW1mgfP9F/XZyZYV/8Qr8M21vf8nGZF7nRB2p
3u0u0XTwmdIif2vWXuw0VeuEbACOTpsvvz4LxuPIeRmEydeddmeomqrHVzI5OeLD2wq2lcGuVVrY
PMNSUSsr2OJWGhfpjedar7dhj4JplgmrYV+GsezgrF16KpyzXjhWsXDwUXuf+UKscohAy+2/7ZlY
SqRC+kJxTpJthnnploxmY9CIcYoHGErxNOJ7w8OM4peI/B9zI2Ygh+ombvvqew4elNJBZ2KhPEdX
/Ly2n65/c3Rv3f7WStUyxGmca5FVdp9xTx/GZz+1ZZobNN8lmfqmFGgVwIrzkpyPkz+po9Dk8h1g
bojCmnlGZY4xGggwPOAChI/zhccoulpbA8CTRrQ/bIHFtzs5AjZUF6q31cfXoZCTPXIZqtWNTzo/
ebNSGkU48TdMp5xXa/jgAyXE+wBFwdkmiVwGfpSBvEQ3jiVn0h4z5T956W+5PQ0Ll2uWURqmJxVH
iN7cW/rAuIYeHAxSjUpYjDOQbXHRP2BkHYa9tf7epJyFlUopEGmn5G4NwX6bxgLm/f3/DNSVBm2G
sF8Ve+o10M0MXf56JI45qmseX1WWAidS0OO0mwH7upseXzbIWbOyahNfmgDs3kpwe411nG6lddnn
KIeEVDZUe3sspWDkSyR+96QiBwEIs0SvHMtHGvl1aDrNsr79lZmUUbmy1aZMNfuTQxo6AImq6EbH
sEBJvSEvuxJM+rq8WN5fGRgM8FNnSCVChyUMigyjVcolnH7VtnUH0qbSf4lPVF0h3l5/r0C4xBMM
ZeNbvmb428p0ndlRKKqqR6AJf1XAGVpVzHFRNhvLRetOYAmFTq2CB6Agj0ebXIK5hU/ApTWYyR+5
IPOJor67Qg3T+sZNI0Z7MqexnoC0k5UsT+eghcylXITDgb/HyjZKy2JZRut/AHcS6Up22T/61Xjn
KQcMQSbXmkuKmDrM80m7Pg8zkIVS7ZJUTKVzk/jexc7H3vFqxZ8dppVtkJRpW1c0uinvyJO5crvO
vCSC/80pHOYKFbM/zwdgzHgdtA10jphhC0MAnfhB/pZ4qasqQLhstiJj/QML+b3ZsSRtDigcBPuj
cPQcqbJbnSzFk71Wiq2NjH1ACT5Fk5GoZl3JWOq6JoNf+NNCaj5IETSV1KQ0lez7IG65FT39Pwom
FoN+Fg0IJqjGQWtec/JuITCo7W8/0f3skY6GHDC/yHF1cvVcKjSm/qj4bEN2D52suXdvblylew2Q
GAl3Gn9wjaFfkItpAEo/aSqmO/tkOaTNWz+BllL34hQDjuidOIDZG98qW1wRy8XNWUVeWJqgnUIk
mYlmzs4w0WeZGAqdLPVU9Tk0XT8YmkdQQrVL+efbf6658ARqnzJyqod3sJmcCIfOp3NdwzJKy7pd
RYNzmiWjm/8sjUppQyX+tNcTyYlJyPkfOBamcVp6mZdsiD8IZwKXEtDGce80IvsohUhsrK2yXClg
jKQgK+AjtDwqI56EaPMRmKspCmuzV9tx7sWMQ2pjIhc/GZ+fsMIw8Zi4mapIaPFQ00S9N111Tcky
nDYCk+PoAIqALL9BpGCTxEnWBVsJLId9oOGcYlEo6i7n/XU3N75npqdRKnlfcvhKvSG484rKH7IC
zaUPefp3GR2tIBkWuvFkuRO6a/JQU+QA9Zdkb/Pv9w/xojYccNqyeVboZinHm+UR9JJH+a394IEO
13SzBAchrgg9NdnLTLQLG68sOKcJIrEdh1f9+ApHL1np4Fp9RRPr3uLvRTh5J2ebSxZZNbhcSVGN
uc0yjV//bwzXWT79ME9lWh1TT7LEQNj/F6SQRDQyFo+gXvsYTZt4ieJJVN1clvSjm+8DtrU1uwI3
qZbzrsCO7RPlMXfRb3cVQhWp2QeYR/+3b25T1qjorEnuk8EBX7AhKX34BOjPccqBRUltzBsi+KSy
AaWUz6uAgjJSbk+gB+qzQcsXGTdd0euyNXhPnZ3FL727DNIqeSGsjOOCBqPxRahFoAMDHAd2HBi7
nhZyVDG2equMJcjC/jvL2aofCFhzGq826D3xaNrrhD4N435lGbbbXoNe8LVkJSqU1HfjOcqhBxnq
BDqtN6JznDFDfomPNpNsKkawPkTGogVsCukh0zUzZ1JLLOfhzMyt1HFxhJBFuxeSVS4H+FBgekCN
UiGIY8/mBz5xpPfi2sZYWpaXv2HtHaOwOucdMf830CltiCVm5bXhAYFtCTavNXAFj6428+NP/I2J
OB6pfRBZI6Ep5KNnjXcuqbmI3b7KiYtwfz5dKPFPHWlQZJnMl8ELmuNnqxie5jvEVcKTEwfGq/ib
LOl90nb4rqpJLxepPWTLADje2fSauBHn+pToNTXQD0cdJAPm8MX/DV3f+x7KoU4hbsV2V13llZQd
Q2FLFDeBdJuE002QB+1AKGlALI1+TlHVeHuzfGVy9ncq1JM9EoWppj3lRDg7sxE5RmvQDWpGhD9c
TprM6yMArGNp+N/p6BOJXdimcNjhaBshwpny+n0Df6vz/4IVBAa+OlTL19YJ3F+lyzi1aKtH0W0N
i5UdgnLT1mjuNEMWTpfezThRKiQsCA15geB07hQpZoA/1iJuvpmtnA0/nxf52Py5ZPyd4slJdyYF
gBVfuVGxJBWN3XXszr1Jv9sLxrBbvaGEUQ0sCyJ+uVhnViWJ3pV66DUdS/HvirRXb6hj1FZ2iGLa
gZx+PmpIKE/pQOOSl1l7mR3LPkL9IiJbJk3695TyyzFZfcI4CKer4VDxWRr+8I1gW3cZFVaUECsD
r8rApVLjS6/B1eh5pPN85nR0FzlF/4vWUlhXh8JtKJo8cblab2J1y8PcGQG78ktwAq7LTsQK0M5U
XCwE6NJpVuacipS9NBAh6DC978AIn2C+ch/gSaDcOjEMXEpl7CemeKFh/q2yKUgHhGMyzabbfOX/
nvF2r5TPg5Rn1T8IQhmj7fF9wL4JCnhQp9roosuCmlhGM6jrf2tbwli5HeVGzq/+ItBoYJYDSGgq
2sgkRhbYEMtDKaaAaduEGNmDdq6nHI6Y/PThJfw+5LGB4fp0hlnqC6o9ANgGjEH3wxII9Oa4bZ8Y
XIqlsbo/fz7tGh9obfjQsZ+ZZVDWfX5J3OqbpH6G0h60L72IiocQJcjI9IhBIfFKpVvIMNesX7kB
rRiZQpnKgv9hT0vcTYEIxtxEdBzB4A6Xr1XVJ9fx/YqWcZXBm0uEA4wt+atizb2hQj7gH1YYcMc3
e1NHyD1prrX1PTKz9DHk+aSsslrtb0I4I1u3S4hv/jfeymU5H1gQLzd9voadbkcr+Xf8ZbD0+Guq
3wy53PpWejlwPuQRNUaWAf9caHkMyDfoC4p5uxSxJO/0OfmNMio5och4H7nRpjR6rPZeHUE/NM9B
onUE5hxJRFa27yTaHbJR3h+urpileuwl1muiLg3XT2XpBBp6fSd+Xwe75vU39Fqydc89r8b4x/b8
BPxQBDBdRHrUgjT7keY1fSg9Q0f0Ryiz/19x9HAQa71mqW7lXPINKZLLKFlrjoDANHFjawg127Nx
cdEMRYX5yRFwGKnPGp+qclDTZkzQBcOfFFhu2Zzz7T1TfipuXrEqsivzk/Yo9wkI00FfnMMSjHMJ
39sdXOzdd7AXW4S3eqX63vnjwpS/kXWGUi5+RmJ/NG5kbi2LrEknZbGkxA1OcynEcJJTV3F/PZeQ
BFluTps9NZ96RD70WAA+WbeSb8r19R4pfBfnbkBriuFeT7rdrbjCyUvKr5ZjsEw+2ovgOZObiN48
KVKhHgt7JwRChbUO0RhCAuPzGBR+CMyTzGcM/zlyj5GER3vBOQ+oMF9pWLrC6BNeXYvi+H0Vbdr+
EpZZHoI+OQIjL99m/NzfVkUTyR5ecHKfzZ1H1L9lZ+M570q18ClErAHoXqTNOX8FpVz+kf9V69Mc
a/GdWuz0hvJoABns+/LewSOuOs0VjgpVvglzYsG2Bgg2tX1u9A/ZEmBwcYRAQd4SmvutL7ciDchh
Lmc2cCkxnFkrFfzQsMb8dYgTRvi6rl0wH9IPvRQxlaotZ+a63sLivFpTJE9trbUuMOLA/8CTpzFv
ZOtBsYDpwGCb0fMys+y8QmslQ98QLY0r6X/ka1Rz82Z53Se/j8IMGBcqPiqvPhypZCbVi8Dx04Xd
E5VfgNY5sASEOailpjlX+GSCt5yrRwtnvhsl2uCTT66V4u057oH18IHcIzbbOEKBNUpnXPIjAVM2
1aCxnOTLluiYIN+7k8b9ePuJfEfLKxAjq5aZtXsUIdJIoyN3XJjeox1D0BgS+vQZf8KR3J4YTTv+
nmMLl3X7fYwrTq2pYKU9LuSMqueWoclvmfijjDUiR/XmTCko49PvxWGPQ7PVlVkxSLM+QRkYTfpJ
6lZzmm38QfTgmrnh7rT7vUnHOMy4zyMjgguQbzHRW6FVMIw83e71rww3fkwUpOIILLNnYiVENaYW
4LFQCbjVk6lrd3BgTsoJKOUZs+UoB6hN5mKWJhOysF1322FzfoPLQ3RoddMTHHBCrwwD2TjvfYep
IPI1f44HPlDKB4rA2NPMh/SAPZJin1Jga0UhZu/7IFxtNBfZjl+twgZRdZDOslGO9rxMarVDjumP
gT144kPg3S9NVnwDNClQqi6ctzuV9T4SL+fWAzJ6wRljWyiwuKuOiXHkCz7RW+uwhjSO6UGlUz3v
KmnJJeGx/8gLN7OC3diLazW7Zy/7ZQz3u5cVzD9oYQpRKalNHt0g3Ej+nRdwp6JOzC28AC5vKsg+
HCkwu6FcdkCjWLBUUbwpOtYFUj8mz9YS8ncfV75fhMOyCjsnhhwj0A/Pa/Y0MWYou5YFtFzVVosL
AyjKvcmiBjWsKqz0T4+Ckz8V9s28/CQzg05SW0wP0OIJixpDKiVIsxMGVrmdhQJIokyCBqw/WTXF
Mm/uRiriGXOKWraBqp4sIOuyAk0Ejs6QaIJupsyeC+eodSqsPbRwvzkyYiHzpcpvFTMQmgu0IKjm
27j5z47ojOlgSnISM4PyllSU5RaAIgVGlSEy2Mh/sR6ezDk6Sx96fTv+4/WNklrtqhjApIPCrLpO
tz3Qyfnal9n3FYnsLGKW6Xd3kE7J5+MEIdKXYT9PdHryEk575RFy+ru/jU3PnaVsZ3NCNJVP1jKt
YZyR63en+6rzh7oEKxYIH1oUl1oIi8jr3cEXtUlEypzsLsagDjhtezu63h4TglrVj0vmvAgO/a6z
Xiq6KSHYW3iO4Xw77Cki1lNrbKq1+1Nm2X7ptkXzhtzlWpcYpIuCzYhRrDOM+o9zKFUpEtnZSZir
gejgygzCIOoZmE/2HIXzeZo92aUpty0CT5GELTHKPFqpEFfSfNm1ovU4RNLaveQWI5YVUiBqsMHD
MKU1zRxH8SjgSP+8x8b1XCksSE1jas9prBjyVpdPA9NUFv0ghIrp2SGO3RlEQjA6jGqq71fIM445
DNu5ZhWUVy0XLw2juKlRnORfMK2tiRYKhmahMCRDjxkX2frvosBZ3IFINhjoC6VmLbwGgkHUCqz7
EdYtDz7mg6QxHrPvasP7+PGYs2Me2kx+ef+hh2Ge28iDEN3T+FkZikELS/77qz7PRsSOVGRDUn+t
pgkM+jhRO5jKa8AjJaMkjqoLfgS/t4o75N9gZkZ3FNu59uu+E46tCT/A4+ixMDyBAM1+Hk85aOlz
MBnzu+iHnuCdTdXTTrY/AMYe2ovgM0HB+bv42p+sxQRP+947tS1g/VhhiisGzWOnuJ/1G15w8T3A
Sav0O5yyh2iWOQtMN3FHs9n1QR5cMO3qBRdnCyu2w9XAxBKTr+qSG8Dmnv/Omsjk47amBIW84WJR
Suj5hofMjqaVTYwMQyQ1/DTc03qpiHoftgajUnqgcvllbrRRtqJyK3ADYTtrnKEIMtRDaybPpDrN
6GFuPYU3ydpTfK6tVpNREGCyWoOcnsdIBHpXPCrrTvJUmJwzYlGJj9CCg1qPk926ZirxVOAh9Gqk
3OLPV/VBMNU0+MOwIxoYjT6ecIY0JBx2Sru9qltQU9Wfi8vqMn+pN1/SSrY+8iG5Iwvh5/4/O9ZA
lxR9y4TQ4+GhD0bv+Fn51Yeamzw0eQD04Z+iQp2NL3TfRYQB5YmeP0J67/w+Ym1axqS7GvEVJiF/
uI8KIYbZzy6BTimkzlnn6AIYUIP3eEp4JGbyJRlfdMb98gDZ1qZ4590OIkEmVqGytOa5IwwB8qqu
FTpAJ0U3dB1s8BBiLfU8pKB//Fi4CbF9d8xXpPkGVUmKYLMLZPyADXHfcRteLjl3/REMNGB9yh3l
Z/UzFn8lT8jSNXHSCTrqIMU2+JN9gXeneHMPeMTVObJauFi3kCGE95k0dDkASLOJlynHRgHov/3B
53mntw+JcmESvceCGly6woIjYtrLrmQf91vglS1ikc74A/OjxmwFKTxQAjX1QbCBSD3HafHG31PO
KCGvOCeLGL0wBAA77OzKrd1ov25kuexJGwBVH7Zd52zUPvq0pBn4PGEVLXEaItlJKm2Wg1o2nDN9
uGy6CC5wjc/aD5bdjljuoKcNu4KiZ7aptGxlLBSrAOwFMMA1RbcLufremDfkOKoOY3z18vkyblw6
fvPg5VZwsOXJHPzf1kRth1b3QZEsnKW6fm0dtxxYZk7eB0hLlHj5tNG9Yah+Z3psOFV6i2wsvedx
3D0NiiMVqtf1COHyGUggD5++vO1cbwoZyQUa0XXmNMqV+eVoIhhOD5GzR7QaSCBL+8O04cCkyZ6z
tnd+uTapQDRSzZNJA9xqFRKQiuf7i8C599BuZstp5I+RJ253dgljyLQTTW5aVzma6rsH83yvCApq
N3ZxkbLHOOk60WqjpD3OnlrLhPtmiIAA+uPdKXfvsw2fwFl2cuC/HSs5mjx+ZvguWOZwOJ5eoXPv
c4qKT/RcQURgGF+vVFjJw+tdo88te3xo+QeKfqkECZLiPiP1d/4n8xJs1E6OgAsJyfPHs1NYzvfD
uDrPInqiQxUviCt82mbRbjMNzx0kZ6V9jWaS+TTv+BgMPCMccaAInSWvOmtHxuJJ1UzdxYZTBp/O
4zEg8qVKe16AGt9tZ/Nbdsi+f5n1ckTRzcFJInuRX2KTenfYBwMT0TLKyzudPIRBz34HaIEBsH4z
UWERCKxYxsDiDluxYGXUcfBZfnj00dsSAFQudi9CMtBGRN3dRHmllnBjvD3o+iCL2FzM8UbDWe69
mHto900Bu+glkqymDMQwGO2phmtiYF4B/6rCVRYhJ6NUlC2514G9njVrhB/7x6qLmgoMQnuSZh2W
L2ywHwoU8p1rhXAn3NtwTjd+uTmLIy85Y4gG6reTnnPXGZtvVhrv9ipEDIjUHzySdmRkgu8ob0G6
CCdl88kY6SKIhH5SgXlSf6XRRxzIzU5Z+8HH6qbFlHjhyicOprot7gj5e534K6Id5Cr3rFy0zldZ
QU6h/8bZDtxJaPPVDdpfunOsTS2v3FjB3haK6xokIn5cyEUsAUeJ9mQv1PAzjaUnbV9eu9FO7n3T
f6EOnUnqmUTunLStrDA4gu8oriqbNWbA2Api6DslcJT6HDsmj1PLYVnGYx6o7L7TvPdGRyGExgYq
gd+2C3BbnT16t1OfRLkxk7cyr0xRoFrR+D3xGfpKctzyMf0rJonOdJLk5bL6CQBJOBpgJZ1V9azv
0Gv5cJbU7CfUbsvEQk6vfWqO1/toz+gIEHJ0eD9zbu1VCyfTDkpmyPOHyJU9q2TuV5AD4UWiAuwu
V/NWVZi33GUI/KeqLJGc27tjde8+p146Q65e4J/OlzkruLQBit0BE+U4FeWmVOckNyTDM6rxOX/H
DmI5VJVs07Gq7q8Mmd0COiP/edRFlFERmlbbxemLKDQ5VeuRRKxsk7uoPq+Qo9O/srA/HPZ0II7a
Jcw24fKtJbnmMhqVyfs1TQ7Q2eWiRZY1puAJhp9z8uMABK9OqY3OkaKHKKl93bLSLsoZsuc4ex67
pjXft8Ac8mNaaRFYmROTc7g2hjVBySnPAA86X0eRjR6B/qkmrmA/0TZM7cLbskBUS1RFq9QZcEg3
cBSu8fF4Zwh4H1z6aIUbVEf45GDaEla4T6jHtyK4LGi1m2ALw63zwMXMl3OZxzAkFvINLQ/PyBVx
SHx3aAZpAeyNdNlBlzbAkpfsXQaHsVzIpnUx3kQuV41zg7kvYV+puHuV+nWP3t7i9lsVwnzRBJ2G
XrCWI0vgoFhVwfTwUOqSG+2ZYAuEGhMgv38BeHvKaHYShn1KtIMCg7hC5g69wyVVuxIAy5pBbQYA
G/6qHzJY1+W6in3JY/kdhcx82x6G1MFh6nfAzzhGK7TQL/s4zTfQwEUDaWMP7uQhSodQhAvzmeEl
b1hRf20ol1CfszEtq4SUQocSV1PGrn0uJeJHNmLE3C7m4esd9ylbx9PaixK4FgtU5Xs5tOqRRnXQ
dPfUIQXv6Kr3kwx1Ejgnfo2RiczwKNnuY/LP9Bsx/N3IWDjMlA/gwPdD9sW1W1NONaY8ySlllYTt
VQtdJv4sP/GArtX799qICX8NggFhBg+2ZJ8WSNwKUqBJY4d+lViZvw8UFQs/YylTXeqrP3R5KLhy
jrOfNroCDdrTbmIauoZns5MVYDMreu6vNmHB2Zu/zw4brQz8vrnUNeITsInB+B2vNL2cV3g7uUW4
G2gHwFTa4929sxWO5xpytu7h0udVJfGngE7xIuQGqlXKzlJgYkZVL0EZMMJhP8/tz2TbfUmT3lWX
h8OplBPs1ZFodvwK96h4vthdIyx0jVGWZVbXXxlABvRAp7xTwXnduP+rw7iLdVTYbLrF30YmOli8
Twad82V9AUjzyZXJBi0qCpz6cD27wU/e9ZWYDnPP5JnM63Uh4QCWaqWrFvuOtI0uwjMbDDMrwaON
yohpKOxQl0OByf7dRQicu+ma3eAqECzPgDPKMiHFS+QXEh6SW69NpSz9Zy3yePOWO/ybsB4lNioj
slbzQ34mkv7yvEgBc2mDIXlKiwEgC1AHg5zQ6CPrZf1inVeM8EGRxzDfbQPyud+XvSK+LG2XlUew
eNQZSdxDnL0s/ArkiZPU36VrubSG1SzyuvJdJYvL8JlyY4FqjN39gGnR9w0aJt1tcZUIPHQDwdPL
6C2Fbu1ia7DBRPLJOgSKqk6tL2C1+gOWwR0fJW4SVE2/LN8iWVcSYaf+P3sOgNRMhAuyFCU3BGhE
EineJVIRfeJeuoTv+V5SxjpPVoSEQwhBERjLUC7z4GQd0Yu3fepNb5EBuTM2exNG4xBJHbVa6Jab
oDjm6BxIotJNpD3VE0W9TkhEDVXTbX5ynYGLMZ/vUbVBFlQYYC4hRZeGK8Gk9bfjecjAabaa83Ja
QMvBbT3EbEukfPWytwpJPVUv7MsoduunafDzF5qu/Gk8D2vyKKRt7ZrqhUmwRB1hBqrEdjMoXQl8
YpyHSLXGynoHG6y6k5F9nGqkt3fkY1whZc8+R00BZ4CW4vy1KanYr9/TouQ2FOuUuoklsAKAqRHS
faPCvg7g4rjMK+en8rY74dYoM5eXozPdGQ3npZPLPagGfAJzq7wa1wsfa4fkfYfdlJ6Ur2VQaROU
dx1dkIuwBsouE8B/D/5nSYp45S8TtQaqWcZUKuyf7APHkNuBSJdnDnF+FaQEk1KWC5sTiyqSIceI
iM3rRCzuM33R/kk45cx0TDgv/rMnxzFPf7/cpQPzTPCPKlZyr8Ro8KrLmmBZzuS9rxbV0Tv4oXTc
FE212/BQ0Cwiu08ZU9BVGtKb4mF47y+23dteO6DTDq/RXvVx/LNNbijD+u2ZHDpEkzE85xI5+iGp
CM7/nEV1/UU1cIFq5CLIE8cRjs2W/SfDlikndlERWCY0DFeWoFtx9LvNlsRhCYNRN/vcsuesN/Co
4qJ+0Z0hTZwVXC6HDYUdWJOkyqh6VeMN3uT7pjb8Bav/0oaDLfvQ5ZrqMb4L2xBgSlCFaDsz65S4
VQ/nofBXvVKF7Li5TW7A952maUQRxg1LtmISfRQSO9j0MkKUfvom8esPjIVVGhXi7TgTbmWLlnz5
pGG0b9u8louM2nMFm+QVvwKkLohiATT8h33AID5ILjB5uCMjoZkj2W5y232iNauo6DQ48k7VDks5
6rMyQ8V4t3OF19Zs3qwNq6H5fKaODz74DMugeWWMSF2QMyX4o58vPE2YSPDsI7S8TpKGz9XO8wz+
SmusV9lqxqg/dXWTtNvmQB4P1UuQJd7G9zKQc0DK+639YS/e/ZR5qoDPRuk60qPpn8oZ/+mrxktS
bgbJAa98zwJyOFbBFFVZYHlJmFi6zBlNMO/BI17Um6HneuzM9VOdgbBbOhcvsOIJWqQqQzzyFgeV
g2Is2AmGavr0sJOVMK6Q53tN/uj81nCGGutebnUUkSG8jJr4rQrqXBhmNcd7TfN6W0Brwz6ZQs4F
g2TE0oY+xZu1MzothZbdeJIMUNR764Y1pqrKS/fTk9sP/XT/R5fcMhAYX+lQNCVeiz7/H1sD0rDM
PgGfUH0DbzF1d8xVOnw5a58rf7x9C59BBVFNy/MIt1xsdq2IY6I17A4yLM2ratreyZSmLl8F/Vm6
QxeRqlk4KNZ2uwHzGZtVzo3QXJ/Y0H1pShRP11JXzdeBuaB1P2JWu27tB2kWx0b1vifJXBEgvO9/
yL/N3T4Xi6cZkvr8ggCWogScwLYaGOqqyvKKUIonprqn8iM3UL4xa7wlZg8sJWJtPESaHBzh3JL9
/pU9g9g6kGGHMCbyxqW0xeLuqFSAIZCWePxmfbvLMToV67rpVSz4KOA01XhljF7nPckxO5yvQVo5
17wP3gPvb7rOIys3W4LC7EGFd4jj5hRw0QHqe+/IUmPc8TRybel55cAoERVf3/NJWmitVD2fjzaa
isrADnyYzNxGtbpNsfp6v572czK/qqLuNfnXMEtahUD9r8am19tihoKlfbNp0fTvPKTkSASxQdDy
WPUYshwRfGQagnuX7oD/0a6Nyei+HAm45lODUS3BBCbok0QKFrteBppcdEdcjN29YdpH5xpv+pxs
dZcO9P1K51xQgf8gT7sMGAVNMbEaS9sKPY2JPJcAkt1LtfntItzMxForag6flv4LWTHGoFDhcGF2
JaOjekdh7XBHFFkkBPlU+EPg+lIZLfQ0POD4Xu/hBpR99TBHa3BMsdQPbDUCiMXi2edUajya3zoV
5jSppJ8x8kxRvKMGBgI3L9MWqeqwXS6HgXViQaevUlC+FEqOOZEtijLZE3cSkNcf1DEW+JiKwX6b
+UJDeNEJoRvPT6ysNFYhncM81d/G+pRllZZA/Lq3CVlu0YYpnvpvCtRRcsLyA/50Se8AJzIFJ1B5
TRtPmyG5fddt0MtWHbEkI5Yi484OqnmR7dyOzDXzXrve5Yu1wM8fjB862yKC4SPoqY5I9Kt5S/QR
3BbWz+F863dwum/tbVzM+j08ll3Q2lvFyj1YgX65Ooyh6ROGMYK8OeoBcVFHS10OlQLZ1gGUVMyV
5KX2ni8zQ2SxjxcVQE01LYQ8jmc0fizAEr0zxrxDoe6NZAZPbT/eCAYrn1PyyJ+9reqc5CAzFvFm
bPep4P8gxEEx48sLbLMXlZydSpamV2NPLT5H0522N/F7XNRB1W+NSBWdFPc9oTk1UzfCfNsU4NwK
eis3hsYgQvRq8ag+bEPYVzKqx1m0oOfkEKr0MUjILegRN+AWbJwj5eAi6o61NB0B047eiqPykMj6
IA+UxRyotuFI+kwH9OvRf7gRjt6EbTRVt87Dtq+oZsU/4e+GclkeWfPCfNtuLee0WCRY9WnbFQdt
N5RFIE3aQTcW2XXrpA+lvvaDHy9KKqxgHYw1vtCCyHMMM0j6gmUBOtHpd53cRf5eIycq0C1K16UX
3lyrlmfn9iTzQ8hO/LvxODwj1rooGcvkJKcEXZMBiqRRB/cyf9FJN11QQKXuTi7vdSV6t0pV1giF
VA2E3oaKmnRoNO6uZa69peU+ScN/KNjpRxoWwKh8keux2YtAal54oLWz4v1tFIY/CmCks3Q+OXst
9YfSe5f1lwF+aIwRYJv7oFAMc5n2XgJFzi/39peK1Yk6Yx1P2snpfYS2bZa66AeijvDHAfAAp143
vSM8Y51Az45C7m13hlF+NPgljsoxNfs2eLO/Go5aLrwd2AjcTNFU4rQClWJ3SMeJCHRp86lBo30o
4ufIgpMkmEBaDlG/qaTLf0mx8wzIiV+IYxzc4CRVj1nS76WjFROpXKoZlNq/orp6oUuWzvVMxdhk
XPqUcfgfgZ0IPIxsyD6j4SZ29HW8SHTacfP1U1FVJlnm5GBdos2yQiNW4UjG0gbAUxbqwH7VX7p+
7+Ap8fZJrVupVXdjWEaYHRjcWXgdbVPiAR+Mp1yURtmh1pwwSNOAiLqjxqez2cBXqANDQjzDnHDY
shJYriEjYYYQwx8hfN60zFBtieI4VUtqja4Onrg+hxrQ3Kdl2ijQjlPLptTExV6sf/n45WUN3ygF
kyuF6Gbzmm+CnBE/Xp184jImENFj4Iq/9dkc3FsnwreSiLALzxKOQA+0f+WCWVTAvIijn6EytsJe
47GFoy3eXXS32xwquPUSbO4zffwsuU88SNElcRy1PKELlIG4ybTaUmZwz34nRncT9jOYxz0Szh05
tSu8/+JTBaxRI7MvPYFw/HM+AEPwIc2JRdY+grOoEX9efumntA4xS2lCA6qclOrIQuO7KI3WCHV1
I+1TQsiBrtVz/FtO1T9M9sMvEYzGcZTQrI/Olr90iFP7toKiQm7bGoNQOpc9fIa56ApREaCEzDH3
OYQHdtIhUXsr7p20o91ackz6IVEmfL1xze00II283r71dkpM7NV0XmZhi+SF6hHxFh6dqPMmqkV4
AMIlvRgMYGMrGAYgVdTuG6mO2h+Z+IONyjX2a9xl89fXx1fzkH51hdOE1CGVG5WVlniet0ZufkZ2
P7ROwwcaZm2xOLHwhItmQQwPVt3HMi7aMlJP5JuV0hbGp+DqCvDtB2nCKFyV9mmD3xHjOFJCrl18
gRSoKl53pcphymwELdpIC9BvavT4c41SBFkQlZhJAqhLh8I2RlOs6z646Cf2jQwOJUZnHuQ7E0A7
pP+E3/cxOUPa42gm5elyzGpx5inNDB19vTpibi0rLOX3pKt5eipkwiY0PxlgHYA/S5ppkMEWF36A
1pjWnA+iDWf4MCrYgEf6rnAwuDn6jRi+Mm1epKeoqpTgDCIv6giWhm7qqFI9Xx849OHi+ZU/cZ4Q
xxol5lqXzwIynX0wQvD1ueLSsDKDU7raV04CXpjUXMYlTz+ZY7CCW0khguTvIVUlohOxPCY2qTEO
+2hCcyfd2NR8b+vpcB2ETVs4bNBRaYcuzUTWuLjW9gjE8rPPIW37ERZweHyrepk67R1pHjs/LKFe
+2IMpaAQe3o8sY0ywcDpJ6aMLZ7VpsE9wpJ8fk+DywbZNx7RhxBSnSH1m3/wOsmh4BmAV/IgeaOD
7TGABFLQAyA1UTtJdU/JsKNHj3OyXHKXno6v9sQuGsuuH+xElM35mjH2nTqZPZRdCQU5Sp3a0q3D
4HiIvvbP0nl0kJVtqM26nubt8yaZQYNulm3Sty696Qx/1997nF2bx0N5Td8qh2P409dtM5wS5tPt
GBiVKcCG2F8Gb7d70Eq6o0SOuM03s8L/a2Ey62taE9RX+1oWF6X22Ovg8ap+ZRmeTQTIeP2JqIf3
kd4H5QF9gpVjtA93Hz7b3PJd2nv1qM9MN6VyoX+KVx7V2S4YdJet/iWzCQJDe0blM4FrzV9YANJK
4B92CBSL0l0TwzcKV0XX0gDhD4C4+VDadyG7o2LsNRVFYjsmNa1zl8RNA1R86j9PabFI6pvopsgV
Vs/Ow3D05lS5X6LR6GFZ19oLhjST3rLK6KkhEnd9YqDnbwDjCbeji1kHAb1mtD1EbHUoA8KgG9KX
15f4Q3a2ScnsJ/HRFy23bS+C1yot69nKLpTJnbNLrn8eTW0fvIFGw7oOAJyRY3hyA3E1M2YqWNDx
VVUrOjHxW7ortBnhtGvu5cW7LUapN8TSRGb59YpFlM9B475qnZxMtb/uBP5nldrYhwmNPUc+JuPk
zKedVFFyjBF+cxP30XSeoBE14CS0Gd9/gH3u21Mj2rfr/vPbq6ch81+QzEhH48n4FpwknjB5zggn
Co9PPLrPa+9QEYP1dRvkErvwUj9XcsSYQtfamyJdpf2iyF0ObAQHlwWWb5bnwf91yWSm8TTN5YVD
7XFVaxGoxpqzvZjyrHFntWCEQz2hkSTmQ/peRFEZ/lQl9JXpov4ag68uoFRaAoQ2FRyPlTy2Ovli
2KvoaJCOe+9hS5N9i0sQPEtiJrDzZfd4RmRM+lx9ag5+lDG2fv1DEcqEpwWUtoMRT6FZTtCGE76i
gGm6pObdP+Uu60y5urM0m37j874st3fa6o4r1OrCqFTSrx7oWmKG2V1ETg9HRfuylRQn/PRBN9di
Z1GRDElQFfYG6OGsxboyma247D17Vq+HXLbNCGdKwI/tUMx0kWA8ZCv74Q9/ZujkhNVUQns8hXRh
G0yC8ZM7pNAawPTgGxDTEdUWc6+IxRC1xwz7HLaiOXwSDRMupL2WsFfmBnuFGkxv08ZkiaFSZRpG
64l7ms1jEJCln7IMHW/CewIKGP1xFD9bTCCfa1dVetFwomRLPk7M83I6fnLkHy9E56Gv93rh06rN
zp7hdpyrOFEAAjwksevn7Wad/wtVP3GUkJPy5zSYAsPAtFq81PvLysiI7eej5vU/cOoCayw78cfd
6myvp3eCAYqbGZFhUzblTaKqwG1NTbFPyr4QwApm7s8yWsyt+MY2CHSF6kWZVasYNAfU+43319mb
Da2iNjVfCj3gvRftkLfXQh3NDWVx67qSRTTthgkemg/jKbdq5nx9ZxSCmfcnkIHk+yQHpbtICJaR
IWuhRY6WJbeixiZKiukkFNfq+i9IPVcXWtwaIk9FzMKBpy0WmDFqNsSbMDB8Tk4xg0Z9WBklQmIj
Ep4jIthhRvX/cEyfb/3k6620nlmovvgsyJ6ZTMO4MF+KXziirtkgUm15lm8zDNJD4IH5Ey+NzQUf
jZwGf9LBoEG7FIULcFX+rp3AFtxMe3fIJbCdddb+9hifJKlfubMioU754xEzgW6g1LuoYDzpL1CF
cqFQkWocEu3nRXh+jCT8MN04tEpz63V+8ECLHYKCfIgDmghLovMBH8VV2OlBuWfckKb3zAm95l+o
pK36u++ZeGLNNERJPU8n0G8i4AbuWQ4jKpKtE6BAIeFdD/lrLe38kvoVIm1aqdLNdnA56ENd0uhc
MuhYW7zOThx1SVJ0KHHP0ctAehqbeIBAke4WTcbKaCI5EbPP5gjur1iQgI+EWqzmyqgJNU0/xfX0
v6VhknLWMy8/cYBNTGFQQEX4zJm/4VOmedNl/OLnekQ6Qzk/Xoi+8JkR/zbi3hRZbQlgdjWqAbCU
kg+UwWalPoyfQupcIv6ukIUUlsINCt2geFlFhYGH90T4sybdOT6E9EaOe08Qab3tuHt40xMuwK1C
psdbPetv4pS7/v7qrLSQIxVc5n+4GhfgglGMOfRn1cMGEoC4nFb1yXpfIJRH7eLxoSmDz+c7U4vw
0Xe5GuJBwxqTDT6KnLYMzeeitX7nwNn0co7CGxZCRFl00C/MBxvhnJCokqWi2su92YhuR7RMQ/Lf
K1pU8EmkIjDcQ+B3SKp+Zcsrw/fXX/OSrKJfBKXUsSjY7J17ezpeFkTdUmJ87P5qywTRAFdd1ynU
Y+9EKFtlkzpWI2qK+g9/sYJm2rWS63LV8AI3SbxyobdHKKCrr1Of9HPXLdiH5a2HkqJfEHzLoQFo
FWeEjqxzEcYlqcRb/f6p4vDTKShrzV1gr43aS6JMxY9+SwAbXsh2130/175sZ5p0rbFr2jibsvxH
P0GyRusTHSN3v4J05vQoivfR7cle96gfB5HV5kNCZtE0roBiiTz2Gcu4s4vSOYnRJbXxgZ+TQqxj
L927Z6rJqjqSKhlur45XvHTiEaRWvP5pOuOSO/rDBqPnfoCo9P9qr/i5De+IAvqQRAL46htiOIzY
LMJXT8v4KwMeVArLGrbFIIxTIbpKijcHy3Wvn079u4lT2uDE5uz+Z3taraWOgsjNUmEJ5Wud45al
f0EVCQYkBk+8NyUOG2nWVAxHUU9QEc/lmfjM+g6b17eOpKX5VG7UEbl55Ep2IZlfX80GhbHj9v/k
LG0AeDY1tlFr/PFh5hYdSm14NyuUpR0nQ+snkje4D7gUAcwJx9q5+S8rU1UnkUtEWPS3corTt7cY
cCo2sHyYiyPoVpAkjn7FhaVR4mUeq4432GJvy69YTbGKg+gLVB0l5orunN3QDGhhSOaQ3+QY7wZ2
9TTwjntPATX3xD1wnp1jYbrP/GeeEasa9x2c1WVaV1K5k9Kax7l+MXqQ+fA3c6nF2otuxy/KHb1u
XztPTDQG4R/ikTdsfR1Ok2KiraJLfcXxeQXpyNOfSR+N7PHbYB/NdCGNPnGsXzvTjZsRWfRK81Co
DinA31sgJlWuNNj8J+UDuFKBc3R08l0Vtr7we1Zaod2bcKz8ZTfZZiIyEcQjpfzaxb4GSsaQPXQC
XkHzpwu8ww65o4Xg3Fn8i+GFrqwtC6YFUBz/d6hYQtuGZPNvnd+p/Lc8kSFHmXUAyJ6Fxb0cy+6d
KL2KIrlKaakWmbBXaAY/KJ5UQYMEkOurnf9B+DOrdMF+ozjLnkUo5rIhdvtWtzkYy+k27rF4YjkC
YPBPDHU+t4jkjVIAdPWInxIKtvXWc+o46aLCBwKl94MIoqgvi6aNQNBwpj0ObQmaMuXn+Ax4OSpi
dwrmMGLiWE9N5bvEQg+6qzYwb1ndqY7XKgIQfY33nlz54iJN4EabvRlK5O6UWv0/KbEqpu1sl53g
3I65UOJ4B+oobrbo4pnbgfoHv0FPkH5QyvEqDVtvDOGA8CM/lBiYzf7g6I0DyoX9M+WOABN7jLRm
h/SQrlJ8L9AjyAeZ7Q0daYOXhpuO/GrsdrSLVx/PNZsfW6vaDWBGl9hcprrVv5R5AxiC14BFHpsg
hdwUOEoqrz94jQA0dh/Jw1CsckIU3EMzQsCopy+JKgNDdtQyoof0bWB7NMTeYDVTsJzLmqPRMktF
3e6gT4PbkUnGtMvUVDhP2k5ajM7yspQPmoHdh3p0kuv84spO1TnuFW0kdeMjNG5iMmpZ0IHO/Ddw
Lwq8e7/1jl6gKrdBaIOomN//7cONIS/CTE/sJAV+tuPt2HZyCOZnI69AX25D477fHm9WwvQAWKHI
wy0lb0fiAjRvqBkfwyviReySLZ+IY1kwK6oQQzoNBB9HBWgRb1Iab7cuY7DgItf+y+guhFn2JCGX
wrs4j6+Ky833tc4P1DUSM+jxl38N19BN25ypGO0KpB2JAWbm9wRdLWkIqN2KoFoMvld9Us6HwmDN
kmXBhZIcvALLHCE7LaODfTvkb7M2K41J6cf2rv6gtgqNXjiRV+rRgTm8JdGb8qCFfSeuMcumorWR
e9ohcl+TMnLaes6Tvm+oqXZzt89Us/8n17I7kaQyoVEwEnqjDjCF5D4UsHLbtSVGHaao+9f3r3oO
p0+uJ7GczEJPnjVcRsTE/G3YCNgfnYm6h6ysu5Gc01A/Zj67noxytBXD5sNCkB+RhKOuAthWeC0L
4+SshxNgK+NpEgntopX9LNoz/s0S1z1H6tbe+ecPJKGZz2mz9RfAMRwzxZjMB3TEjMG+Q5tQKVKz
srhfTS59hJgGmojp9lSnIWpTVrfZuOjQj3vX1xAB7irWLWsCMIJoPY41KdGX2FPp6koLF4fU8SW+
t7kraydXlyokQZhuZDaH5vfgW4qyYMuHEPQwmVTU+zpMPh4EBTIuGTcLtMgw7XHD+CHtXbO3bjgL
nVhlQ7oadC6d1VVb+LPLoYvbS03XFNs2b/3+b5BgedMnN+jAt66VLzmayXFy/aey9iMOsJXH00vY
47faovqy6tVjXB9bpx0Qw4ex5et8vB2faNayztmi5sueUjFwptL2fl46+g3KIl25MZAdLKJh1NU9
quwf5Ddv/4nymGy/Ai1pHKPy0BpEs/MhhoqtZTsQGwrLkvd71/LyyeR4pXOUSjyNCu1QJtoTAcY0
6Lw06BAAbE1CWVyS+TliJ2Rnh8wmm7/MaZwOzPEHLad2ToJ7+EOkddtfCkHEKQB+aTjpEAgwiwlr
l+l3XGp40JiMFkdCR84qaX4BlcLtySR1nLk/MTvFoWU5ZTm8DE+E1/ui/O16y4Gsn1szDNDD5HqL
fN63PlO+7njYW2PtU2BQ7Rw/wUogo80UzUISTXYWZaJQjPUtMesgEL9pfni/BNan0MYuJJcJ7Q3w
sJeLMpHCv0oG6VtrNzlmurcbmQJYgJQs/t2FvoqwcCakF88y+2K+v0O+7VMsElcbTabFWaCP+Mwd
iBWoVFtUHoLzABi2Q4OUL6tN7tO1WSrNyiwmZhyl4SQrAN86jCQdIX43jgfCmntFjqaQKY9GV6Jn
+4jwPKCGdPPtHUbGA9Hh7v0WOvzBe04M8axVsDI2XjQW9NyG3ZqkPXb8CUV2KH56pxhGI9UFqo0U
E/tOu9ZgLJyGwEBsLZ7WYzz+0ybRcVWjEYRioeY8uCdRQgk31QnKVHzI30KrDqglWZHWopzMNPPN
KAQvZISbFLDlv2P8/Gep4lDCxkxxGV2V4BoKwY97d3GlK6U93B3mGkawMvRIaHAdwsi8Ilh5Zumo
H36paMqvUw8PAn9+G4MYdRTAX4l8a3V9Zw59RfGMuxNQyt32JzaM8BNSfEhwFkUbl0eoouTjk5ql
EqcMfIJygMGxSHxttk+ZPmdeAWwBmtAk/jn5iYNheO7zlMcol0KIZw5QfW97KdKqURpAzfAV7VQT
yBBM14iXNeeLFaI0i4+ZBaOg3K/pORX0RNBaAK2oGsXk5lIVF4L+4NbsqhRx7gGqABDsYFcndvOz
dyHz6yiC67jpx3t7Mc3t/ZRm8UAwu6Q/kDYrslsa/0fK5dZFMCz1Tn3ljnSkQPvCKxuvTgN9K3ss
ubmHuaWlrwNpEB8SYDEeSQXl76FLBfhzFo8zU4RP3JcWg2Q/UBChS9NvRz+l3XHvOvD59pTuCrlM
AlLYjpDKKK+Ae1+Se66f/Lk6Rn4bQsG7xZp66CJDIdU0S/gCQhaENWHJPXgijq0YRBfx57PL/A72
FAwpuhKZbZZEZ2LWrIVVGR1Xxl6dj2I2Nad9bqxeP+16jioMex7q1JYmsGUQkLKbvFsxAknW5PCK
PU2H4osOp3u9qDxBld/Xw631xg67IfmHSNfbxOx9HBYlHYML3195rZ5AQsLHqbFR/KS5hh7sIBIp
lHTUxX0eSZG+aEuVF24awQ7K6PoI95y0qErqvWNwrSv0azqXdlo3ltX9/65llupq1iEN6cLtdQjD
NueX1JNk/5xU+SHIvr/rGfXt4GsgKl2MUhyJrqajRc9FfvHt4pwoeq0fBcnDiJxbGfNHpUDZwhYM
5yPJ4Vn012mOcHWvrLc2j97s2nQInkvxjPdEyPIAGuDOzX1jbD/tS+OoDmxjexlKb+uZLvqyOqq5
xneYxy8uSgIxFZ97/9K9Fm9bAuyiNgYZbB07C9cUueU7tbB97vvcFGjpWn0uySUXkNPjPv73hk2v
sV1razvozplCrT6+GzVk8fmosoD4MUC1P7qkKI8swPE+Z37zxfV2zrZ2TmuQRzED9UTzXQ/WyzU+
czK3mtwKpZXYiX4SNtOAmHmKlJTl/238Xa9AD8QaqABBiBx7E4i9TOSEnTSuoC485pNC3UZc79SN
WEceUUPVHriFk74J4Tvej7Qdy7edQSwwfR1HZIpLsZEayw2oj4hLqfLxrVvGMoNU6u1aETRQnWf/
MEJwLJO4TmGjPFMaXTHzLVDzP+fJFZ13uT8RRBhxtBclkAKGbIVACBwIZnXHHEgN2iGUQj9vRb/l
ROTjcbU/lAvoEmGDqFi5wQizD5fHZb+i09dwNcVYla6gpENWCMtapwusS9uaAvAwz18OnPTUwjCq
ae2V7HbBPhp8k24SFGAo42JMMGQgDoG2B5ZxStAo6LNpCzpB4BGVX8CapZfSVgl1EFJ+jAGPrZV/
u2u2giJByjvDdsyD0GWtqD1vdnrL+ws+GtpvaAi7uD7VOvI0jevZqxAWHJ7izv/vgXZQD09MIWwe
Wz8qF7d2132J1rzC5/n/ZE9QHrHt6RWvw1MlE1LSZZleskMWivLFB6puXNzVaxSymxuJWzFIyLQc
CMChoAxHIMsCEelb+u7eEqiv3eW3myeeO6UgwwU9W+lLwnYSKfp+0Tni4BtELclpCj8LVWuQjPe0
yheUrrdvXASrnEO5pmxOGdqSMgkUs3z8EJY4RUfmHQQFE41yoAjxmq0BAaVqsqgt3aL3t47eLiTO
5X5m3JUSKSY2ZHjsjL749tFi0sK+NhQuf8ekUQvdPvf7FRaK/22NK/4l7eNqdjQzFH5NMXxCif74
/5p/ox8cWmbx9QQGc4feMZcPEWN8cLsunAor4bX9/weO8wrt5skC3HdYr/iz1gP5ttNVmZcX/E5l
gqOKIACLswmMgO0CzzVhfMWqU/uAYwjCSNQWRERIhZC8d9q7FHA31pfl13f2EyyD5LvpgeBolzdj
Zc4nZd9q6xBg7/9EmFiuj35LCKByqGqthO3QUnYNrOGXWgDr2HJfP219d4LSsTIp8Su+8tRwGEtH
MeMxzs8FM/4uXKekNyZBBs59FCoSQXdXEa3sD2lE2sDpN0JgM5FIg9+XHUr0x+HPfMvfPsAqAeLI
2l9G/iaD+eVHvU0x2mV+3O4aCHlszOPv9fPQj/I746/INyd7k7AUuTU5c8036IIfTI4Zz1ZHYDO/
oF3mxxBSKPMeswTEyPJfGE1aGG7Ld5ZSbGVrfHWbFU5FzdxG/4LTBuaJByw17Oyw1cmodARyObEh
Rmzy22BPKlDnxCfNyeletYL7q/7fb3ByRQN+DjqV/wrLS08o1m0Ws+vLcl5ulpFnoGxfhXsItnwJ
C+1cxHDLrwkfdBMI6tLyv9Q/RfgknLpcIhvXntzVQnf1hUULo/kabM8CU7DpK2kF696szxg9qBRU
bSxOY3r+NqhZp6ZSvCdjcfRfM2R0k05t+etJs5wiaW9Cu27z9SOFbiL+qhnhmVf/FioKCmpyOzDL
BQ58WfPI8GHFSE221toCwpV+/vfFEx5EzyshxZl7bhdqA8ZIIhzuwjz0Qr18kF2G30EuBpCbd8+S
V0E6dvUxrBz6ZROyZKX+rYTZaBoWLdRsJcEJlNHICIkbg0s/qpGP/hkDJyVh2HDWuUY8MgowGoVg
P4f7EpCrX4PZ/9mltB65jiJcOFX6yyrORYwhNFyHIAyBuQ9GiDgX5qlX0/QNOEW5EMWPR4AjjaMJ
vDL5lKerLlT0EMr2E21g9seYPh+b48kInyjSNSlXi3+ODDX48fIWDhEVmfFpvEY7GjRC7p1wZxWh
eQ8UmMT42b+lXgXJzeGaOVZ1EvRug3/TMh6bqaHAjTLKJjxiv6vSjVmZkcqL/zws7U59oyUSwzqR
CEZwANpf9cBxztkGNGTB+IVSXbyhCsgE+MPmLCjkA/X4yeYQXvlMFnq/EIUz9pTuaKyPeJPi79CG
gsEPJsS/Y9BOnd80eLe8mluDIJKjbVKOc1mDzFcnuzc9LeruFSJa/kkpeOyV9Eayd8rHzPO1ULtg
330cFs0yWKdFoYTQY3KKweixCzmDu49qBTMGjobLIHTdJzLAcdigttDpSVLYac3zv3g5avYP+EEG
37PzXEHhG9p1ynaiCUKl8mrR9Zi3FXTYpclLbphzyXi7e4citbUGwACo2JGDTxs2bI5TpNBRDnof
P29WUskuZRrJIZlY8lAdzwmYEIUQd+Ko8SRDXybqEXjEFifg1p5yPPO0eW5RMMri/tcOKeY2ToB0
buJXlI0eizQLd18RWzYGHusDn6hmrLHoG7k7n9ziF1z2+bVZbG30K/XJsqRFHXwB/F0x/0GwHCmM
+zc37IdP8ihOVeUohOj4DmWAQ8Jv8/AYvS1G9w94gG5NloQ/q4d9eoqqmhvXDsFXuZG0adIc5Vnm
AWuQTxiaraQgCi79vntH65wLdoTIwTJmK7gpzPwDQkw+w6QY4EH/2UZNKueSFOJX2NqFbBFVw4N7
aUHdoib2UvUpCG4Ip1EF6IayzyXixUZ1SUVqcRtVSBm02fMLMdsqILj7HKZTZ3McUI22osZS/Yhy
P0Gc3/QGX08Lt8h6pD1jpZG8dY9HutyO8WDIC1zgZTQUCYDYwJD3PCsCE+D0t3JDiDFfQALRgsnz
nRarB9OCwfGn7qdwlbkMhz5ZaoWktJSisunVlvkzUvXMfKsNTpShGP07rCVZlF0SQMEfZMqGtQFp
Qqeo7gTLNJBKDMmt76h0q8hbjMG3+UYqWaaNNTMFKHBoL95NRd2PXY9GxMQcX0AjXvTOgKs35AR5
jyVQoo1DGzMZYgj6gFxngGxhmxjTYN88kBzykWxibOu7ScZdV+MoWQrLynrqNer9Tf7hptFV/99/
NAHaA/jziNOXd/5gWtKn0YRec9GegJC7C0WVybymrzAtUzPryEVTCbpBRMfC+g36q/bXoH2Ll5Jz
D/uRfarnQkeGy/8bIRq7zhqjPKzQtB3TYxVeTzmjBEZBnh6RdXxLzzvYJMZARX7eZnZR+8XvF0af
3ZCe+vY/vV59Z77bhzATikxgxr+BEkBTjQnR1/v6hAnA+jR0GpXLpQKKidoV4XKOBNU+/qKua16J
u+kDurJ3szQYcFmSsqzf1X2Fy1x7+RqWN3ZG0ALsvoSgCUaCH61+exiapuSWt9+7GfWYdZpp3w9v
tcT+xIOAeK9xZ6V9t1ZCMNpa1hsjbSWNBhy3oYJANrZMjn9w+snDZ0Aq5AefeRccv0IZGZ0P2ULf
zeiUmXv95SnO9LmpgHLMHHoSgb38wc9kTKlm8ZxgmUvmK1plplhoT/jWZR+BJNlxrsz22TGuiy8t
et4ANiRWtoQRHHxMeNG05DPhJis5acBeqsX0GVEh8hdrhE688KVSa8v2F4Dqhv9h2PVecj0oBsv6
WnUKviJwM6lFiJjm0p9u8v3F/tq8PcQSwkt5udqYBt11WYuSGOGfUmjIdUOs2VgjSGspBnMuniRx
0mIB5rlAsZdQmjPYQ9ygkZP/eLHIVZ0Cd4fx5jgQV7VCtYe7wCkBS9Tk6Cu3EyblF8K9Vo2gFx22
jDi8T665dblVMwSncPvQHNgwsqD7xrxl/h2t4QsGwytb0bfELBAjEzE7UuaBVOFrhKHhx/pRjpI1
zSYgGa0zmxi5gsTrCk6Nylq3gFidZ7y39OOaN6Kot9DUPCiGmeKiS1Le+rUxKcc9cLOUWwa7DxwP
mxOla8fTWwLONEJ2/y/NOt3sDL19X1MeiS6rMbNqdPlbalD2e/VPQayf9pT89Nlcgjibh8+6Qe9A
URTlLoRGve2SOi1KkSM6+YaJsF0VpGR34qnUch17NtIrF3rZJ5v5wuHU3YOFIFKHG37sGwtrwTDj
3tOh5pdNKaiHQCI+UGIiHlcg6gfFGjnVcEJpFs598v0fW5h2fR4/y00pUciL9FPXZinT6DHFhthb
KUDGUrCyi5G7md4gYG9DxwaBISTQkOE8o7hOv9a1L4BCbDAoowNe1dFHVYHjlI+kp06LRGETVt/U
QVO7Bn10nCsnJSQyTIiPjvRTaPFGr8gjV7Ct1BevztM9J/4Fm4V1PBFbLO8ohxf1aP4wIjhRFpiU
WZtl8+rmOVFHyc9yAWkIYvSnlqpmBFwzyrs9tUbtf4hrk3OCo6axBxIVz7So+aNaXvkggYIMOs93
msNFnIeygGR+OuyjysU4EwpS777whvuT+ito7WsPFgMXv3psPqjKroL0//fiZqD/7kVpxevBl8FK
kBhGmB1cgEr7FpgYbSxKOIQpzNHDPxqa4JiCEtQ5ruRoRqlHSBdes2K0Vbz3nOoFisWiUHV+P6DY
qvh0TeoM7OYInSyhVpXoqUszDg3gyf9Sz2OjuUUJS3fjPVEoj8R4QNwc/+GMGZZIav2fF9i00NXj
yvKpxyKaBG0+pFeYvTVh1zDQbq0fs87dHts+6Fl9yCEskQBQ1q1+TfhW97iyBNV3OL59FVOgamPz
Zojh0eKzHyDXobHm4cJczJCGickgPfzB9dIqGN8YwIePL2j2Gpt03L8r70O7hZZjmDNSQqMtARGc
33VHpZGutao/bWhCLBthM1bye0oVcfbBr6uHJmbcFBVHDv+aavzWv+RmcLs897v2eOT+5lgdwo+/
thgj57VZ+lAxFqMTikPEpbMTejDzq49pW9My0ecKffDfvniHuEh/rQirskR6E06VN3Vm1xyXBKn/
68jv7s26dmleqrtETuNsWF/ciKWJDr4y+a/f6C2PxhgTuxVj7unXIVV+urX3YsmAVRsQd7asWJDR
GkNtI9TfKcP8FUvbOOVNHX0IXcrxEM9gaGiFH6X/4YXA3Chyu/6YS0w5G1QLFdyfWihl4ltpII3c
n/8IqKC6T4qlEUS9obHrI5Yu5TsJXdrffp4lKU2jx1PfKB3wt52nY9QzCORHAlBAqQQcdF2yuL11
rY2OqzJ6KHlL2Aun0ztN5tKJKn6hi4BsUAn0WeSeny2aBCip14ZGtihj/YxkxiI6bx8eEO99xcgE
xW0wN4yxXkqql9G2eI+K99Su12K0E5zk9yhC92DjB1HUv5rbQqlnvwDQcEE7h7Pf+IPzFpM9Z5lb
Z9iZ5aeEKs+aUBuy70OYlofax5FWPpPN14Hs/d1ecL3/SNq7Ge6AoNBlXjUPdsa1KJkZOV741uE+
3iBKDi82rrTB1AK1A+gSI6//UkX30l8r2f5lC/E2qOvMLepfWqo7X4djX4YRATo68zJK0e8ixpEz
N7NW9lND/31+3/CUZG2MBNe5JF4QT0qBl95H1DDAPmMKQSG8MIztvv6w1LNEOVFd7/EsFft4mRd2
OpxiB0Qcka/2BlUoZdkvHO7/tgbn/LsTpdZkg69msn9AnGEGXQiBTgOYA2ce7lu7bwI4BG/4VffY
r8l1hqHKZHggb6kV13WY6Ki4/Y0v4exbPk1IBINUD1NrIWhBdDYFsZGLyAJJ13OYErC6a1BpDvCJ
5wSuGvnv2pslVyySwLSXD8pTrTWx5RcEBdT693Ozj+ia800J/VnwWO6oOtevDe32CxtIkJ+1h9Ed
bzcqvYzBDS9Dl098plOiCc66cPMg37AUdbqq9agMuAUf9bHtiH5HF03fItZh/L9PnRxZMiOuKohJ
gJVAnBLhvLajAuKZ1crReFE4Qk3uflBQuCt0FaslnFPKNr/K2erT4qZaAz/dNk8wJG3r95REQ6Ed
9lJDIy2XddCbPj+ICh0b8eyp4nHr/J8hOr742vxNXryM8ambaoa1s423gincLMqPS8okW1O02YTa
LDIh0ZH5Vmh/eqKz2XbBWCYEU2p4c8tq89kBBLAnJNsO48y9exW3GRDcVmywTc3m+QXoMmdCBSQs
sE6228963U65wnTx3SqltK/t8YgHa1jEqQne8jNr4sgnqPFFWcg9T1WbcWroFpsEUM5vrHlskmco
Fu+LtSkxPRpwP077HsPQJIUZXRClROg8muNhKK7+LezXMT2kepdyiNv3xkWF53lVWBuQC8xk2Pm2
6L4WLH0uMPeiyn409yOdnpjrxzbkflo4WBJ7yRemAVEojcbyt4nNKJHrZi6o0WRGAIouxMtKF1yE
O7RJLkXwaFdVB9eECCYDnK41DX9GZPIDEsZ4reyNYEYRHpxdVqn0sHJETCSZoPF1R6YArLm4tqLk
WpWX4UjthzPmgNf8htXxzY+BQdO+0LHoh0JAmH+9cp6Yzmf7HjnOWZjzCx1+xtcoG5jSFqsC1fdL
iPHyYA1n8lzp5FeZFzB8Au+hQFV6uiA+4lYGZxE6gWetDQYr1xsybf0WOsZUCWChzoop+Jce6jQ7
DP+ye5YC+R0MEnTsKfxuXZHWQgr/FlRBTRGsIwK77zIXRmEZQyry/2bDEAj7Cau2OlWyHovpe1EY
ppd3ZEvqzov0K+FSuOP1RWrEdLkCwuzsS6UQsZIWB+ckJ/0vZ+TGqTvRoO9nTPZMsTyQj91o5o2g
gS8OfEFPt44Qqb9tZH3zteuXk+lOXAUCN724lT69m4ymBu2LvYwmQNEX2c5LvzbVSjZfkzX5huIi
EhLrJsWzoVlhlI1cFT0HfgV8mpB8Ae4Gcy1dYhlyyNUnxOmAHe4AhjrHcWislY0XUFfI79WRr3DM
BS1FN+innbCY1offfZ49SJFk1M62T+9rK87cmRa+mKyxchnWt14qRbhJRKhmNppj/cDkHH0qwN8w
r2vla1OWPj+DxJxwoXcS0XkpyyGdlX2sBqv240OaN9eWOFLNl0oUswtVy9Ne44NJXwx0Qa7TcNA3
DzdzNU5LT/jWwI9ORhZmkpcGU1Kzg7F6k4RnHUL8Hx8bWlfmRcrJs/qNnjfR7wdeRTwiFlhksWkG
xiIfWoWuTgtCRGwx0W4zEhd6hvKyd9tu4XYNdNx9q6oADCL6GVdTMifsV+xynP7o3CRtB1cTsuq+
HpARoYcu7e7HyzcxJPWWYAe49k2DN7K8seJEv2RfIei6SptbZGqlcLIx7Qt3gweuDQqNxU9vxvJb
o02p66VAEE0gx68KpbqbLeOhMVIejqAE/FdtK6vkR2IM03seJBbBtgmDGoH0wpVaA2EH8VPCI1hR
8bOJL6AJY5nHkAAxiwz8SEQr8ZRUB+dFMBVWWArHTdR6RUpuiMZMd5BfPtxtl+paNIXc7rSdNMt/
U2e2SOYNLPdJr00nSbMrDqShVcHI3u4NUDM40GE7GOcLvzKyO8LcOjzWtoUTU+1MU2zb9QscfvlL
9GuXfhJpbvCsZeplNMXQrjz3gq92mbV7oaHqQp4MrrGCkHT1peiqZXXK/poMh1z1tv0oB3oN+n8R
THlQkxxfJ2V8+j72t7+XKZntb6jiRm6e1z7vXIPfcAuf99PbHrOfebwozmUa+U0q9QUkkRUyVOM0
Yyb/YQiZb/8MZm7kVgm6oFfhL0ICnhQC01lg1P2VU++ThTRRLRBq1Ov3Qr9EWWM5rZKlAD/0nHy9
F+eKDdDWvKW7z683697pIzTxi3CE6uxYt1a0YDMJ4rC5rVoxgx0Quqdwa0mnAZP2Iwrdm3E7JMFJ
ZWzI7qjYhROyKHSJKizPmHghsLaNPjfPl7i6DVsa1GO+KdNY3YAe3IB3LvPmh6IxpsX9hsdQXy8V
iGCblQ6WPLlqq45yRcCSgN1QkQZYCiZtRayhQpCdSCpKThF8mYG4aEi+OdvsbNNA6eaOFjwVfyYd
zY92LmAr1nCIRdYVyQWgchnL8QeYSOVM+xEQyL29VLeqoZumvx+mj4Hxx6ddmboNpL7HcHsc5WgP
ILK0IAHXXBVOUP2bZwfR/6lxZPR2tQCKH3EF5bCHzRG1ZYoFGxzmVAw10ag63B0ckl7eliO6NjGs
P4BOws1Atb7otn+dA7laZR63O3HDhuXN1ouNNsgm4O/gW56iinKT05OOYBpDGXcpYipDiFc2U8ii
sAGnbsW3GEYdWPu4ioW8DtIfNl4EocuqbOlEr3Z4L+5+l1Q60B0gaLns4PfDmKA8sPU4bkQwjcbD
UU2wKm7MwVeph2EZVuo/H8xLNqxrRw4fg87JviMXINdXeGNPQoJGtGdXjp+WNS3//5z9/XIg7Cmu
9UBRc1exoz4rrHkEm2XZIeh6Hw1O8C8t1RBgNfnWIUL3eDhOiCPd0CsALOYd1iQlizqDx9+mzk/D
DSWYfoRha1xG+0p+oqoYXaxvwqxKDM183grbiZxgTQFh0o9VFxIBq7lw085RFOUcUs4YHxASmZeX
3cuV8EhD8n6QNnqUCn/tslMJX1qdPBHyzClTE4EdCfZ0ZNGrkxanOL9/YDNPUO6Aia4WhsfJPa4A
BDOGhj7SLp4aUrbPZQXz9bmpkKaz+R9jQNqyP97LIcPJkosEX11SSOmLRy6F4fRCcfth1ZPqnJ3V
zGSS6ho01JacnqtW61X4QwrHpVpwAvRzdJZ17TM9vwNz4yYgfFpoD+A7AxrIbw85zrOaCYy7Bsvw
dlN+X/z4CoVE2wxW2tmeJV34ArDoRn+K0mIkFNo9U4CjIqy3WYhIB41el1kgbwECjfd6BQT18i6H
r8Zo+ncH/X5sVcAm4fOZW+J2hFvMa1veiyrwXuKGLATM1Uibt9BBBMEcHpUQe1KDUHCdwcIOLc4u
EhK75s4k+fdaPwyaeAGNPKeSd31r9/W+LrAB7ONg7qzkE+nmoPTeswpJSRIl1xPWBMnuoKmOC+cr
vgxbm65bvdB4HnBVvjd/x6Qlk0Qo1z3vzDPieSs4ttS5OVLlVMVwHtEicLRdzhhqKqIZ3kKLnk4J
Vx9z/v8DEx9ckbuupS27KuEwudiiZ3xGa/wdZV00kw5oKQhwcrKxHnUgq+9Wi4pCFo61ZHQ78Tpq
vpFWerWwddK74Ok6N9YRsslYRkiE55fjW/4tPVWjjHXge616qVJil22QdebpBPMZ3AMEbqNyB0E3
zHHuObwZhd2FjHzDIJ0ytjtoOk0fDuGWWpVMTzT4ATvWogwp6hWzEaQLJpmJ6neVbgLzNx5PrWVe
Lj290fJUR7QXZWaNQqaE7gsxFFDZExlw0NIYJ6MqjWvYvc63oz//2CXKE9cu8HLEIrRHeqfPfow/
X+wVzEtSDSG2cHcLpLPAbHYJCTkz8Gg0itqIoKmQ16zsdG+iQkXcCeMBMnjQh+bQzLk6VkO8AdNq
D3GtL6/o9PmrR6N8i9h7/SOO+t8LuyxCWYOaObQj46ErPrV+bOMkZZdKscUN9fklYlejXvjXQKUn
1jqPVjQONizYlM3/G+uo5kF1V9zmPRuYWtuAXY0yWwKTjGEI3xMr5m5/GbEK89l08n1gNtDCQWgs
XUADKpsyy9ppFy4G2zHKv0zahsQ9P8PsxMOe1D/mJRsU4rjsYIXdMItrnbVUlinNwTlmOmZdgYs5
nNA1eJiY3fNdMXPBjWcASzl3qMQB4jnc+Uyqo6LT49tDW3gEjNaj/xFMoKYH1yfDzbQbznkWUJGu
nvpTJI8HHocjz6WVsoAabRL+UCw5CA4iHn1WeMVWCXwpSx9ay5quHTjAtyhtxzszNUrsOvhOQJwY
KHVR5OEiGr2u1tWdDMwi4JnoyImz23U5HwthxLxtPlTyEVWPJEreVJ+WyK66wTgu0t34z+yujhcO
eD2qQxrSu1cJ84cll0VIOicvrR2xfdmbB29iOE/QzJYtb25weY7KJF7dxTe5SNIuhqkmBIZOCILB
tIUnrcTIGVo+JaH3y+Ncn6qHBLwi9nSUzQP1Rdu9CpdrnVWvM7wugp+DKmLMKWM0fhEYUZfYdPLg
lUpmW2UcPXWCFg8xXnOnWXWR6COyjYsWbNv14qu8xDtic//Eqk7tpOnqUFKM2F3zdviTj/w5mhDG
Vbw1LgmI3OeTs3AfJ7GoGRgkDUe56PC2NKj9byin2E6xFGXu7xBzT7ylFjy6DqX2sXrffGsqeshC
owJ31+APuW4IzOEafHEvObkTi2c9JBeJpN9eAKOnWpRW0KYgqV+XCtw/1ehi0CAKjjCVwbvILyVA
o3SOEs4Ty2sG/UY11v+Fql+c2TYr4vj0HfTki0JVI51rAhl+kiaIrjGhLvlekW2IERsNqQW4BYCg
Hlbx8sWyDsveZUYOIVx63kdhvsSsQSlrX/lK/3zL4oqjeN6oB5dXSIkXp82k/yieiYSmDqp4gXGn
NYGYmsKZdUsNYb08uIWg2Q7x8XGN3cmFxBvNX2pSvoyXdHsfpjOOLxAYwyt2aKSYRHEtVMEBoAgO
VdeDKacTmu/iNjA9RngUeO3xzifxhrEL62bHpPdaCHNrh9aKcXavyyVh/Jvh6wYfyuNgrPc0mfYL
D0ie8dM4J9kasp0SRqQAcBKjAZIvZYvcpouaDzjcBkrQbKscYR5+Oo2HAVXIVhZGL441SqAOxWXU
RHf7px3vXtn9fFNIRIZUPCTICr6B49mUVnK5yY4VSScU8wRgv6xw7jLjDOK8VF1Jogr6QEuAW7eh
tn2Qg8wpVcs6y635+7qwpFSWa7IiQ9pv0HtjzqavYqnHlXb8lVHUqGR5ThGtJqbCk+1bpFK2V1V0
ffq6zfLG0/3yPeGVo+YrZ3CAF7WKJDJ2hLOuBo+S2AvNZF8t8mZt6TNRjab/GgS9YkCHe8pRgj3V
ViAg1Ywo7w8/JkgI9hewN7pgrKij2ROjW1X7yXAke/Clm9tG/hbiRfzEA6ROb7N+lgJC7vtmY+Dq
NPEdWFbW1NiYALBbjiqy09eDzQxQ1qeHdn+GybyHHNZS0hTyrJNHolZ/k1ekdJjWGy8OXYnYHEI7
WcQn/mO1TKF5fTMrivh5B1nAWsa45bS9KMDawI7cqhW4DWHxi5QxHqrvm83vbwxY+8lTN1/z1eYJ
CKvoUkq0eSjHrEktfzUvhmoX2UulSauTLA1w2cjTiOuYTOtUcpo5jn6cGYtdkn2AltYhnZyq1J1o
iCfYgngBzFyaSqBqfCrehkeGWEzmCWAMOzavbA3A70O2X3vyJnuC/JsvLahQ/2KdhCIio/E9shBv
ZefF3+y0ltLsmdbD4CEbWcuSQCqnmEhGQN4pr35BULcxW3zE/9DPiZYS3Am5R/7GsBgdvnYlflJt
1BWEAh0Mz2a+bONxLjHtfIyI0Ettp8mxqKSYdHz0bM900/jqAHvZbDqC67Vun9waWzU7XQCxV9GI
y0XgOipsYDqs6US5TCk4dPvlvxZw+0DF4V+uPfWqYDQql4L9R7eTRcF/AsjuPxEKmqSIbbfHiJn5
4bQ4JI8wywN+We/3DRNuQNg8/U7Z49zk7JhQSUUCYO5p05Ki+bVpn1zU1dFe94uODHVtI6y2BG2q
jkQIiVNvHS5G6r8dIY+jS+ehXWMwzM6vkYOZLwBYl8gmWBqPJ2BS46GgyGceIkj79Io6BwtMMnTl
+8Ur28/GtebQ2zHbc5EU1c6WfWO6dwFwK8KrelJNh1G0O8BKv0J6hhjXzSoVj4UCeG6HVq5f/SEL
ITjs5Mj7C96oHLqs/N8KH/27UHHQNdYvXPtcmJLV4EckjpqvtsGTBXl7+LdrsErtZSEJOgsSDAzZ
MdBkqsYQ2GcaQ1d/PCxswhdLCY9KFMGz0CozpIF6YhS7F65CxM9ePjxu0IuelwZyN9ZWdfkbVLX3
zo8El8fWrzCVqFYiWtn0NXeWrZk0kdrSlg/k3u90MwvOOXgaE+ul3ke/8sR02E6CjDb9mk/GLEgp
isY5lNXJMsKijGLrvLxLM8Fp7ysMnLP88WGEhwFyPuoLgczJY5M79oFomVjKhW5frzlSB9H+hDRG
sy5oshymj88Zuf3/ee842Iv89Ut7Jjsfwbezslf2BJKFtJbsYs1L4HKKmbxWrL7bn0Zg2d1EcieB
MgWcSd5IwcqLVymQGCWm1FZfUO/niGJN09TYHiKVARe5KSZ0CfwkTeanMXNE5X4/61CHSk7HxrWZ
rniOKKHOcFOrn8y3iiMo37f+xG9b6upOBOLSDcNefjxTivpky56lGWLEl8uNvTLus3XpKVNLthGS
3rsPKMdOI2lp8k7EIYUtVFBaCkCt2/Ly+vHcwXvzH/TswnoI16gJy0TGfUBuL5e+X4MbtvJwmZ7f
qQIBuzh3oauvJfON9y+8lsjOWKXyEVCG/+Sto1ns2H2L8N76rCXUjNv3iTBfEZtVeEMeI/wWWh8S
WDreRgYciVFgK+4spOTy85Yi181bNHQ8nxmqswDuAnbT3iF4THEK9a9EnXiClt32ynnX4CGhh32U
hhPEs52Y+K1FLpqcZbUQPvZu5FGlIrVtGDues+iW+PmPpfQ/4GbJNS4Z4ICr4fIQpvyp1Tr1W/eR
VE32HCZiGMfJtGkqkG3vraSt6zOA2W3w+ZHaRBGmNVIYhDLiv9q8B8Wf3fyKKBQHFVJHhDgM0B3t
xMJtIxTJyDNSE+1odS0t4v0yiizvH16SCvBugaK0eO46hOwDJQ4vsYmVw/aVYhlM57YCLI6FMUVP
phg/Ekz0kqtnipwFUGG4DTS6sdXz0C94pwB/ndcUVeezO/alVQ5pgC4mZ7QaO4XUwMtxqXumex0z
Uagq7mKrQbR1hdEXGRgoW48zZontoLMA64SV7xcyazjkwvJJb7oooPZeSSilkOvvQZUZ/pFQnQi+
fyxBtwwiAcLx4NPg/7a8m/iqamcIiYXTspf3ilAjd0tOGMW1t+aoqRnHapP9nd+HxlLuraTEo5YW
6HSPo7XPUy+YUIpTtFEwK4OCuMnH1mx+gWqf8/bn1JzXOfZh3nwbRVZI9N0oH5X0codTiGdHOxv0
WbC2cn8dwjSVT4P1aRgC9pYn7CHdMKyzrpGxHucrfniTmqTVCGfosyScGzX8ab3JQEoY88r37Air
8S/pht9C5ps80Rc+QE3axgL9Upw4pSjd2iGWI/zsBFMXTG4qJVtcA5dDZYGhmMszRhx+EYJjJB8f
8nvLWkpnkjiNmaL+l0++MYS35FZ0BirCVHjjWL2xa/jrUF//qa8NwSHxWyZI7aR1rYgsO9PHCmc+
dhxpaoiQXykownO/LkGwEhCY2KpXaL9wMvV+UI6IvXSo0iwjppTV61yq/WMlMy8V/cULJG4leCz9
IOGrWx8SOJGMHAoZBh3nsWQrtJgapw27d55xfxN+cfFv50Jh+XrDfvOusS4UmaXmGrCZSc20nqLL
SbCVPwpy9HVQIIGIggWtEx/jl2BctDbmvZrrgWRliGRnQWuBaaI2GFIhtl5JBfQzXPmeeWxE7mtI
Fmz81SSyPl5qkiwj3sADTNLLUT1n3yZjN1SKmGCiPcI8YarcqFlUNfzsJmrg99U97fW6+i28eTLX
jRncgmOSedFyhAKAlbdwtqpOtnTc2dzCkJEDqhCDAQBGUqnp64KpXRY42ucwIaM9OLASTvQ+O2rV
GiDp8gVrsLCPkncQcXYGNEu9Hm2AcGd9TWzXPhamJqoglF6Q0NkUNm+FVUDi7WXa29IhFUsj8ULb
dwQLlW+R+Nq1eAF2pafHoQCYKGZYrTS7CpLmKdYhVkZtRo20BgUuKwoKHPnGtnFzE3T6/Be1iEaZ
VwzISWkwAaes+15twQvVra5PV+yAsWQpdsIATfv6kMD+Pl1HYmhoJm9vls7EFfXhVJWLoPS0Ppqx
ww2TNkDp4QZTvCPm8IH1DIJ8nPpbay4rQyl1QP9xee50T7N/dZADk5PHYS2B2CkFb23wh9uAhqsy
rsDjLVHdzC/U7wojQWFtrvK/Ve6ArZ0goMDGEv6MD+S822/KrQ1E5RDLgeUb94jB9opcn65vuzKD
vQNA7Jzj+rzDVb+I2TEZNQrmtHUSn3ViwTRmz+VT7c2J//ge3AVpO2E3t0F2aNWOFs7HeEb80Y02
1byNZcfZGAoqbLAyGJ2mKvcXLV5CsGhGaAgR77LvtyUqL0ic3kpcfZ52L7Gu37H1D2tiDxhGiomL
HLYydIZL41P3deE1jSiXS0rt6hNsufSXoIB/IHY72O+KbF5xhPJg3QzrsX6c8dj0U+71OCCBw668
huc5uxf386sCTiOV9YOEc40TstwrLNPszXyuVbQPJ3J2YrJ20Q8EEkUb0FXE04wDFua21H9UMDRM
NxoikRYohLG0wfpD4eMVGsTLvsQbqNBG3btx8ejzcrMh1O5HROnJqRCbkwPBtTzfk4oLUbm4KDZh
4QpULto5Ii1qZfKm6UsYkVo/NGnHhdMfugQnNKR8IvgNw1Ww0hhmrZGCueBkA0gHpQxEKpdemZEB
xYpuhddk9A1z1E5CUnejudlOgxt1PgHe/6fmOyRRyBHSH5KQH224A0bm+gweq814Q+YZKYTPGCkT
QUdmabCvqpWJLyFUMsOAtZcZ3m4nHH4iW2oDOg9D7rOX6anakDQsrZDoZeCSVDWHA05SGJMCQ9dO
+LCb7cBLl7GbhvHu6LXOg2n7zNP6/qvz1B8rCoNpb7vPWQRFH+MnY5ksjdRF4Lg5+98OMmv8R8c9
XzV/R5i2ficTezNGRlq3lNtFFrAudmHbpy2JQAEEYokGO1lgWKkKB2CrRM8J0ktZQVE0W3RVqscG
HLAO8e1w7Kn1KjX296n2yNiMkAa6pq360m7ZhNxEzIl38eHyD0Tqez6FU8auolAl9qzkG+ZCA1Tq
Mq4gVD8KiRETRm8WDEBHiWwuVzdaLfknBOPXYfYWa64EDJhe8JyR5RHqW8XjCaRbn4tBlooXDSYp
hN/tbeTpnNRd2arMlecUktOROvGdw7r+xTJZx/NcBjSwVAddwq34aCeiZcYFkoJfrjiJHs5O/4G1
SRV79NzfHAHAbzyGZLSh6uREWck2HaOoh8Aq47t1Vt+Gc0uiVuW0ZqqTUAZPX4wWj2hGbxC6eV0w
crnH8+haLt5Os8E8HiLuUCg2A7EGuszTaSUWM7inr+Sa3x1eYy3TOGulZSWmrAGQG/VqUOFjn+P/
YqYPvBiDpgcIkuLbWmgmUYEEhqWhq9YRxIGtU1JKjOevkc1vTTT8DUJW0Md1rEa+FOG4EeifaE3h
/tjRzDSQdzYUXgfW6bYR+QJHSpJ3Uk021SoB9KhAfBg99+GEpzh734YKB+KABtzZhQtgsQMDw+po
RMGimJrBlCNPpgiAD8G90G2XCUzTTxn7KlrUfcMweaaCEgNiNzyV7UdLLk5QPOWRYdLl0kfNhhJY
bjQCeZBXoiS5HoafW51f9o/hIgDgnyVj2whODTHVupNQFSL+5mqegmwNZ6c7lnxq/r7erx2qpSW3
0v7byh4oz9DGftnvnRmNYOtqJRaerB3/jlv7cvfRUArDhu1CZZ6JCDmGcjYHGljgp9ARqPtxlFBE
ZQJCfGCWa94LENmcA5b3Of3WhkUMfiBCBTkccBcYJvnDyU5n7R0eLcaGqqy9nFdkV84tM1d/I8Bx
fv3AcWkuKoFbB999gKuQTRI1kZ8WC+rggKqG/NA68oiNoZCdWSTDYbuh8gTYgDSmlQ7wfqzep0kR
Cmn6Zg9WuYqs96vK1mCqeVxMI7cL6M52PsvEoh8JUYH0GYfTJ1S5mO4UUdaY4qmHVfu54VbHXLa7
EJl/2hh8knqoHYmWx7FwU1L4M9zNfUMRueux9WIBjV05L75tFYE1DgxZS7PyXsdPLDMwBFZZi87/
3xqnknKadSu/UEFENUC9God+FEK73Iv9bTf1RPRe47zzXZXAUBcOCUERj6MvxZXe4PzDdH78PktY
wjTlkzhk4N2So8cq4gWT5W/Cx7V+3y6QVU3QP7hROCnt6qDPa+eV5vZWtbzA44Z/K3UDzcmlTA9Z
UkghwYQ7tQD6bxv1ZEVAio2888sRQhJzFB5bWDmQMm3qR9c8sRT4BWP6LJB5Y23IQzkpTFHaD3Dp
8/CXbZzQT7a5EO9zyWjEqEsgf7Xz8CpY/uIVYHJyRF06bTF4Ivoj96aZ4TQQHznACFOUn93XNSJj
tQgdkd4P3z9LkVD9btZoagtqBUOS25ifKytmt+6c/Hv0G0O/6UpwCAfYPMUETaMvuYgCwgd7UQhx
h+UdCd3CbZ/idGcHmhWpkKTBulfBCoO5VCHIAInvBGfME7LCR8TgWyi6zbSpSw6/KxgLluIAMyp1
oj0hcJJ4vpBNVT0pOmRMQ0YLQwSlEaGrcAhKCdzYgKHfbIE+NdmVRtRGOxnxucVkOf3DYRgCA97f
lfYYufAJNdQ8GnMVF2Vdat+AFqAtW682M4NTXe6xo6JOQwbFessCM+cZjqNfD8Tg0mvWR7QlwCiR
0H2XnTRVtt0TVU+86C53rCfGIcRa0bmrEOW2sD6iwzenPwTJVO7p/Ba1qYXK2WEisBRQ6a9IH6iJ
IIcJM3kCRkj2729HhUksRzn6nnS1aKvuHZdG6lIfAFuANyZlqDajPEjY+CHiff830MS0SdBJnO0I
gAMq39fKIwhTIEfsRmu3SyxXb62sEMttr9Le8ZzYqtiILc7iLpBsuuIgIh8QQSRUatwH15N5Btvn
tqifDwDlnwUPiHgum/xLCWWjBiaDdi3lchI5rfIIk3oo7QlBpJtWkgAKehRyC4dnQBvGkhpCwS7a
ycNR8BiFERSZNBpy4m6pEqG7vzhZscykSncghunzPGI2E9dBl4eXZc7FwdjMGs5gDcN7ArTlogjN
pwfAsBdgjUsokTOiI7I1AqsjhThDemWQznU0ZC9NslaTYwBkkQj8HA65WDzK7jS3ujRRzYhk3sbW
Hje+ju9+spzsdDmkxxAADvfd++yNmHZ621CqdFpS7s0QrJso46nW7ioMTpeKzkWx0JwkkbAiPuzk
ttCkHmAw3w2eeTdcnoT2+zSTiYt/t+9sm3VxvqeYbFug6vjEfIi9mruQZzfTfnr9qpwp5EGsKgx8
GtgoqbtyleKFMAYVMD8jxT/wra0eAWPDfm4Lxrtw9i9bYbyLGczvWQPXdmbWapoBDVRKOFYDSeNd
CXRhwfN4H4ZL1LbaTX0kLbo5fPstk+ApKv29SqVHhWaDYdH6doRENyvRCtKQHzgtYo4xpDG+sAGm
WaRNNYq7P6Wbe5M0eTdFSaZMwOPxGVIpJ1QsSxQ6KW0sPZLa2YWj0cfTAqH6UnN/MArak1X6eckl
BiF6yyHStL+q7nr/j7RJSr9Bb4mLn93u7SQG1EihUnD+lE62nw2M/3pETZXJcLNrw2OVAFxbyFWM
NKM6s0tlOSrIj+/M3KWPnLT6sB/y2MmjYHe4tHOBDHnEkBN0sDs36j0v2nkWijzoeJjdggSvBui+
faoYMrbsPARYsBzJS90pp8g/dDw8OEgCrheVNrC80PkaLGC+4UI1MmtW0EyocJAe4hMg9+l2p6tp
LanoP0hUBkqXgOP/aUAz0UhIp3j8bLC10BdaJ0SsUSLQt6bX2O2F5/vurniSP2kgiE6mwGMTkdUj
CKs2oDZ/vQlKEI8ZUkD6oEFE4JSEVCjLkm07/b/B6o3agg6vXV0yVk4w5khckYaRCTLHLyh1cxI/
1VH8j/tQme3QBQIn5H/0hFAmqbu0JUQJy070jKCNXmCP1PLRpH9J0JxoQgGq/ia7UIAUaiPfESRL
GxPElls3JjFTQsJ26Vk24feCY7VBK18D9QYqK9o9b5SnDzfVq3KXIGkfML4I9qXBMLNlqObEFVSP
rdUU0p8I+bNuJdmjLbSILCqM0EGa9Bz37+hUwrdDiU3wIf62xPqlxHtzGLJp2cbNtnykeAQtiqRU
NLwAjZ+WfD10/ABt2FBGl+O/+nq1aDtHaf9njaABxryqi3Kgn/cj6tZK6orTKya42jlU95kPNUiS
zL4zoMa26Es0k3aIHCeXP2QPWFuzfi7ZeLr7VGxK9l25CicTpRuWXpaghVPFCWc4s1779/U6uJE2
7heL+g5gEp/O5DJb2EanAR8SR00cRRFsGOanjW2/ohgSgtJMBmqNKo2CBUmsMalI+QWInxZsnLmz
nSOQjoIgRS6keC9vCWfGQ3WjPJhOBaJNjjSFGM/MNnQoozltjxoPDaFfgUtM/SV5fUsLJisqYM/P
eKfiRclWnBYXEDWhu81IUhJE/JbTLQrbcIS0m+2urUKz0YYxKZH0YfSg/vwUYqNtOcw16jKSyURt
lSNI6P65ex/XW27aLeVELZXxJwjg8VKTeSbJq3l72pisI7Us6z1hBjHzTKfUt1Sx7q6m8T1qjgby
SCzagQvvm0H17oWA/S1+L8imZdlc+tmHxW/krexHmQMOcfFl6f5K4z3HbT9QcUXHlu3M+Suvcgjs
mQTWhSyDQ1o8d9Cg6iy4C/7Tb8Yd5MFgFYG4xEjAe0VVScWNhR5X5dyrTDQ0kV8bpmHfYcJQ597X
O0FQjqp5dobWp28dt116lq+LaFt2WZCxTbaYcvzNRaT85Mgeu7gnRXMbscJ7EhUviTjIjL7n0DeZ
GZ7gKigKLowDOO6xVycHBcNQUok96OexG3giKYXKpeBX/jagOBWTZK7AOdVwdLFiop9j2wLQOTXB
zCaUTM9qKqqZJ6ODdLGLDlp4cLKQ7k8A9VPFoxWQhDdXnOJzJCQr9WkJuPqh7g9DlXBekx2I/8+c
/n+9hskCWLbOPaz1ixyG9jDqy+XeV7H4OURwdB10dMlTqW6e39wfJU8f6T8HIZOpgzsKQrK7OAp8
neYUgAagdVVS/81mmC5C5dkBGBLye6ueh8Z0mPtNy0DXlTQi8WvNzqIRTvn2EgEIv5gqry+Q0Wy0
CE6TLiRAcEhTNDic3d6uiIrIlD3YPIhR1ZcNrHCqNx1CUC+dwelMmRLcFqvMiKUAPQlF+XkltF0n
GHn9bjgVkBbzahOlfUMH4WS4M0hrlrq4LUGn4WHUrBoTD967pbf7tVU/2qrmSh/4etc+zPogrmvD
Hm5vpie1OQ+C2hNuHMHekBNb/jfvqz73Vn28PUj3vD0rr+nDZm41N/bVyIqsgAi1rBmyQuMVUxyt
mz4FowjureUJMdQMGbjMF4PXuXXOJ5JHFr2Qlyvt50nsy4Id+F2m8rBdG2NkC5e+zQNbTfkj8Emi
K42uPpAyJQv+T3GaYHc510zaeUT1Faa10OhDpTcpjSAq+367ZWsaxU9gezUWsIprKE67t1687avi
ystoHUQoUnGJQ3Sqip96z5iqJ1eNqZKeWUTLg/7I81RBCkXMulBrpttnsJRf6yDSeHnhPUSK+ii2
jNwlhoZuP/rxsMzWQ34/B16i+zc2x7arnBv/Wme9s3e00sRrB0XRIg/jYhGaDs3FADXV3BnEYQWy
ea9oMuMxiONQ0q4sU0tgMPmOZusUqBsCVuPgYs2Hs7lm5/uvougnwEVVQNjw2X4mcItvmFtzJ5YS
wqoD2JQunf+36GfDZxFkyZ/V/2fqQ34dX0Rh17IGNxocjgah3ShEj1YDnq6ktob1h3gbk7mCjraf
YACGli/f4e1OowzFYn5EgvIxfAaM/IVQwjUp/kkAYMdNde2nXBQMHVI5ZveaIwnzAkVmblAlnWHO
JLKeLnAelzx6SYSd8qXqe4sjT6BeD58JiDKi7YgwfHqQ6oRCRLh3GT+Rld2m3LjDQUAKyX6ScwlT
Fzgkpe4G1lW4eauypM4cNEkQUuaLTYopMz5iXI5Je9UFbnfub163PUWnGMyQKLqHj7d7d18VRzQL
ZY1gPMY1RYiMH5DMDP2Pp+OSqvzNwqwGqdGDOE2E7aL8caPmPy+2EBnn6b+0epP7MbVbU0jnIOi3
qwA4RLoUgo3G59bSXdPnrwG0ynoybBGPl/6wDusF8DXLT31gS/+6E0yDGqvmGku+nmas9PBH+cPZ
uGhiewI1Ob/E2enwU+maBN8OIS9vyKaw7K2EBHIN5y2BLQ+hBlE0Zb/hTAxvKLvCuSIkjlQNC2GS
dl23Pj1Gp4htnnSkSSDdKBs0jjoXhc7iESPlUVcyrMTHsBioCowgIUhgjxjoWdKI5+T5Gi9TqqC2
K1SujSG3eD/uRkwwbouCT/zGiM1GcHuAAAfwY/RqvlJ2SY/lvuPbp3+pbSG1TFnRII4hwCQ8+nV/
OdcIOqe7hQ1vAeqTCgDchHEcq0f16UUx6njYU/WTx0wf6CoRcBBxeu8ksiMEvmOugV7FhBPRPY4i
rIBXJTJ5d4QDZNRGKoIBA+2lY6ZciBPATqx9lwXMphaO8e3glQMRUKMW1oimMXVTVsrujEv4ljjg
k232Guwk7fK71zbYSPiO7PR1xbQcHBHAmqhKlkWMl/gPztx27ve9gY0PnC6KKsm5r6LTUR35v7Kg
zbl69MEB4B2ZZJEQZ30NpsiwcjqSUT2rr4tzdfYt7dBFsM9UmtdTtbsU1L18UYrcNufP23MIlnm8
shjc6x/k2cT59yVo45axR2Wx9VSHdlR/aYGC+wBGWdbN6ZDOsHrG9iC8+4WNBpHLQQmOs0WvjkOc
mEeKZoJgO3HASE/nN1pzj+KEPObQmgEoSkr5aSJQdxK7lPznVjfk1yDUbOuRrwz8f1rHrEl6X1cm
lDyBqJiAI+3wb4US1W1/0ZMXE3w64cS1zHYGQA5wjfpvr0ua8h+QEoXs5tnSP40Pmm8AZ80rEnsQ
z04aHPY16kXgLh05KOFpMSMwKRrciV2r8tJDzxOWE6nnqmW5FmAez2MBitD+2dzseembhgAaIt6w
lPSEKdCqkCv1YdbbZj5sGX8Dsx08QnY+vv9cJUFPE3en2x8h1XEB9wXNcj9EVA/6dZ/P/MkUkZuh
x7TW1+NrC+6UUgEPLQ0SQC3Q6Jf4TwrismrUc6Bvm2Nq4AMUv4HcZuNLPkzEKeWmhdzmd58p3uO/
bnoxXWX3mIK4wPw+QAZkcyenkwfp718NRv8QPEHDw2iNoPcQpaj1SCid2+Mg+5s7ZSKi7xyZm2OI
wRolVcNHbR8p2xSH9KLVm0p8ENMmggfoXIf/h8QYX0BdDoJqICpPX3GRplOlYKBTyExlouEtZpAw
366b7//rcBD3yi3Av8hvk+4tW8SKVHJnRqVO2uqkIluCO2A4K2m2vpwXyH0GigfJlb/fw3AQ0uJ9
R3Dm6mWe5WDuavWAxwGz4S6CN7H3M4hDI1OtjPjHTj7tcbeDZOTVbQEwrVjfcuS/bDCO9tU+mBsD
zPpQjzUrGPwegaqdihRvnZVZ/eOwr5+Na4qemqCqVeLLEmbW+p7DhIOCPWhsI7j45ffDRXNay239
9CKRivagNZm7tuRKKQFFFowXWMf0cwiZaEfIy9tH/8SpfmADgr+KH41Lsemt+6GQHKtS/xgC6vLH
44g33WOqNhkWTsMEdFV5/67Amgv6XtKl2YOSGSz9G/n7MlWuCp+3eACvZCTU7QXXgYk9Qxl+ihiQ
F+Q43ThpNt4kKp9c7NVoQrUorh+sKajE2Xkl2ulDl1nrv2O3J/6i3hP4QUcFBCuDmemryM3bqmK1
CIU10rsF8Ip6swjLCx6ba2yYyLQ44GizaKoRhXoZUSQFCAsMhaZdxl7uJn8kRxfWsKv+IN++FdCR
ZTKVO52NCU2BrSxwnupfHq8O4Neev2aqZIpzwFwwQnELLGYTBA55dggKN7f61lutf09NOo9w2LDd
a+TNAYK3GRdo0FY6V+ioHlRQsarcq9+Ez+y8Zq9skYoVxz4ezW7Q4kBRIqRC5/kQa8gbmIYzLvq5
35Yu2yAJ0MrypHacj2K+XjsN6uytPIPRuAy+GetDKMeeE4eeTdjwsGkYibx+R9s7m8gAR+Jui0NK
mvmNKosrUqo5h3BnmcbgoIVfDd6uGu82KT8L/Z44S/bmDZJ7qAN5y7N4sE2vtWGKZ3pHIUrvbnZc
hJ0FiQx5x2uuYVkOXbxZS7UmnLVxb0IrpywQJXbieRJf8OCDdtj0uDQtlVxPX6HqSJnEDpDkeU02
JxLqs4lxSvure8XdAi83tMhWmFoMoRnP3DdDjbJjt/LYBMAFLGas8nMmkh7BFEuIzqNfn4UsxUqY
iH77n49cEDrxqxBcnM5l2vg8jP+BCXYVF4kbtxvKZeJr0xCZVmoABfLTbjLQIYeprmB3rTSPvke+
gYGsWPB94enmXgohAOQFcBSz6ZetCj/WYsO7FXcV4AhsMar4tgq8ejhrbi0y6porYWzwSOgBqIQ7
DMPFhX+hv7C8jogwK4LOLJBVwDwXHlbCbiA7PLKTTvizremgxWc63XUu0hWJKDgRy69xBA4O4p43
JHGLsrhntkIvPZMnVa/bSDC0usVN9ycHN7jHdHBus+s6ARTnUKsnhUI2NSAEAQkY69idwhVlGi5x
BDYS9iCbFkk6zQG7qn+Q5PHG7uvd5UvzNUnMgO2mlGh2/nEwCjpxVxCNFpQYf0SJa6GHrNHxLcDH
h9B2jrwThbVywqZlYACxpQBLXym8zij3hEW4uzDiFTKHvDvb9iSdprXgD0oQGzia8fb4MfyFl07O
EwmnNS1+5Igd812suST1N6ELYMJZUTPfYnAoXMS/HcjmLCsSNuXAOBx3VcgrO5Z8jxQWdB/BelAg
QYDTM/FvhNtMD2JPG3nK6Gv5+9/X0z+PImtJzDiE+wS9u/UsUma4IyOrSq3VhuhhZU0KNuqKEZC8
AuNuiAeGHyVo7tnSGrq6z+YKsaO0yCpVWQdW/nvf80hjOdKiGcauJM4hKvGla1shdkDQvjDtg0Tw
bX/s8+eYyoRxbN4OpzTVRu2hFmeY+ax78T+Y18Sfueu77taxfow8m+cf/+BffGgRFyaAky+4hjBp
hFu2Cwhk6Hpu/nb3AcUrWRrbfJDePObwlLQhsUIapCPCxVKaQilqA6yavenk5thPlRE/TS8OPx4q
A21U5CggHdfcH6UNGSawXCu08xwsVTUT1+xQB6qj1kBXL5aAVk1mZCyI2DMWlRkBBKbQlPuZYalN
5zbHzGu9UdILosyGhrMsMugG1r1LZqRBa2L9yWj72scf1ZyYIvXmej5YaJYsX04g4VKJEMTDfmP2
V5h3Lk3lD0lDwLlKfqkii9E3W/F4dmTt/5UZ6eB3ClTOrlMfmJNS3pObd7cAP5Tzr+M+rZFmF4eC
K647ik7us6614zTZxRrK0bHeXR6eSet4BD/ZM+32EjjnoxDdzVWebNlRBXMLH7Tk8ubRVPw8fYb7
TkXOA/DsD7AWP/EP7wKiPkdAydd0MsxSBeaHFpoSc+/iNU76+SntYHEdmWkyPk1RuZsSNVAEeEwY
8dBTrGGUBUeJjCOV/ZkIav1ZXoRbawjYKRG2elz+yZE1+S0s02a+itXCI6Fnl8Iov9cwX9ZyBhXC
8McUrohUhQi5XaQVyO0R0iBC7DQroc/+npheQgw7w8429pDrYuQEr+tjeGj6GXw6BEHJsXwWSrsc
GuAyPFZ277UPLKCYn09+y9mnCaKWWSKsGxztpwD2XHlEnQrO1dQGeIMMlCbeluTRVoOJKbIxO1rW
evrrEMdCYMiEFMInBs7aZzm5WidG93tHTIgcwiDvhB6kwXIy+PmlL9/9WgAGJcHU7wWDJEEKDH4w
/nwhR0MdOHqLrHMaVd5gH52hmzMmf9VfUdEypcPUMWR7Jr/vCcBU+GD63dYKY0zUFpwtbZZ1pj2Y
N0v7tPYP8GmmvGsURc78joOtXY0EXFT14GBa5Du7UAhhQMqQRISi4u0lmVv3B9Yh4Imot4Y+gBQi
Wmp6AzyFouYRdkWwLSx7KmCHkaWepLlTQwogs4qRyqGvh2ZPHlWQ3DgzKrgcwTO0XLRb0kRtubfF
z+4Da2wThT4RVWks1mUiMpbwX7OzG20AnFMXR168Dcg0XhpL3GspvqqWST/IagmBPTgnekkIPFt9
urXqyOyMxlVrU1k7MB2inCd2qKd15Vi1dflLTbgTgJzOdr/RIiKQwzznNsBaBGCAGTlxMILSNhym
5CGw7NFKfv1oKsxaN7LG30J8DTCAjFwQPABR70NAckb6Q2KO/Zpmt73oejktpnH3td3YwaifGMR5
4sA6WT7Pvxmx6YObQ4XR2M0JohNtzG8r7QU17G103rZwgBrbpybXplOOd76gwUZmu1rkLKccnYYh
4tSC1KgQHQBf+vqYXXGdNlUGLCr0E1lw+bOZI0T/TxxNLO/ZMxUFbY3oS8bprl7nYuBfIEcXocDz
6P8mJE5ZpNiXX5lWpf1YS7UFRuRA8jk5Ryms3pLNo8dLl/APbDaibSm8bSgPhkKGeI3xcQn0B//4
1RhUYAzPVxjKKZMFg4gNIhqFM3JziNx8uxH07yDckzXnaDOWQ1Bdis0PD+9awna6VU9sSjizk3Fl
7hagVIzBCM1qUokbb1JyfIN1bHKj6WKRXobohZqoAI9UTXmtPmjqnyXsp+sdDeOSGryaodPLdObu
JgOpOUHfhw+28hysb5yA6B2OYCeWN7Hi9z1YZ5J2eYIj/abWGNjnFwd895CEY3+Qaz1+Zcjpe65w
buy+COczsSoq0ZFHE2znbb4n4jIUXCnn6a8AbfkqfWTVpDIXfn0rnIrNSGxctcwuZr54rA9Dgc8O
hbQSV65agVi1ER63Ljutuvktudf5AeXHvLFm4TAIuccXmmv2WDycHbMTHN3fbsnqRRW9ge+OQKME
LbD7DojEZSg1ghqLezwlg02vbNHRj9ZmuKYR2HxQTxHIZNZ4b3U+D4Bn2LvujrfgDMkf0bG2tq4B
F3M74WmtOj7UWze1S89LfJXWDAfD2NwZ3zk2Qv6gT+N7JfOlcoWG6+0Rfm6eBAws4f3vA5w3uEpq
akhpCNH98ZqP9M3mDokvzPd4EMrUNCmhxgz3L08GbFliafeSq33y8lwc87wrxZe3sjD8Vq9qf2/B
jqmE+PdPaEqT2wP3oJ1avngJO88+iYymn8opt5WEhI72EvR6NLV2HK9qLnrAjzXI9qRNWHPmb7D7
AA1NI1tP9jcC7AZx2PThPhqKU4LhxV12XObaYazOHw2OL/zTJ0qrm/vsI4L1pE9MUIn2laxRm6oP
Iu3h+xO51bIe+LWU79cF5HidFaqzHnW3KM0lptvbC9iA6+c5Xlua/yQVrxh5hJoILmximPTjQuzA
HZjbcrTsra4zx8HFU0e1eVD1/EJbLFtH0gHmYvzuS/9OXIBRBAKobsdA7EseiS9blVcYQvZp4Ifj
JwlLtIIJvmLnjnJgcwv/LYgfqAkTT0o0Ub1D3PLhlqI9A6xQsQiMZ9i0D+sPmArD5rnMBytdLB4q
mydXZkHqRp3kCV1aNq1Yffyz/zyoygrmcPTwSDZtI+3XtJhBRRX8LUvnsLT23p4RELApfN7JIIZU
75tt1SQm66E4W9XX4P3VYJF6NkztZIrk0eYGO8dngSxf/TnnjRmw/yGB4A4IdTvEZOWoVo7+SzsA
xqCuBexkgfYLkvAMYfd1zlLvv+/ny7SfHpG9d6qlh+cfUhefDfhQjlGSsjDzHlxfUM8/PlLT4WCw
UubMiouQwOF7wNiZBvKEk/qCNh+f6vOFfSfG2V2SpqMfCw2GFGBTu/eELSd+EYLCDvqnu1XxgiQJ
JN1FcIBjmGpT62AALxlSc7vlWy8ejODXQtH2M5NFmFSYQPPNNQVaThgmkQMeKn+1mrwIsfhWQ54k
GZgs9u/fWXY8MdfpLUxzY4+pj9uw0Z5dUV4xGAbK45R9VuewhEVWS8a3rbXAVQ7cSMeQIAixPi+y
HnE33Py829hOBNYYD0TGJyrt2bAt2eoaAXAozvAqEUXi1PpvuOzxGc2fGECrx/Frs2CAEJf17GPS
8Q9kVMW7Fbx9kXlK5a87TSDJhu35QY0dHH/nN/d5oF8QxSK2RMwpa1/U5bq89+vwA4qeYSwJyEpQ
Rh3lOTCzrHIqi62is1gnE+6NRxKa0k1WdmvBB+0AgpgJBrPUIFBIxAM7vwk07EjZ3zoE3+NgV9v6
4JCyfQueJEH4ZSIZYMO+D7Ci7HYO4ynfpOKqmdMRl9IAlCvdhpwe0yB88wl+r7bexiAD0sr+pBcc
kzfGzfEfhkUFT93bNlYrtl9KK8/CUzqR6JiNEgp1c4vr6lqTPfNCEiHY1YXehtrq/ek2t2mAPZaR
SH7IMdV4oBsTGBqlfolw9WVelg1298UfcxeOpxAxpbV2yNVhIxcwSF6FI+flAVfqc6c/p4dXWlSq
QX1HQuDHpvuGBwNiJc2xWZuy3HQLvMTZdOYpTaTTJMWSSQVtrD11jkrg8RVJ9dxuNDmK4zwMjhqX
EfbSKyrUPPBTwlo+p3a8SXHz4YEv7+8ZAuTOpO1QMrVacCTalrruvH7AEZgsl7euy1YXpvexJZtn
SiuG7qdFlWLpmktzgft5ycghi3RsRKoSqHCYod37SZeoIUaG4h2is6Tdz1rJnmdJ+xveCXjFHtmX
rdzCeVYn5yoFwzUCzD53Ch9p2h9TXd79XAwZu0B2T+f/mbeucf3XXy2J1hlV25Hj+1dymp8t8DrB
S2+W8ATAC/ECRY/Xhav5DiCDlSoS6qG633UflKJCNQEsnxlTQyq5ygt97hQ7PdFfv1UmFLF5uUyg
Y3I+TIsMIfXLDPfJuj1RMCz3TextZQ/OGeOfKmyS6u/rDaypl6lOhTVYirHTzxxU4Ro7Zyq2j1hr
yplerzy68eKThbEQUBZLqvae8a3ebCn72dPIthEoNZzRpHjplp813Q5Wgim9XQFzrf9cBQP9W0Df
6m5WfSIaCC1e15v+GyxO/ayfhzJVToIa3WrAIQrDMhCpRXfQP24yd71ulb98ktG2ZUUJeeLCSfP0
7VxyBn/CLmfJNJHi2SALXBpGSUgO8DRMgKhb6qsB3qgLIE8+pWXb9/HPtm7SERumrXFJlaNfEb9c
pOYEmFGzhqW6rVjsJp8C9olkJOTnXrXJFK5y2tax3xqxWB6smdy9iSd4lKIImUHMTxeDAfM95NqQ
uaF1rD2NT1L0iyXpArR3DdgAVwJmdo2W/kCZwUad8uM7cjZWEUHS5FcUViZDpvhVGLV0OPJU1Q3E
OvF96GtqCL/VBC1xbqSqOEzl+45+mLFF0Px2qFIkVp2arWSDC90DvZ4vM7nylSNO6R6nIXFD6Je5
yjhi19gf7gsTLMUMw1Byr6bBbuB88xxOyjwif6dHoqgpCKljUjo/+/PMOg52gBeBpCKnUBfgCzia
XlGSTyOAyKHbc1MkDgPS1qWmt0iacxRCHYL5G5OzglTYxt08ApdQHPtFs33j1ZaXGrxjl1SXeScl
G2fSmB+83/zbZIES0nl+2LK9mav7fw60Zwu6fAaoLsxTvMClbg2HXu2+ACLaPuJBv2P85LMoDnKU
oGVfArnLwAX9suA/wi3ROtM/h5zX35xbkqrR43FNRtvhyd4s0usUglH5CGLnJ8X+Qth9kxpwNVuH
EmQtJwJd5k/t4m0jh7544Umseeionyjz0voh5kDl1MScembp8mBbAYJ0gnogJchZU3jR5nAZnUCA
SyByp7TXh/3xZ4TMLQx+pFaghZzQYmh8TM9H2fPRdl2kKzMu2qSessrMetWMJV7dqdEGakcr1AR7
4wHOPRSpfQsP+wHLsjJc8JTMliOEiWaS8VOuiDEML+3DK+3w9VmWUtW9GXfm/GQbiXZGi2Y74Lkq
KVCHnhnALvvIHWPOpphk56rN4RwZzxJvl5G0S/qHBb1DTGNSF2g/F6SEQjaO/Ymy7dixtyWdQQCS
EwU4PYvJ8Pp3kd9Tl6RZGIIYPDwRWPMra8E3D9zRRQXj7D7MstHwoJf/OdgB+qlc1GAAG3XCWO2O
gApZZ8lGhxsjkTwe0yEGsgFuM5lg48A3fUR3YmWmP6mv9otdvWLv2JiS8QhgENq+an+72dgJEXNQ
zReja1rdQIw+pyXz+fz6DVML0+pGrJ5LpluhJkQFdeNG63q+tH2aT2JthLBbu/pZFqy74LOpXCT7
wJzoFyE4w6e+nmAfPZOSzRLwP58vgvdjz/e+mN01ItugQpiRbAOtnmdXzLjjKVwoVQZuUSjMcVQ2
aT8uQhkWCcMIuWDMgy3V0llw1zG6KZDL3MKHFAsEvRSYKwA1Hp3Boud7I0eHlZ01XWK1KpcVVuCm
P4/e++xCEZIrUNIxWNbAieujVMTNpSDRhIvMrzk8cFVnW559GfIZMVzFjymwpgrt3qAhsvyYGHMe
mk4iBUeGzzTU/JNbhys/ns8w7OKewJHn2WBLlPaPJM0EsUVsaJy0tMVPd8lG0m9+/cOKqBAZXImE
RJJSeaBDegPNYbMEniO2lO1p+B9baqAoybU5z0cKpYZcLYWGg8ygSqlFXXCo4KLONfXVutxbmnuH
ZDv4OoGRGnX0WbYnrmMpn6sD7fbjZ3Tg83IV7y+97QKgmuqu2zPegrwBGyTARJp5o7pDm4HBP177
QV72MtW90otJp9qMQCTG5oPaQEtn3atk3zJhSpMYIbBusa4KScOAoF1fV1RF3sTk7FQV2MR/zcNX
dKiVBqC0iHW50+iISpa6zn8dsGuQg0V47DauJKHTRuFQhM8aiMBFCb12e/MA8C7zVkfgaqyQak7m
0+89Sfi/jhEb8yEBMrk7rpfahnHJtDWxr+PRbRkl/NxNYqVViXd78XTJdremsBgausHFX/XCusq1
c1x6sGobb+bpNmdKgtHu5wiVTv8eRy9JowfkmZNA+N71M8j/XMSA5IFaxp+yINdrw4EzGvaqNs+B
O01dJWbLnKYk/T9dUZ59IU2PgwBhoBT87zYGCyWqnOESeLnJXuH02uA8CeKKs821x+h300zZU2gE
mYP8Gz8YXl3hu2ig/9MjAqNl2Fs3NGd/aeT3C/xgTq2j1gkIy5ukOANiVFiU1K7YQg3mqUM3nMQb
CTsjgfFgoiZZFsUGH/8MyJV0abqwVbXYCED6zJZiRbWeYns001Bt6+1983efQWM8vrmqTC05knXQ
AFjPVk6BSE56N9vLfskBsXMDf1iW4rLhZz34KkiwrScEmKbGHgVjUqDCb3bbBTe5VyEYU7c7S0U/
0/pB5nIuC4JJEyueGVHco3ENjOQYKhWE63ywrvkl5hG8epu4aZLjV4Bv32/a+tJFuO6wTpeMTGtp
swBdAq06FWqhbAIk5wDeyA190ZnS3Oh5NnNtCxUSzqS3wmACOb0Z21qt/00NMIdtE8mChpZbl3Ye
OApUKc/3R3ltydMiEVOUljzULVeTmhUa7c7Wp1DFXjOylQHNWwThfU0T/swj81nE+/hUdl6Ds07v
OhcRzihYTjw9F7DMXM8YjzM37Qjl4kmnZXUNsaAcOsyTdaMsFlkGcT1AW5tscEfuH45lrBlFPY/I
xC/kErO6f+b7A+hs0xcaNrbVOT7BTy+a2a4CIn8ws0BbjvhUU9m7vO/SaRnWC+NdLh3MK3ceoMJh
5J00x2mJ821Ur2KAJp4xuI341XMpq6qGfkodVEKaOJs5XQ8EQIQXDhWtkI4iGgSet3pGA8Kj/gSo
GDwsaHk6O2ccYtfwgYFjGWvUwo1XRb+ATXIgsaHPWf6OfanTQAC0Wx+fy+BrNW4DnqylVQ9xiKGR
kCKSGt4FXdDScO07oBWK0ysBihKGvzAQBqmZRJ1pRyyMv2hTvnMis9ae0qPm18yl06iup/XctJos
qfiXsSEfhrc+aC0DwluctBXc8jqEjVlLvZ4yZCL31/e+TDQ9x3ilivjM/NS2vidWqVS/SKfvIOnM
WZ+YcdpjlIQ2IMTkaCRvJPQL4D+C8d+lkTRn+KKrz+Vv2LX7OiFrAeVgtXHD991j6uR75edy9Eoq
2UwI2FPbGm8gpm+LsCRLsYTrgHt0yK7PYG/AbJBVZERfwnhDgU6PY0F//FLld0NcdIxzMdbc33OD
nyqdjfjfqcfmr+DR1HYSQWO8/RTDCOmaYtrfAtSdpAKJ4UoxelJn04p01AcPnrcmna1fsYstWeSO
B79P4VS/7ykd5It2MV3nCj/g2NHZOBYPQaynstip8lfy69vGtYGB0j0khaduD97Mt6VrOebiNXLp
9ZSShNW8SOfeXzTlJjaWQSWVU9SjV3dbRxiCCP98pRFQrSJEd2Y4CnqYn+pd1wkynoBYZuWxWGra
MLhHfQnlMb8hIIIyH3wD+LYHugxk6LNerQISj88rRW7ijm0mNn3JyLASjVoXMLtMfs7nvWkGkZTa
OgtWU7RA877QVEc0kpmTEPev48C98r9nZnJPv0zGac7ea3uXck7z2F9q0WSrh5I+HPBHK0LiH4+F
8JGP10xSjc0ev1nOAqxUKQqNTzQgwLx9VehlEMJ5kMplVLwkuvdTl/Jq2r+dXPYRX06HRFTcKlTA
9+NHk6LCPWYShzh9iz0Uk+pxJLrqnCpcwf7WaqMb1Ukr0BMEhetVBa2jDBrJogJx+4k04kLmtcih
vfHmdRXFyXJ5EazkEj8Z2VH6dbe/kPvOgzi0hKVXJ5eGmtoAjpHASsZzhwk7vHafH2ujGvG7674n
NQM5BgRA9IEjMsMp/AId16WGf2THGjcaA9fxNU5i6IoXLhtLhOI32+iWX2SuU+Ai+AuNitJS6zxy
ws5pgakE97lweH9tIq+av/qBuyqKP8RBwopE+5y8r23mixmx0UfwZllosOIU9gPvq6icxsot4nzE
cImgF9Cg8ApqdRHAWi/fj9f43PDf6j8IGfZruALbSNX/OQgQ+6voD6JziwMVjglWCWRJl3rwzW4j
MKEv63V0/rwv4oZ/DeJsHtKZ4gQiAWgm1awVYy8EgO3t8GPWOH3ngG6xcskslvSgMx/hQEvSAIU9
CAggXjdhUFQr3XB4qAx5pFoxtHnginxT6z126Al4iDOWR0Ei7JcfWJ2opcd9ZqOkCY80rkhzqOTc
KQieasKmT6SaQaEg5v6PecqAUQpYXecKjgShxmCk6DDp9uLdlTr/usjZwp7GRoHWFLE5U0KPjF55
D5ZzfhVw1Yb5zBFnmfvaQUWN+wagnIQJ5T6JShHRg4mzeRuwj+v9qJjhPNZCdL4YdQQLHc2Rad7Z
SbJV/4czGPtgb0m4CQnw53Mm4aDvFyRGA+Det6j2pEL58s3NrHbb/EAjo4SLblET71Hy1jXaJwYF
f5Y3A/G89OUHI4vbg+Qh2ButBYBlOijeLf81HmX0adXYH+wxAqTJ8fA6G/u9XJd8Zv/IBxLPul2Q
EkztOR096QFDYDysXppeGSgsLGC8vmVadWDPcnY5aHNQsIDbB0RHdiYj0l7kRjeNzkq2xg6Lq93p
B1sZaT4flJ54u4OeKKlWKTOUR8mEG3DbgjTbMo1/mEC6DvMEHIuXa4+arLI2+EDVVMR2Bgvycxxb
SLj6qV5gJYJnfWhWiT1IDw9xXzbAI7KzrI/JjbpffdP05VwQPVTEd9UemCV8KSfC8RCCLtyFVUQl
PgniTrRxUscXPdnBVofyvS8AsroG8XTp0Mur+SJgpaMk6RXn0vVUQXPWH2b0lQYp1ovTAODupbkp
zSkLMJ5+Cx8v88G6R03/hYO1j7zdl1Qj2VvZAa5vBnU36SaB1bhwDeBxYvGj665u0I19Arx72sFg
89NbyGUwnbZOj7iPlpx1zE3saVCRDgmdjvNZNtC0M8BGN2ez3nsLqTPe4TC+Q+cy5Eahld9cg+4X
0dyA/evcVNPMBDt1RnmkRo+byfcypTsFUOTpOm9uGDzjNo4yI5Wx7V3bpcQaiaGgaIrJvutG9Pp+
zYGwRSAfVbDM2+Ow39SbgS5LLuSftX470u0w5WsQrgzdoliUSui5VxDbkjN4mTZwu413zQ0ZyE20
8K/7Aiwnf2T7du8aVchvk5o7Kj24S7yWVXoJxzg6mYpIs7ijy9Veg0PR1PNHHOOqvvf+VkAoEy3v
qYwPiJP9SPTatVpEvksj4QZhBq6y7I2wyZsDf6nsXKQdquLntb6Hqz8alSJ/FM1P+9cTH9uZJbm1
TK1wqoA8cp8o7neVMPS+g2XEhaExW4AhLs3bfeFn3OL3qhpNWgdYpUQ7LXtDaXg4GGS5KZVNhavE
EmPdHtwJzBSLGMyVO4FLqrknMwbHIJ8yeDERfFKcNQPm8RVPG5VU9i4IxFzE56l8mE5fS9mJJ64l
j+1njn7IwYr6d33juBkg9FZMJoL6/GZ3bsxADIuyPRwDwEu6XrLyYdqjm9l60zc3snm+cr+j4nTS
Nx63X0auTclIkFEg+onQiNjKXVHdU4cOjjn69UzPmvLoOVcf/IahgkWbK6x7gkyQWLUnO8qysVnj
I+9mTK8+pvp0ed8GhjoLAQ+B6bYJDtA5xhuhkUrcVibPG/UwAOUz1Gl5K9EVJQT8B2kn3t4nhdiW
lGuOGFJqUujrSeZ9fKeF9nEHIeTm6Rc3kHWxqOytgQZbtXWSbHw5fvGAJEdPXu0vSOHE+XbBby2k
I+aeLKld/Tj5F5oLstmCnP7ARwuHoUE764I80SXxlDc0qQ4bYUp/DX2mKCJw9E7Nb0AsaHa14XOV
rNyrWzKeAm0XZT5UEkxZNhgHgoM24e+nkhSZyRtOs8Sldw1B4+rfzX60JrbnRjwtyDzFGM/FILPp
vU+oA+7cvm6AkdDB7vPDk66GZK63oD3TlcfL+seUAz0l/XXA6v8q/55KBu224AJflz8Y/JROL+sn
T7bVpgX6qJDHLc9y7McnGHkDokjMSG/CaPlQKWAKo97CWYb0EipTM1uyDlL6f3v5URCYz/Ffh0ly
hqiIoco2R0vocjj+dpf38hw2ASMAeu6m5y2ldGDRsLz6r72WKG2rlFkUcz0QGFbpVm9d5jykzFaq
tmyCnD/7LY9m8zi+2O5X/dcpKwjzbsa0ZhLbMPBfY+rmsd0qeuIkdpuzuw5wrgiTBGmnUrKUG0vs
ZWJWNw8tfiwbO+tKrOCASs4jgA/OqgjMBqeMBg3eNRl+IocoFf83vIhCClp/dcNAU/sz3ixMmF6i
GRCD/NJzcLzvW7Raclt1eLoCHtRSGFlg1wOK3xWHN/v+sMMwfV3QB4ih5scy3axqTMLFlNvGEj2n
nnI9r2gKauzeXXVJPHYGpCiSXfQCNRjct9QGuQbYhSTKA8ljoDfvEt6oFG3JtalPEEz+HybBfNCJ
mnBG5XtBhuYz2PkGDDZ66kWkf6K+8c5lLCY+uy5Lkc2kOX5/Hq2dKNOCMUGHSGQjIKOjyf+XBNHd
NVYq/sqt5wc/fgEvvcPMqMMGWBlU/r3RcknGcHDiry389qcFcDMdXZB3ZkGZVhNdlajmDRWa11Nx
t//5xNZtCsK1XdWXFJXQpVnisoYniKSdWhrxNvRvh8xXNCocivQhotIFIBuygeutmh0cJZXFXf7o
M74F4sxW45g21EA875zu2s16K9CCESY+3hzcAhVNtnNVi5BgmQN+9I/aW0LAPudek4gqED39Qgj2
F/D15SSx8eYa/Oc+uMe+YpzZFj4qAjMNT3RynSIo0yD/vAOa+U0MMZoU+t+OhOFUIInm+Z8pQSF0
IFZMmzFjaa6VMw7KWDoxDCWjvljDnXQGBWhr9/o54nrBI3z6tjaXZHRqV8fH0hycnaFYbzEAd+Wf
US1ntFSNK/GcFU7GcZ1KCueDd2dQzVRNL6fjLIklAKmD1hT6dKOGW7qA54OUvjuXVa12qKIT2goe
nqImn+50mAWsUxg7OHsWYQP82Vk4e/QjJhUpFVSlmyJ3YQx5g+L2XzBOJ11Qi5B8JzEgqK75wvCL
LNNhOIn4Sr3d+MYHjg8/hxw0C9h8kvQQzGu4DtcY16DT+wIA/QY4e6kyRf0mpgTMwbe/gdWL7SL0
2IluQX+EQ6qjebP2amfaHB2PqDlfHNN6U88yVVum8UBeKDqDC4Vf6IU8VB3MZDAhXP79xaNf2jEc
lykGc4f+kT6NXw/fhZa7cm6Pq+LTc7/41oUHpZ1IX95ZnVthZZZ09fefW7unlsJm8XSeibXnva3z
nCrszYgjJFx1chMFW/BDcIc5KR42RkutH7K8iQPLpvDh+NIsmeIwe51+Mq0Rg6TmQyV2qc2zwP4A
sSbxuWRJD/QGLzYVH/Gn5kVb5j/89mcR2CiUva5vOJOpFGtbefuaM4OS9kzWxSfRFQZjrqyXE9WE
/fZ0zcXGlvUTVmqjJ2oEMh4mGPVxuAmlAD5lCCOSl4HAFbV8MmF06d6zoVqsP4iCsjFDpe9jHoKE
z4c5leGhyWczYZhgivBgmtmQfAbXSwRj3DsCS9Q0tvjQ4hl19EIaeqDSUk4r6mOwY9taUPdpOVKi
KXP9QWUKSF3pgcTbHOCatbRvnfVlptP09RGy2T3yIByhuSAWy7rF2BXtk1vhn+ZHdY0ymESIZxDj
EaLlwpD51lqdlf3WfmIndBU6z+QpC0KsWahH1HObAhtLZKlbdAGGYXD+IYM/g9/k7x3unLr5eOhw
vC9kWMRgo9CQcd59Gh4z+xtT9WXJJSxx2auKMMtKYHjITEHj0UwwiBL2INaWKglITBQx4hfUBiHg
E19br/mGalHcjFDrkCj+0RDmyq46dATG6ZMOFRI9F2iXjpIfgFC9cu04CItM2g6Biybkn8uulRFw
3NW3dB0F/xOV90m24X2eIv0fWqC5ouLPkrTwW7ym+baMTig8kxvqUC3Ny2nY2GA9GGaBrgI/KZfH
5ssegxYWwE3gX2u+YmKFqI03e/JFbfnKPQ0HBWwAnjjK6zbArTF/iiSyDvOoTvLn2KUjGMdZJABN
ICHncGlXk3Kmu4bpar07PCKFJsI2jn9sa9x5TS21Gs5TMjcVFnZvZJdqa+Jk/tuGO9NwOUlQlsIC
FRu6jNxK6VFdn4l9KYbcS8atkv3o/cUyGHOx6oMtUkMYJBax9h1ktjj3jliTsiMuc3rSPzjpB9L5
6uXJmVMEcoMCC3Glg6lyf7eHwy8Ohbkc6SzeINArZIzN/UZsEQFg9aB0g8vDJtuMsKLaCv+ZFaGW
D37zy52196KdTE1/txFqGIZNBHXzpLdEwLdYUw1j7PRG/AbqMtu4YfqYrlPZbe40SnQZPFPfoC8G
AshacmTArCwLpS6LIG4HPgvxtIjCM4shcBexTAs6CUU2ArNbudr3p07wQpsIZFs7KZWqqhoaAHXL
SssYUrXcOXUfUBno1PxM0ZwjGVQ+h66cu7fTEipoGun8hMvGsW7v/mmWr07FodKdECjNNrMLWZxj
VbNiYTxj6PH1CKYmd/l4JZtmUqmwAV05uB077ZXBcNPNCoEgmezz+Fdrfx9cL9FSjNJqjs4k2OtE
iIgjPvZSn3epNGWR74BO7PqhiorC1Z4LhuDgeeoPdj9gfreMD7A0R/Ok9Y0KxCPNg+BV7gJEK7Ky
TJg3pK2HfPL5Gemn1WkLJb5CrgErpBt+/JypP0WT7MVo2VT9BkOSYyAYMXonYtj8P7g4zBaBEMiy
ANIA9vJ+Ir/6Y6EMDgxp3tqYdAjERlUk1dXWyt997dcsdBILPr1Jy7+/bb6GANeOn7OfD8sBILgN
CeEFP575XXX5Siegec9b2JS67EeJmuFM27vQqQw/hbjL6+sis1Qw3A4HyHSmp+8fnaegoJ4qRr95
RzxbqfNE1FieyBoXyQ5DEF9Eo5EYmrecj5EqykJdYKI8481UCXnrkW+VqZylY4J/QsoG8Ra2dqHf
/Hb4RgQJRdRkIyklkDdacgf9mu1ARji2ugkdov3ymFmfDSuqW9LByPSmk0WiIctzXSEMLhpBpW6Q
XqbLgcS2nLuCUH05Nn5s/NgcDRhwsb8v+fUA4YyevLlfLaSdhe5zlclfyBdoaIzrGYjka5sWfugh
0Pl/tTOGWu6uGCDP7fLVg6640SQF2LVkjupD0bRnNOG0UREaCCX6X2qJnwG6PLZ+RQtW/paQiVK+
xuSyGFZic4C5QA7auucoZ3CM1nxI4Kn8OMsATJ/52NrqZkB/tCrx4RlaTf+1KFxYqjMw9rizFkcF
ZfMs9qjZQ+Zn3CBfzigZFY7EoF60qtCOtHJ987XSQHf21yErEg0X1DTdr9nfoFrdh4Il5jQxjE5h
+DC0Z+gj6oEzVKy5M7h9Aq0aEvThTrsdhCsAFQT1FURxf3X8UryLrv46eUlrgxsf9a+TbAw4O6nn
JyRfBFMI8xeLOOLnUfQDrS8WJnxVbiaeb6yXIqzod53AgtNv1bharS8VrfwsKUkpiBfosKPeJ1/4
8WWQdFxA0vjU9b8eqiZg5za22+FrhLPBQfiWZhqsyeSrvXDhnqJSvQy2lFIv0BCyZZ1iyH3PFoRS
76lWOSPmUM3SEUPFLKG+Kvl3BcPEkVkqr38KzRBBJeHSi7lpvIGna5uirLyEZ8AQ5JmQzKqQSPLT
A1L/bMZuminqTyK079rTivgAcJ/P75f5BoCpZpleaNNJPFB5OOQBPp6ZWLkErJfid6a+o/0wsBB0
xOPlN1qq7kgT1kBgOpZCEqynxX6qvuGdmdUBx8EdScEls66w40aEZS8vI9bZ2aaV5hSlKvKNpxgN
0aS6PultxePnULoWYriQH5cuoseo8aDj9VyDELhrpy21AGu+Z13mxBJd7A1pOy4ReAfOiubsTlOV
DPG73voyEUQsX5SKJr9hnV3uLrherV9pZzFcbH+fpMsx/cR41fuRLmuuUgUn0dfrBti5/4WZofJG
CYSQUt8yQxFsshpeEISEcd/4s+8phL0arCFEzXI04AsuWB2CsJwKj3kxpNWGbMTr/O1fRCRJsT6X
bIsYB/qe4D6i/USPYbWp3JiD3b1oImoskTR+V3yMKC5VipdorAu/3KtVn4bGdozqeUj08mrwR7mF
G2dsXYkuTKHTTLbJVVFw+H+7lVcu7imreyvQCPs6pJFS6oJK9NnAOhK/77HFRLy6aMnDgck8dJ3N
rWMvMeW9ZQ52mHNvdeaG7WVON7xJ6hGweoK7Vh37rn+kvZo9wnzO6Rqi8hoUTImDWwEkPKJg8D3h
FcJFTJbwI0ppeKqf1QfcOHS7oLe7p6gBdMSfWzRjBpxR7mAfUBH6M4tOztgE4ixKWWyNnfJHQMx2
MBBzVs/A5iH9ryowTGt57/twWE3dL4QeahPt6VujyChqpr7RH8eiDEXOzbMHa64mHiqEYHpLoAzx
fJo89GS1PwwvkQ/8IPptK4nR4ZKY69CMDJHk7Jbf39gpR2B2Rp+rbvgLXjz8E+K7udeKx4BKbbkO
KVyHb2UU9BsGlcuKgfxwIxaDysYBScMd8MpGcdf3jVSmVaFKnwk9FlYU0uVQeWYb7jA8gYed3TkU
WMQJssZuBUGNDZAoU12f/pQDFkJLKMMC9XUYexwx5/7hfC0WdcAtivsf/CAVV5TKRWHiZfBPuoR0
79vSvmXuGvw+/RsZz/o9FoEiJXe4CuRAWY/gDL8tB8AoSqWGqFJmgxnIp0ly35RFNdKpjEup5rIr
ZwK3CC7s0KRmyg2aB9V2y4dCsOdMtgr3tZlk1f9vvYmlW8FHmGkAjbWNDPFphldNOVN6cIoxsDtx
Fy4DY43BWvTLAJ/BH8/jYCJIEDwr7BDEZg2b34qW1uiXmdQOxhB294IfZXtyd/gKuehP3PvrUIRo
XQGf8sElEtepC3VAHWwohgJBXDlcoO3M1vxVBB4uSYvyzyreJIeIOTs6Yx9wyhzOUolow5eXZDQD
v4BPTlWeyqSWCsO38J9VLGON8ht89MVQwbD+aF5Cw3Nl8aGwZfaRl1+2kTJInQtoE5Pc3IpB0b3Z
4+w0icezTQMDwnh/aVzE+ZlJkyOaaCIJkXKr+9cIptxw/wgez4OEZjTN1LAmbpiQp/xif/MdmfCl
rJmFP+O64IMJp+KX7h1C5vQDraLn38WIWquaLtSvSeXbN2LxHpXxdoDuxjYU7Y2dGdXborLyxJFz
SlkfhS6GEc21RDaDG/rxu0IDUSAwP5GkIEQZgNVAkxNvQ7GQSikxwUGLfKRqbh5hq79fJzP8Yfda
ODbkM2Y9qfnCwptBgwE22b9kSixMbpHbgkqPpW4AU2unF0AdgU6Ukbae+McbI0jrAdkcIzELA9jR
j0DE1SZfhGhTTsZHafTbBQlRcRiUXXlEjKJDT19t6ggv41A5KSsJimn4g61XsSwyLLYWFNDXtGyg
29gG/rbkOgpSA+P/93DR+nKh04zcNSfDiIrGbCC5OXwpwp4Y2v+6DxeDeQfAflBIAtwygxkuF+DM
41YzN+6zBsyJBtnJXBk2V2XbVsD913kPMtcSVBnwRyOeL84EimA5+XPACQ0/28a46z/gBluuO8HU
nIK5Rjt7CKXhuyMT4DlLyJSYkrAfsgW5TCxrQwV0nBW+SC2dOTqeIj/+TYxcL2cZ5oJIUNnXYWBA
ms3mu1w5vCbmn7ed5QLfhobZHw5/r0bWvMfFUDiZNIrrlzwlMFiqYbMyx87coQP6yaCerbvzo8HI
9NqbX3m5sJ7DhKDqaob7M50fk2y7GGIUurg4ribdI/yy9eY+9NoEWbwsMtzNVONJmnmHZteIcMG/
WZULZJk+XCxACnyWHOR3xsPkcuDOJ/bj7wI+vM6lzyZuHrMC0w73HulN8V9ELRTxhdNbtQS6WKmi
tdNDknLeCW8HZ8wG2KnPOrclbf24i+dKShKRRTjPrRkMfziHzzXFmsMo06abkyM0Yh93vBAaB295
jjVbvWFr7SlcKZFrL36j+xXkGS1yvS0gGYoCxy3CuZLvFDM8aIw7gKAdKTcDMAedEh4pDtYZJHcp
CD+Ld/WRn5n6rxItnUX0a0E3NV9e6VwKBTJPZyI4B34JHfhQaZS5jKERZ4jwz3A6VgkBSCol8Q6d
Wkyg+bZj3+M4Bxv1ECLtcJaori1ug6NSHPgY+OIWAxqI/lOwsS2QswnV3C7H8S59Uby5aVMUCTpK
AD9reYKF62Srn6bxKr7wwdqwJF5BEFgsDsEVZIYtQoi0WiOZSChsldHavd59rTyrouqcP+qspxFF
nffK847O52U+EERzYMcFmPWaOTJM6XMjM5N59apyBQpuOBCvmxizUVgBsdLruTmvExxEIhFXebRS
PXQ5FL7Xo1r6GCzL9hTP8JT8xxl/pN78gq1KFuqxChcM01Fwbm2nqOXD+awi+rmF6oOtXP/MvDom
Xz8cZuD9rUONM5n7V24L/wZbwYM6gVoqUS04x339zOM2g+RF3FrxtSU3Dm3eyTCp479y1hGzZJVk
S8PhOrTeDUkXd3f7TIOn/ZEEnCxozrxmll465Olk95xya9JzKPEn5z+wxKcFSykgJhEwrFthUh/I
/DYM7rJ0/XbRCxVprDVUH8Xy6wYctTrAS9fHtmWThBM4/q8a0Nh5waGnMJ1mIHXPe//bcj72mMoo
IDiQ2MI9MeHKDInsOo1M6e1CalLtiot4gP4hTtPBTGilRe5emGP5pYL+rQKjTXNILfkM+5T8nW41
Tj784AWS9Otjn/D5m74JLDOqWcG/z+FNHv1IlFXicQFsGZleBVijRxOPoid6JwDlp3HUL3gyeqZy
oUxh+gMzVRxBcSMAesqmz9u4zAs3CHBODoIKbAIacLO9GhAM7V+Eneo2W+9Md9MQSzgy8gKzW8M3
1dpKYUfOuYhtmPvNU8V3Xf79KcWGdsPhtu5jOsPG2AwpEcnBuXmE41csAxBbx8Bjf4xBN5gKqW3o
MA+nyf5k5hnjlbSocTMlK7VO9cdpODegMILYu6Yr9DUfvG2MPuxZmjU/G2XK6abO55ZKtMzzdAVz
qvpXWpIwwpURG/Rr80+D3aRh7JVhOcsEQoIWYZZJQm/0fnXnS8M1dXnGvkYov2ACrhsiDcPCNTEH
v1lRs2UIsicy+/1Ppa/BYSmcC3Q3MdUt5rmVfttIE4Wpckc5WmawHCO3QQy9JjMiqehN1CqM2nOH
8KAr+xkMw/Yo5fbLbQbtgICmUupjEFt5/DyFaQkbjY88hRSlPDXqpagSruxPIJNY9Qx9jy8j9nHm
86Ix1g2fETsErmzekulLlj32HtTns1UV2UNQh515zrJD9J+LaiFwbzIZ/ZOPdMVDywsbJpCguEE0
qdKczGbV2LFjQQFbvpFnt6C1FCBRpAViM1HEk/q461v11+L4BD2TZsgl/g5SL5Y3kjxEumS4f9WI
sgKmhUgh5QjNj5RlJnRaDewM9a4rM5Ng54HgFdV9d7F6ZUvuHfNxj2S/DPRLbZrYJ5Sq7Zk9pzgd
bgJfvitxY2wN6FfTBPLmcEOHAUzj6V6IZbSlSpNkqYBQXCWAr4Mj8S9duBcWDvggCn9dm9TzJfC/
eNMqSWjulB1rNW7c6rT+bHN+t8E5OYiLH5JC/0kKNLR88YGtTU5y5dajNPp2p5m6LKoyjU82nw5n
pzUp5jq6uuoMB6ThKTd+ovTWeO2gJ2DWN2AZfJaU6o8MD2gmPPEnb4NHM5eUN1b2IMb8D5D06GyP
wtOJZUjw+6wxLY8c7/1IjNYrO2n+uCT87rYTfViHL9QQO5RmPZ/PrW80JEK0rm9B/g7KeosBehk8
jHvHBbBkwc+pckrScGAU0KTLYDgDWL8jG/L2IcEeW/9YN+MCUJz0dtc06ZKLn4HCK0hiA8RAiNVB
LuwsGNRasFthf5/CEJ1zJpq/Y9tBQ2Yn/m3JY8fpW/dIcV9oYIDxENoCrbVxuNuNQkQYcL3sV1uV
BBzyCWyN4u0oWAGWB6RI5dMHNo3JIEnY03G5YCuCfsJRinEuVktZb6+Ss2gd2gW9rmRzPrESCHZL
Doo5VmXa/rlxNNgUMPRpSyplr0nHPAIBgGUP4vLJD8/RrSAVvE+NDRNTXHGTTDPVySqNPabTExuK
Qu75Vh1eu12NPH1D93ZMkTzsbXfZy5gXbv2m7kucZEd06rue1X1ZpaQQ5OJd38rCXoa9Owuggr6n
KdxEtnN+lmuCUWwbn4HcafeWwYkBw3PoOUsDLWn3HJmUFv7WTSIl13jni6PAl5PuESDMRAoGNjPx
NfxBindbZMmEG6PV+lZu+FRatzqv8ix/uey6qOFhIPs99YjJ3CMKvdVZJ75Y7yNQfoAJgYZHNJmH
RhXc1aLgSyozUNYZZPlOzdEGoTKUORx0UguwcvTqRvaKgjSwmwA3a4tMS0wZA7fmPs+bPX9URZQZ
tG3lIvvWds6jmpuh8mGQ7bkZLx2V9H6aPbvGTXCZruEkX+vUKQish8+SDgGFhRQ5AqqCQo9kcefR
uQG+HAC5NEoIIlu7nUXNjOH70rM6WKkPz1wlbiJLcIl+PJpFQNIDvHCm5AmPzA+EwWwLFM4NjuDS
GVx5DHc+IOuRflSQ2LJqrWPDFGx+2/AgvFc2KOZpuDkvS5YW1Ruk8sJ1aNRD4bvdbehCGFQyXSpi
YNIeV6fNvUe3uv0k/c0QddLDPTzHHqW/iI4bgHfB8zJ3T7APupgYu27SHrJmgv0s8AGu/xuZv1/k
6Yo6m7yZmBZYcTgR+kjOWPHMEO8/lEWUChtzg7l0n6gLbSWrAkh+wDdJi/CBrjV1uB5R4loaW/P8
gQYjeScvurXIy9V/mPfRGua04pwbgyvcx+1AwXUZiadrgnkm91oWcrT08p16vAukJvXOSeEHXB7w
MAYLOVNbRl47uybR4hSVvWJI/GW7T/PTU5hO8oobNR2ReRQPIq1PqgC8WzrmgeMCtEJsftZufd/M
oVtwkDRjzmRexuLh5MZdAPZYlrNRf0c9afX/DM5SR1Dt1bvR7yXy5b218zOeLmR2afXq1+oHLUyO
Cp8Fn+oAJOiCHu9eUhc2FY7e3RHL7WzRNlkBFriGcg12FgumkaOa/99rx1nF1vOzYbkENYY5vrnG
89/ft4QyL/Uj2Qjfq70tYTwBHNun/iRJxFqOY6luLLVP6k3KfIwnY/MfvQVFlJgqWuvHr1OANhsk
JVIh94HAIoVFQa0PN6bRJTUxh9Q1DqbzosEVOPh3XDJsSU0BNmSE9XBlVHRPQOi/J2L+OdpzgOY4
Q1zJhEStMEWl65Rn5epTPrxwpjud0FXG2y7q4wRXQqYJUEkslIldvUIdikfsdCHtXXNGlc4d1qyo
GPl7AZoTuFaoMvhkOR40D42cjRshKCKyWLaIHUBtvEXWUmp7Jtj5bR2unzxR9tEUIe2LaI6v880O
eKgN7nvbL4spfGQov9UBDXu/uGwT5li3BxGyw459vkN8ZnrNBELVTp6X5RWUTMkklzTj6U73ZhYO
1juJ0RKdujjhHSc4O8C9CQCB6EpX57kvGqg2LmFdD+BPoCusiEq0h+bvfX7enJuLe3BDmj+1pC/P
70qoJQKtA/XUI4KLE0brjeXa9BApAJl84lc+uFieqZ2r+F/Zo/MNaZkfqd4a/8liTFIPlmyWyGL9
P26nfiadhpmY8Wwkz7oucQytI3nO1/MY3vf1ZiWZEsJRF/J4QfTjnkN1I6iXkYHV+wAB/ARiByA3
Q8A8vg8v7OcwhjqTpeDuIhOhfSNhXjLORcy50Ib81EY9mcIDUKLvnz//EsQxEuUwTmBEyV674j24
NBqdFbcTMOHqU8U2PDgvOwaucdh/WzvJc9kblK1uKbRuwwZM+bJLazSwpw3HFA4J8MX6ATKo2mT0
xnX0jCFu5DEcWsZEC5hhIykJvU77eTWbFVAk041/Zs09tyIV60uBoUk5IZIKo3vXpKStF6nerYJh
Et8W52xLEomicgW3Xipmg1VkziNJ6n3UB4xPdmNgMO0O0PF5WCZ4bQzWd7qNY8OHp2PnG8mvciBD
0WCnPrSP5hnEZRcQR84P1BnBa16dSug77PHf9SBR0iM7rS/a4nGTP3QUQTsyJMp5xTyrs4Jk/AmC
AMoIP43+/qNawXtvkpa7/2DQ43Y3NmSu0BW66mg7KD28+6dmBifh2AU416cFZBPjWw20cAhgxf4c
YV3hfKJPUzgpH+dw02sVp3lwoLG+GeDLwLT3zj4GKMB3r8/OFf7R+QvR96lB5wdTCy5UnNXZx49w
d8k1a1PfCi1T5AlicUf1spEdcjrgp5/6/pip8IodoeLkK6QV2YJo8SEZf8B43uQk3fpI7J674neU
Fa5qV8HS/HH8FLNFoL3dpXBtrMBElPci21nHy9Ccrw8EkK4NYZ7LV2wNo+1YvvuOd7KPJEHn+iWA
IEnzkD3VQl1VkoYA83IbjFnYSiFYYKPXSKiU7tfMfGjRj9R3QyeAx9vsxl6+YTcDS6XF0UyosJ1C
qcAQlhVY3nr3Vy4ADWzPdsh8RBJErIXc5h2IIP7nPx5WBxVxQ2mihVt19eE868W1dyjKgbehd5jt
pnUJs/4TPUfUJq7pA7d5cvC8vK6Qcj68uBMacW1KGT4WObQjVLoc9JpaBdAofLT8aHk/hAlNcOd9
K0UZEOQZSeSyHcNnM3g+rHqIYZvKOWyjM8IEVu7Pw6GjF4Gl2SH9jlU7pNjU1Kt5Vr+WDenTfm5T
shklDT9vkB2i0ooXGfX7BkuQ2GKXF6xhD3eLGjpgT/+Ok8TyOj45M3mRg7RJHKlK9ZpT1MKdWXc4
kjrnpvPUmZms1DIpPjLt0UIrGLp/sEe6/qzvYxlHtDB/WXMD4JO4zgA+jbDBOP41tdaTImnSdLB3
PYkIT2hIK1//E/L9WmGCksdchEO/dHOdJWPoex1reljJuFqU3iDKw+zmd+RH4NGCxeT45UGR00CH
Ur8mY67ZDR7J5jnuZIrdXw9UM3f9I+MNrsTwQp7RDLFsr0x9Ll7c+R9BO3+ykMSAik+YWF2pOUxM
XnSo7eaRFFbRi43qP4/sP0QI9oKNEMoO/O/pNoV+lT0RjKGcpEW2scS46Un/MNpoTp9gfbMRQi36
tXpkl8l7cyCyn4P38/WOVr5aEVijqkWDgPfLAciU/7kRGiMHU05HUXb9QoBeJiEPDU++qQC36ix5
0QAQgBawOSLLfQG2NPybuVaIKKPXtMmlvwHx8JAXrZbZ49X610cP97wiEHCXMdIOIh4oB9yNyiWG
p67cahnG2eAdBPtV/tKqyaLwuORb+GdN83WfwDIrT4IpVdr71IsJiVA5kcrctrdIuxc9gapfhimQ
hGL2WvvvQHoqgMh7p7V1xH5OeIoUxndsoah7UqO/LIT/IuTgRt5yfuRKph3JEmxu04N/dDnQ9T1B
eNazX5SXt8e1c7pGXvs9kc4UaJcXSM3lkv1M0aohU5+DaMWcEmCVnx5crJvhqCWolR+9GZACp8tw
QNjDq9pqlGxHXJYDCtp1X0LeLwXklRE3hlnlr8t3fP3IfmYnCUEXsF8lp6j0iwIwAXL296GdR7hs
zmYkPnLIE1psRcxLuDkerh4wIhTnoakmM0aPsMMhmFB/j5Osy8x4V9Nzt+yJOvVlt6iSMl3o0Amp
e0svVXsI27ohJlQ8jU0AGdhgZ+Cwb9dBK9IOlH7fk0m6sMqbw3Oef+ilMrMKOF9y0Y39dNST71wG
gRNh/AUM6+CP7qnGX/y0iHqZGMcsELsut5GggfDRTfgLeCo4XpnpkUX1lr1QrED2xhfKP/YAZAnk
wQuXj+SXoMISewnxPIHo/nog2xkHDDWB5JDMkxg5aMuZkg6ewHOayP6mUU8jw3Gm4sBoPRUejjMM
ubou4UuxXjnBeNfD53L4iy13wnSb+xW1JT/04nWHESTkoSNl9/rgcs0ld13TPZuLED1EQEqV1SjB
swr+5M8GIkkbqqMyhUO5XFegqFPolRk6s5P1q9VMfiSv0A9T71esnHfDWhqcUL03OjuXN2D681qO
lqSDEZ2wowCQA7ClWy7bwkTVuS1PZIcjNfRIOQCOjcuz4KCVtPMvbJBkkfyC37TWE7+H92J6kchD
qAUmGBOPhOcr90QcvFiuC+Ao8rDGveGUTN2Oi+WKFkNI8qjQZ8X4YhtLYCDsQIPOupVqop4XVTrM
L9z+JDYEeu3nnFUj8jY0LFbRwT1h1E7bxu9qzhT3LvzQy+xerCglSFpBZ0Kmye1y6Lk0zniqXy+7
9+F/ZWw6ZVeq8z8xsFujMmr9kSPph121RLlTwy5l5FzBYJny3eOlVRZaRuMFq1JF8iSwBreZpLhm
2rL5R5kaoRAAHzDMLi7i32NV9aBhEyCBymbzc60NqxblLGa6U5B39HFEnWoiLsD5t2HKxvoGxcjY
z32l1F8J2QQpdu4yazVmKKiDWm8MffdDCMP40BWyJfBhKq9ZqZRbhMgpyzvBN1+bx0UdINE6utJL
tMVMuLH1Tm8kjuMJhrSao2WD7uVxfwVLCdgVB9Gxbr/Z7rCMDFQs5Y84ol9bcIVk4Y3FwgGN2hFF
b6fqBKCcCTMKomxffnF5ATuqmy11gGeZLCxM2cKSji+SgFXCiJDguiyyo55a6kz91W2rJi5UcfPV
xijTqGkEwUFTwT3N8jbL5AMeD7R6nT/tfGULfY5s9UE5E4+lCUIgkl3182krjCzWiKF+RGIIFKSP
iAB8M4rZwrzhIz9dbLzBC7fB6wgS6Op+kyv6d3IjBazxdN0laCJQSUlT7z9Afd0D0y9jHhx8Yfwm
BbdARlgtVaD4fuiszLP2GHYxXfkGU7n3YTzQCpLWSrq05Kfq7AsME0lbtjghPPPgmKIIsPVeuX7C
IqwJKF9udQ0kwRjCddkpyOEzvq+NM42143KIxm7V0Cg2N61+qm7E+11QbVUJodYocMBtZUsTEanc
jNPa0F3liXoV0jCSGYCQSZMGRF36a1yhRRPgcie4ojFTCgYjdUNsstwk0Zy7wYZ0GGUV7UWD0A1I
1DT2GtdyQasu9hAmkgPCYoP4b8HChUiNQ3Q2v9aDki2rvS14WxygvEBYxK3Zc6IxLAGSfu3iRCk0
2jWTZn3swqwjvbThbFEFqpzbCk/uzEvzM/HSZafq5ItSdS2M5Sp4kA2MIZmpih87J6H0ADMfwc4S
TqiOtcUpDMtvu0xK2GlKyQedgBzDUI9UN1bkQQ/ZyBopNEdyO6uMh2pj06NZRVAWjN36A5cSJdCL
cJFYPbyaEiedQK1aLgcRPZvA31efr/9kc8g7UgqzJ3j31EqHsZaumSUhz6f0ll7CDRbGTS9wW/ll
1s7gc/KFsXJVtuRk/smZvMEw+kcrsRlBR3jPo4v4JkTNkD7Ay1k4cFgBqZyyUgnDHqb2+iVXzT+1
83nwe40/IiqQe9MWb9ttXND3LVIrHv+R7BSEJXUmyq7/0l6tkjyPQhMtBZrG7/WbaASlR0dvNSH9
BWrIhgQj7a65MvS45sH5wuEEOs7uWyQcFiudz9jhW2GyKV9In/eIh2xQQlC+TJYMHyY3v8BqYoWd
jSYcBoCVs0/ECOqk73MPYOpF8EhRy6L0c0RAEpkH/TF8nolhfcPFyNhQ4OOQeAM7+Vocgp/2POGz
QU+c3xcf/8mOPbj8guwzgFhioZKsFHNMXG4ogX79UrZzA2yQN7fxewkUU1HHXY+fULarNHvCZvS4
8dMmy3Zykg2USLsCtNFnEv+0evd3f5V1UlBANvrZ95+46qK9AVU6fzbUpFQyEc/7FjQn2UK7Z2Cr
NfuejHvcdceGLoJbbfeIaN0fki3yL5yEAHP71PMwJ80PK6+MxtnkWge52MRP3WiiZ1xe7fRAf7hA
QlZB3rZy09TQrHH+LtS/ZRIQbqI5XKytvQhMSzN42w/Egik9OJeHqQ/YrhF2jXLiEaBc7eqD/ifZ
0twpn6zdQOYeSG9D6vz+XamyQY2P+9Enw9kpxigzEvHP/6iIF8Lsbo5Qn4h4P89sF1Q2c/ImYDll
hbUEeqgHg43zpV6ing3l7Zd3Au90WcHvz0HPorKWj2LjZK00tWOKMzIohIwPjLMxheW+NxwIYFmh
Eo/lfD0/F6Trhm1Zb42E4q5AisMLTshTUxsr128N/Yf9nqHsDJb0cM5fpZyE0bRyN84PvgAg0Cnk
5TTxv9t6PJW1FF5ujUauWaQebaqEUMwbCU01AazE7s6KtrcnnUFiD1IKFlnTyRX2/YwTR75bayeH
4dUByH3KXJdvZDbfbD7iTwkhJSNHuguotBaZQG/7fKBNSVPxjbKYIeblHD+ArN7olSTGW8Deh2MQ
VrDet1X2D0yzcjOqLas7f6ywSyWRNgaqRsDBMZslnK62DlXyT4o+iNjnpylWg8XARZ0IKIsU/gcK
S77dIPuQqnU9H9IbQZDhShsP53e7tZ+BdVPF7JvSX3r8C5ZL/QIM/k89LceQIc82Te6PkAVR1dos
zSsY56lHo9NkLDDnZClFkBANQNmsBdJPPcfHeE8uNupYKP7StBQjkKsZdlZVxuSjmsTiw/1eq0NS
Vb04pPQ9QcW+sDnXQxM09gfjCM5nPeOcfXChimpJzxaX/306ebLWOcCvbawcvFCcIagEiM66uWQf
MT7mQpWUnSPa85InF3e+fVNVXslYar+2fyrbFFv+eqCS8NYHWa4l0oUFQa2Yz7SX5mbtLHgzFFbS
GNyfJvrj97AmlZnhMiOo2AZkQMu9RXbee5BRq/0wQonVKwGf/0vV0MzkB5SqeW50iglLgu8eBKer
QHMoJgkOQ17pQ+Cm6Mr8/Y1e85dvxvRriRuMFztZO3DrEwMeCY/+3zujdQEuBaCM49B9sFEmfH9w
9AP+baJw2i3j+a7xi3Vv+ihSBta5+lsPUoisqOEJ9B6mqtqJPmPMjcInL9eydfB53JQ9fBS8UX9l
THvn2H+5VQDMswHDTYNFfcIZ/g4EyhulzKWhQ3u3KYKRXbBLDE2N3rl/kkbqoeKv8wenLret1wWj
bfqwkjnyM0sGmZispfvjojopwCo2ZWotucCRRjr+kyX+0o8PKm6/UKS4VagOw1H0EWzPv6tUPiEU
tSd+KwS7QtJ3/fwE+71yBdDgm0Jkr94tSL2WsiTdN65zRTQKzpeZkkze3v384aM95N8XzsF4BZlL
G/bUaZeQokEpn49yxsAtGoAWigz35zzQSWal0sULeiOjdjsFPEcoaciRs4ShwLTCBvdEs1OrhDOW
UF6FIoR6GomjZLfG1fcGHrmN26YaMzvy/sRWVqeTquNCTtGUWduHJ5rSNLKgjV9c3zujifMTQ30b
8v+7OQEEskPNyX45gDP7RSDwmFW5gO+GBEFydVAV4ncwuLENO7Hj4Rz5FF5wPvsa6S2rv5xn99vf
jH3Qf9OX3kUjyXD0bC/0X7hxptLiqxgY7qjt8qhXsookqk28lQ+2m2akxWcahpWVVptDBvGoW9y5
tNgn9zMAGlMPrPkjjtCZOto2E0upLEt/puxQBRSZdR3qaDNA7DR7+te5ebU8h6Ih+IHzV+WLMqD5
V0HtccRYxUenGHEqOxGOJLzzpymQQML+Hb18TVtQ48VCeDUGUrIody4k25J18su2EwU5FkWkKbl0
izBMllbY7SUydsE5Lcp+gnuo0DojHwZajqIWg+aGCSXu9Z0RxoHGT8lkObVjG7W9nbTOfAVcATiP
1TqUx2VZ9Dr7J9AbMpibZqtvV8QRahFL8KnjxzQXT438G1Joh0CHYHVF4D2lShHU7YHnsFMDMoaq
wyj+PSHyPcVwD/gtdTjXlvIb5leslOZ2HwLdHgYLMJx4DLtdogm+b+Ck0f5qFbDhX/ZKQTRutFrj
R/FRZQRn006BQbZvjiYVgzwA8D3u4pXF6bz6fH6Tuh7N+nwuAbyWPBG1+AhPiiuW2dhOeTvsSrL3
czIbCN8z/4ENydSeKnOk+ExEmz94RiEU98v98g5fTlVkiG0T8sRrmQophEGp+g/LENz8jPLrDVNG
5m/OAIz4dLC6/nLsqXmjDTgtH0WlLAZuyLSwfVBMOyTB+MIAL0eWozxYv9WUc01fI46Z4ZB7qnCg
4U4I4UlYwlj1KqDaWyW7tZfbEaMd3P2zjwP4Vmk5++I2lix9enEF+Pnk/bQu4VGivYtuUiAszUSr
2t74EeOIJhtIznXRi7P24pFEpVap/JlI2K8zeqmmTraG3J7+YUBCoT36f/DKWAdIn02JyWAFHdik
UOsTHAkJJdOIuGhQ0lPl25qKy8jb7zlbbmVUkBJvAbaJXpBhqlVvtk43gXxXnXCwRlcBNyBGQxam
/y/qdgpY7KJGOxEawMzmM1DRF7jDfkp9boW+0HCBgbLefpDA/+R89dUpCNbw2QKp7t/v3AuOyIEf
GIxv5ym5s8mbnZpGrxubju+7vr6t7IdUgc4WMcW+aOwr6Uz/3AOMlu95YytBDy9yXcjGN9WsLWEw
oRNIz9PblojY9J5hDpj/8yNwHXk2wpKaAMdjHTWQsYnxtawF8C8sR7YsyiyMMKtrRX4I43/RMO9r
cfByZHe/y50cCc2skVnWeQCk3X+T7vkjSHNfc1VbAA+FQ10El61kCkhHYQHxrMiYuwRkp05WyoF8
W0QDpuwPl3Ay6UCH73BLvOjg4b/lfnOZwSQAWhBIVPhG2kmKFStCO+VBUpbzaXGM9WYY5HJN+LDw
OuPY237b/SBnC5d4sCLeZzrNU8FQp/FRaU7aeZoVw89ztw9jo4m8vmg7zGVeuECp+o/JeVRgavm0
BOuhHdiwqDZesz9qPo0XooeN6WrHPrIF2wkfo17qAel6b8ftIdzcMPW2zp52WXabJbSEPBJ08OPB
fsyx50671MxfCFlt2ge7bcaXG92M9MXLWTKgn6ZQ6MElhb5lhFiNjIVeVdcpjkWpKt0VJjQyqfXn
gzXZTuzPophD8zf1wKV1/Tc3ukr+2H68wOpVy0eM8gTZYGbk/0D+9jIepq9CkGvT5cThwVazyb/h
gi1oJMMaOGiwdthBS5XuU8dkwhp+1pBHXOm4cKJnqzMsu9PD/Bul7QuQccuTURTdm+Y2eR5bfpSd
TKshe8yC9WFMQOI37gmNwM/29Yxs6FvWTlwAOXvJypE86CB0ulYf3jkXhnmrBmJBt31jsmOlqkJt
yWULtvpIz6ucY9lWWylgCOeM6+ulYLXJOdgEYPkn648a4DSITg34f9VtDRezyqnYmRcOE1MdskXu
t1q1d+ZXGGybMnfgrm3lfOWwAHM4UJuH3foj6s7j1iwGX8mPfv4G7fAVWogm35IKjeMzjgLq+Ovh
qbeI+vlkmmM1BF3MADTzfxwbDgwNiXmXKE62YArn+e/zuirAh8oXQ//AU2lKJTsxAY4sgIwVFiRR
LaBR/KG6sXBMR2ndlVpFF5ss5IzoUiUlxOY8VIJ6s3rJVfyBnE2IzX4K4yPkBUFxjJeELy0TXkIH
9GZg5lVO5O2XRHEjzUR4EMYYi0u/iGVHcBDSQa7eF+iJi9w8xvm/zcyJl2boAi/eKtJGg6lOFMJT
gR79zuNC8v1Q3Zfu9U+NrYGpvORMR5w3ev1MnZdMLyzceksvk/ODhw357/1g1HV/1iuMbAmQ5Ywb
I/JYzreex5l2P5xKox/IrgHnrbFXAMaWnP6e2cplKK+zjBf7hBpDIirgJpNBjT+xYjhl9tBgbTvU
S1+FcX0uXfUxXU1PCV4AseZXyfbcn7raggmcbD83eYD19MTdXN356IJLx0q7a81gBiYinP/ZrwjH
sRGidwss4Y2n1JjXJwkrW2DHsqp5evstJaKkghw5VAMvTajZquSyBFTDt35MdNHsVdUJcunUdWpL
jkmAyLLZWIbVz8ol8Wic0436W22I38GQ1puqosTgGIVfECZHwt8nf4A8vXyb4N668512hprByRLm
5jntFBt5Zl8yaueUQWutb7jt61jiqmw3vFxVYiQQjWJAlskXnbG35mBT/XVWNdaCY4oUCZQyWEwF
zrVfZ4gVDGCwK8gq0LcHVAg6dZ2TAX0ldqwQ7+ekH2G3+bsvlTnXZGFf7HONRjOIo2sfyAwcjQ1v
66VJ16zq5oxSpIm6+jwd8cCCL1PXciWkpM8q/r3N8DEdAiBubi0s+xPFbhbjm3jtwXrKDak9NOJh
+3eXpkxZ+KWl1digB/n+191i/raJsvMGtU0X0eB2cbSPEDeScmY87RuTb2o8xK4fdJ+iDlMgt3iq
Bn6yacaj4/gkgwKg1iluFDhQZo3RLgBsYAiKuQ/h3PqBdo8gAbK98tx3Kb5NKUmy24QSS0xFb5vo
L1gr8uKN0//BsNf3/Y7AF8AAQYQuvprSvvMDRLcJ4e5wW3jue5sFJ0cGNwHkcDwxdhJDFcjr1auW
sIrlC3ubi8ADoy322v9OtBcTlxqpYhJwltllP/2+UFr8jGXf4ZDQ4uQsyNtp+y9Q61hpdkJO/Mbc
J+wt4gmw5MMqjK/n1L99d/8zZZLlDG+rZy1CDOEbLvza7EHG1y2Od0fjoXDjKhQktZYnG7zTwSKQ
5LFzG5G3bDjTN+1C6pYMK0wTd6JQmqDn3j6l5mQN6lrw45qSyDvdXBx2VWhetge3aIrf14c554Da
fkfpLYdStfJJiZlZtJfo2+qVfS1433G8ti2QyZHyt0tV2kl3RErscpPSuabX8pysEZKsnpNUdo6u
u7pViLkkmVKg7gJXrRXUILJNgH5TnERLmHLnmLxQv5exicIO/aueYSuAf37BMwEeoB9pUclPSy9N
vtZRaSNX7uzETa434QDhGMoGjgKkgXLRa8M8uYsAEXYbpFlG6ioANMRVKXfamK5Uzx2CueuJHlnk
l1A/vxlQeq3HRD0YblluPPFek60j+De/lSMDG5RQjNuw0eaJv2d1kMlbY+b8mhoQRccnHXIXZYLd
1m9P3hYoVXAAkG+s9fDT7j799gnSAgY0DraZnsaGiWP3cb+sIUk51je2zCetgofjBqzmMJ/cTko2
PGpYCOHodpeCmgEjNoOT23eALAFC264eiDAiexxj7PpyKbcekhArWLi7HvU6sKzhao7/VvSw16OU
SXzpkW4sSviH7QxaOAyWvWCJW6WDinLiX3Sm6ShxlzG90VXqcaSgEPpK6F1NsoEgqnwMdGajkP4U
xWv+c43ZP2oyqD71vjAUgase1Z6PAye7+PTMckBMZXFEKSHE/r9FWoo5rMwhbkmnMRt2bmprESGb
6LkC15XVcwGHVt26m8MaB3jDphCWWvAg0nrCvn0C2NJeyzUz0eRiMFm2GybDIe+QKk8z62cC3+ev
ppAnkmPdv1+JxJQCTu8zPq+h9ShKqHTX0wlyXrzvVom56uiU9c9JE9eCUtJdx1ZH8Gys+FGhJDyw
zlVffJkYGSKrWgOdXkjtn2EwueX+08fqYpgqZwgR9fBOw+8IepIPRo0j11pnexGQ1QrGJkTbS7xm
VRXRoVW/F0gUENg2qt6/8LxzC0jua2RRjv+27WlWSDB7aHrX93nDMJgvNqOhuYr7Aeh/t1i2gaKD
0k0AvSCkvUqy0dwjDWg31TIo0WQBzkjIrZPzp6gs8N0fJg4xPOzrnhp9OfVJsp5AX1L3YMvIWWQ4
QDJfbQ1KGa6GxigiKwjp32Wmn9eOBNNbRi1PU12ZUC/j7VMDMcwYNacaKK5qRlUV9UbNqg0mngHR
G66DKgz9gr8/Ikc43d6e6oHNgcg8jbxWIVgyYdBJerwWSLXz6a72JFDfaDKL7ew9Qa7A5xsLVzs1
wxRclzqoGSZ/VyUWrIZUyhLss5Ybt7GKqLDaLsc/T3KvmZBbxF8srC5NwZtgb07QsNyLAJnGeLxC
LWzvdHJV6nEGOatTyPibZmXEqGDBob4SruUbA8tHIVFm+4Myn+ilyAQoYkDPILJUL5aLr66f+t5y
3yQQa27rB3H8tuy/HFXS5v6OvYzXwZJluLU1ZSl9LcUgEiwEVy6EegSK4TsnNJvuDbAVm1d8K9s2
M+QqCEE1N3FfVgZ6DWWXMS2RYC1/3Fv24Oh1oitS85t0N78KyszCn4nsB0oMXcEH/7E94FT8qp7i
Hi9QLkqzFNH3iFIdEZwJ1GwMc+NJwB/H9LiFFV/IIqr0EblzUdW5ioo+ApP4PIrA+6Hxq9Hwh6zz
q2OvV6AhuzO5xqrZ50XL/cbnW+K+QgtxbqWhCD78SaBIoYR1akcIUA9oFnsGHQL7XBYZPelLX8hI
biKKfOC3wY0a+J53xeMnzHk7EpcSzyES96tf7MUsUqKok1MG7nzBtIb3iWHnijmevYkVlxNvWNlA
fxJLW9V1qegUFkoyU33xw70AudQx1BA1DFikaALZRABhOj6yaBOnSEMM0O6enPyZJe3TS6XYys6p
L1wAFN+2XcqKYscTP6AjOrZBZgrQsKpEYC6oVhuPqqtUpGaQYkcsJP5t3fBa3YhbqQ0OY8xzHDNk
F6U0bK29PA34ACKy5VONY7rn3FzqnmlT9ZID1chR0iR+25/joLHAzFazaHToaEt+J5eTIUD1wSFP
iSn0vyWz9FK1QQcZZpMm/XSczJL6a+21J0e3e1qcgGzTCvtQGKd0QCI17q8OBhqbe/7h5pg4mo8c
S2LrmMwKkD8DATiuRtZr7wU0sobh3Qc3KiBXLAupQrLtPRcUqHY9XHqnH/42FWnDBHxryXEus1XY
E8h3fm1oad8icJkvnfuztbY7MMc8FxkG8aF+FRBDSd7oy2xeNYBQVe2SMZ/DMwYDqowS0cGVMMJC
KYXzh1r+MXi8TfHoms5Wr8+1RGWbgbE71frrDTztUB3ldwgHPe7k7Jx7om88ow5+vZy6ZhLHpPx8
KFrvVJl+0DGNIhdpgK7a+Hb2mzIigljtojEClX0GEF2Zm1RjiOfyG23SdpYVMVWsoBNVHwVds664
Z2S9/8LE1feXumYNlYsDBs7jPpCpJQtBezcA8oE1RvMO65eVvmG/vQAjWnEZS87iKZs2uMa003vJ
qO7wiLrK5atOUsxIgz91mVaNt/xDYH4HBBxgwJlsCTm2l6x3YiZ7s6z+7oSo1PlIFjdkk4A3oo/h
DRQwAtvAaB7t+JbXJMcEj/cFV15Abw0AlB5423cOhCkDYUNyDxiuO4TTpzAWSPArfb23vLqEbvSd
SPJj5fY4MhojC0gLq37p/IIRYB6Fnkwwlvh/RzUwffdZCYLigJxcac1eD/9DqfTAnPr9tedJMEGJ
M0TbPJsJ7Wz8Rvp+uWGHVFR9AlQmADwQCSHxXs/2BuEV0Y0dGNA5plscdS1CMRbAJ0fuUbquaG96
ELI3EaYpPYYlTVOhICQ7NNN9YYljcqzvxdS0fu9W2NWsh56p0qYs7EUUn5gCcgfA5Dq+c5zJJCnx
lVaaYLQY1lHkLByBdMRvfvkD1nDxMX3q6jSUqZflv7Fb0vjCF6Zunle2YFSIn7ZiTtQKUgTFSJGk
vebhy5Qo3BpGblQ8DNP6TsGkBJzdgyEJNRRoaxaHbiEuEi0u0Dy4v4Z+w8zCcE2YYsW6H7GWYEMz
wLWrxoEsB1CUJEgoeZvLkfnd1pvgi+4mynQPvkm4uPtV+qgSGTIYLw2eybLOrGbK6J60dsih4UEM
3rQeDKrTJ2fpAy97kiX6ZNUN89u9e8PZD/l2Qw/Vw7ugbzvmDLWRRTQFkQ+3wLGORV3dDV0aMJxX
E4E9lHk570sTAZEHbyGg7TlfKVRUpPSF39I9SGGVMlJrVupk537G0EEkDNki/5nhSWAj3kkjy9zi
KmG+mMgdayqhQLrTna25mJ9QluPJwQdIRoLkWNhz0mmRCLofGanH243YynXfGM468/24tYBb5ia/
sfO2umPOlxqWb3aPp1zdWS3ZTJe9nDC48CnD06GqUN9OYddvLdpBlnbYSA5ertVC31nVeY1/0KT8
D1kZjE7bgm1QO5GN/uL6Gm2yu1WuCOm86zv/uePWO2XxwBI2lSHigaL9658tFUAYXYzCpD0SpnNU
h7CA2hEFeDK9ev6hnUcPc22/mY22F80iZuLYQmuIMipG/lFH+Y2QS8P4GUCdbpjcBmUrMVBO5Nrn
ThOZuqt+E6zki3JJZR3X1BrAmaKA+bl3jBH5Uc6ECzwmhDkYH1FfYbYOWiJjFh2blB+1VHzvNMre
JKPrImTJzzSrBBT2U51ni1ERxBnGMm6tUN++tnfjfbnceM/UIdiOnQesHKgxjh+wvxFuxZSZ6QMk
HXRDd4Mf/0GKFuLTJlytbgRhFSAPnzqHMu83gWJWh4ZrN/7mU2mGJJWS6UzhLK8xcZWbodp84E4L
L9uLj5iGvx3bmEwAJDY5K4pyFmN50p5ayUOW58zCZK8/1BSPFU/ZbWekKSdaE4XEuKyilnFjJTva
ysw1rQDhl0Aaz89uGeV38VxlJRhql3mFKi4rXDbB6Kp7HGRNmtl+XZA/nXrsBXPSHG18TRAoLTFG
3smviuCNoXlSVanIQzUxaoFsA4fbnQamdutfaB9WLYs37a4KzEDyNFkG3m+ks7iHeqXb+rbp9MbB
3tGDOGQ5Ud4P26ccOnH538xMk51YzT780KILBBwfs3d5jYG7MVqI0nrCas2jdpjhZp8NIptuyLgr
hkgRp8PHLIMAoAmSivIqZ8nHglOeQNjB/CKk9le+svRn42oMH4bXm0WM7FJo1lUtVczfeN/p04Ay
cGoBrciDcrpM+7SdZQFu4oFxWGI4ni/jyGCQ423L9CwBRdUQuSOcLFbrApIsNUEvAZL4qyYa5l7j
X9TXJHQ5EAoxBMqvm5Rw80i/lsSe7wp8QmngfueLh6V3Heeof70x8TJj+4it0okK/KYupQHta6Sb
nnkInRnnX2emiw2RC2swvsiJ42iHiLKiqNewARzhCIh74QHozaw8LK2u00qU8yi32Elpv5mnXqeW
ZewBppw+J1g2ltTfbMJTLo30SU24mXg6JMLWdgLKIBtdh1alFSkcXLX1U1GVkI/+I0OTfGMhtWxJ
QOEIwFGUt1VSoENEV7T4t3kswjz8+G9CO3j2dDkIJ4U6fqaYfzKTvDuI6R7VqTiNradQaehSdNqa
639ntRJakNyb1xGun3oRL9eP0zZZFmUSbumT4+l6JHHo+btNvVWBkGJbAHjINZchZgJ0gowIXh6E
4XzUR1SqULlERJs009zQiTwbXDUpCRzIDI3iXOIbyuU8TDoQrxMZVwnmoapMsIVVljRx2xLkVrnK
Lmtjx2UWFc/zMZa3TbuxUjt7E2Rk5PMgKodF6LjhbxIHxNM2RAEFerLQX0dMC8gsmQTlwGGgc0G7
0Zd/4RKBVcpz5AKldhrNwFcYx+ycowFaLfds2njGXRqh+BanHcm3t7OTYp1/T8ecdNDHVS92w6w2
zbaD2Pkhe6ZLbvlaNQCcRQLhQJN6E3UFGpZm6KwxsBGHGun36cTKEqK7md3XREHxNyogqGQ7PUNh
/3JT1bbrxozkrgD+y0uMezcQTHpDVnwgtGv/AgNfkyobn5uSuIzsVRDdF/4qyqxjzG/EZ8NmIiFf
F0+CHCtd0imYPmrGRTtKpQ+3N8MOqHsZpdbSd5KyBGKW9pm31BRd50hHpSSd7BJ6Y4SVLb+yVB8O
a3vxuYs2NbxLCP7V+9FN/BL38AdsDBCx2Cvhr1vQDdYNkQq2wY+EEIK6iVJvi44Wmlv9IMPRwe02
73N4+Tg47kvVW0UxeuSpGqfBcktDD8GYbw6ekrnS2do/1JOqs0MVuy3YzUYEJ8N+4x7HIlTQ9L6/
hVcqlAtD39KfSjIfDzewq/taYUVvo40JSwQVseb9x4GC3ZKGupfFAYBCslhdYmRvYS1LMZtOiq5o
FGKvdk9BHBf0z/2Z1XBgs3g7sRNuhoYpYLAmU4AVpNqLMXVLBSg8PWNSydQMHwg/kJCOclSTnkBA
DBJ8bKupv/GNWYnFwfvpiIBpNKDB+xu6N2VbR1Ia0eX+6E6XTPoHL8nkVwXGMtJ5ACO4cAEvFHcn
GqZrawbtTigbnaqzlpmi1eOBqSx7jWRGsL3jWf3yoyUM3n9pPjPLwqoBRd3LiL+oSBzRt2jHo27f
rPqgur9jAe4LB9xJcVG1YkGatb15Z2uTQooJlW2NKm13rgb28y35Rw/ZrVOokS/wfM2Ffepa1ScF
8xy5E12tOGLzTGs7nCYx8zbN2N6Igwsy7lxMa6pkVdMxUf3wuoyIZa08SIlFKW9nPvBkTh84aYIq
88Erwe94+TNK08/G0PbTsWQK/W7GfYrr2MeDb4pV9IWZ0FMDepJXyoouXZaH2pYmZeAdpP0luWQZ
YgGuGeaRvmebJdQpSDYPHXFBXcpZW6+xPo1ZdAgqywxK+uc6PMu/nJti1l0nVKQc2l1KPdCny7EM
+S79MMB5bMirs+z5EW/vURubOsVdnfm1NGzgGsl6X99FLUkf1zAFbMN0dceU4IDNT6Myw6VkaAq5
6shleRHNL5muVI5sRIBFYJUosvLwzo7mLtTmpF/+lB6I0AQ/exe0gs5PGWFTYQIVx6LKrb6F1C+h
ROxFCpNu4Xukv2cJ665fxysMMocWupjq9M3wwZTEH0xvs0R/1UurldSmkCytrErniyZomck6F4lh
ftW8eM6a6SU1s65je4WgmJngjsM8aZQT6hHfF7rc3IW1l4DANwF/keU5NPcvOgTtljDa4H7QK5nu
3id/beZtThIO4QFeCXUqNEMKlex/xegvmZBRq+U+1ioaNhopjUswsMS5rKAnWdvE/4r/hy+Si2iT
18RYTGVdrSD8LYP+PNJJ02ifGwy7wsfFYvhRIyZ4HsVH4oB9gWBu4PjEB+sfyksEkejbtd1AUY9N
HH5jw2mz/+Fjr7b3Elio6R+hn/Lq0PsuF1i9F3FJKTqm3HD75yfcERcYjciH8vMjYiJ+D+abdcCz
+W/+KsgZ6H2Z2oPN8DGDj9uV69guMixzsMy3HEIRpX91vC8ic4h5PaVqLajnBPG29ABD8zufYWvx
yJDlViHz95AnrfP6VtOlLMG4P73JLnyBcjjHtiC37YetR9IvYqYcDkrNSZ7k8R5RIOnP89lZyh2I
Qj8zB4Adln1sJH3RA6//izUM23BTB2Njby73QhvAz3ad7yxFBXiBJf7I/DLWiWbLArpW8htB+O+8
4zpE6mtrJ+PCfBcfdvB9J+774DwPz5KYoF7p72JXL2Ply5+95CN4I7zsV6SrKU09Hu76aXHhnkWX
SV5ua+AovL9uN8ePeLoc1CLaHqMQ6cORP/HCSCWBwjHhZHNunwit2B8QX9lnF3jkVCotA4qFaYOc
NcPZBCMcYZjgqP//UTL/LHrSrUv85/Z4OyJ7amXRWlQR0+8lIhCjK4jb5qscWSYpFDl7nQ2Mq5Dq
XRt7tIwsWz8WNuPt135MiO6iYnyay8JTvd0KRqNVFm2OK9jQ9KrczVls+vOPCHg64TNiTpsZTQ9v
O40n/N3KNkYAbpoD2KurdgYy0RCz3wrMUZD9XGEw2XbvGXAXy50BtTcRAduiYQ6PJGztBURVjklY
tXwAtCWNEEBV8NUpqfzqy/rul/oCYX2gNG2h8pklt93+RTG8EX+ErtvQEKh38QabLYwS+eeaLREw
hK0r//gy48VVFCiaveP5valZKW5AFWaxt+OciejKf5uksGrrgGeXF4G9nUQZ1xkiFQ0mtzDE5R08
KiBFybznTIWxdj9RUDw5o0Shl1btOqd6e4N4lc3MYEHP2PE0LMxFL8ntePGOIDEk048Zq+0u0J48
m2y5DVMd/sFSaj7xO0o14V4NFG4/1keIBsTB5JIOmGJjF6GatWqTw48AAsuAvuDaw+Px8IYtxgOm
glr2EuzQ4OPAcIw3zKqxIwiVDvyFT0vuLqSEhOLlsr9tU9K0q7id71o7vceBsIspO2NwkULQR7wY
rrBGK0H1ewmtE+qG6eUpOC7yE6vFdmHoFQd9c/5NnQsDtcj5+cpRfAerhqWMOZ6or5+GtVwDQXyj
zAUSFezDWOayj5lZ9ZV1o6jwDv2rBo+FCIp9j9yzJQjo6v2rullUGh8go2g9uPFdf2kt2n2iaTKe
IjnFEzOsCn5pxmH/NB8H1BmYgWgcMu7Qy5d/sicGjqxcByxf4ePc8SherlqnO7GXsRiyyY8pJ9W8
quv+CwPJbsleczsiTubGsYHrRypRjHFSt1IZP/wg0eI6Z4VQ9JQIhHq7Mk6atDivS5FrNXWwC9TD
SyhWt/BjN2D4ULoR6wRqMG+AWX6t56cdjn2aedTDEdiW27uqCx/ZXyJZEwMvXV5Uu/hFoSpUyaB7
S8YN/pvXUc8X16V/hvxezTaWeU3G+ANbrh4yVPN0tSNsgsqd+Kuh0FqbG1MN97tSsbjjESD9+PHa
iIfUd6s61kaHX0ffTHS99Gjl6KyqwRqRs/C6YLD/tCBxQ/oWxDRkNbaYXPhm/RSOVY0Gb+/pXd6O
EuyZAyIa095of877a+IauIOs/BOHh86Q9TFop6/WHC0HmChuUDZMi3IvBlojFMFnwMgjXxcGp6je
T1qH9hUaBILb2vCnrRiiV0CiPX6M8z02zBARLV/Tu5/rzhY5faGJm4gnGG0RwyefuqjXhlv3Be28
UzI9Ipw40SDyRoNoMqrS5kxAkBVUWNRiS5iSIstD/I2FqcJ0RM0SKo4alLgZkby1shK9MLARRHKb
OljNwE8DS6QJ/VhUr58qo4pSjB4QbwGVkyrgso4Ym9/povYjwIPSuo01g3Kn/gVkNsHayZZFf46x
chPBoQj20BDoQqB4IODW+yoKrCh0bGEJ4XnESciNTmFyD0MEavkwlXfaYey4fJzS4kLzr5vSVbYh
riNlxb0BLu3w1b802vadkV2L3A5ttcAWEzJSBnl6oZZPMrZi+pSgGGrua9sVgsrsYJshRICEnPno
zxXys2HVHjEclkYf9ZSU5+AK/q+HVArk/LtVZ4sKYSCyn4+myiyQVQQhDjVjw6nFSRWo1pwIBxuT
FoEoDcU7Q/CDwgVKRpjm+lAH3fEja/HLzoaLQCHnM/uaw6ERx6XiHAoqymAhDPKhp/BMLtmGRYNk
1ZxuTCdvJWmJskmwpQbT0F35RWdeJa+LL5Zr++TN68yDYFqAqahu/BuNC39kYf9X19I4mKoe3QUt
V46kT6g4YV8Z8JcPXtYeILaXdceNIjrvhMG5vgwJD5RxZx+sNKDvfxuVcnU1v1vCB2nJVFSWXuGt
huZVfuwSawKbaFBA1BMbb1UgJlfsYSmRaXAtv2Si8gDhMMS3s1HTJMbWSmFilDgIKD7bzyYcGhXA
RsCrZzvJEhRvr3ESDeLo5JPeKtWBcfR/QcCpnpFELoLHOL1PX+oLJbvWNXbb/xGlp2UOA2kszl4R
aZsOk3zRB9yHhDgXa8Bg05YYMiVUS6TFZo7YmDWRo9F65EHQ8UXn47rQo+BSdBYAijcavQsQfJNU
M1faugCwmo7iN6RL8+HkV8PCeAXWCflGTSV4A+C2/dfwk99n5dYwhjPmEXM7RTMSgZP/ZsSucuMG
vxcpfUhUYbx1rtodQuwNSadC6qFsuZ3UajN0TxDiXqzr66jhDIaLUcO8cc+WjkT80ssAnNmgNkTe
NzQ0BsK34QGsiseVAlGJl9Bh+3rmeO0g/+dCE8FKV9Eimu8Hz4DTQep2YVuHixOY79BjMj/XLCQC
+6MM8pT4jVYhN4ad7o0v+nyv5YyIn1wnaQwpndWub5C+GmusTIPH6Q7bbE3C6G4hR8jwkhsmh0l2
RDtXBs69tzHSOlM4pjA9xeLO2oCgymRf3fitl1DEMzCiaPVHHuj7yD5hySdhTbJacNq1Wqkwflq/
qY6sYt/1Ut6j4p6DwvfY68r1PCaxQBysvezSeWxjc4511O4vmqH/QHxST0Jy5zOdFu9r3w6yw6zr
kWMawDKwk2yAxtAmJtzIL2P7N5+xF+CrZK5FOr62wT6aoOC3eujvNIV+kz854pLZHfI4wJMglNiA
Q/8Jp4VLi94pO+RjMQ+yzn4yErq0B2CWhipCZ+YY4fL+jPlNAYkaFLiwT9EIy3kK8/+RCPhzBfzI
JcM0/k28zZFC2lql3/p3wFrUfz6afpl54z7SL6T0JtjHtE6WCTsSvL2sdyvRcEI5mtTuVI49xGr/
nuBiHzQ83U9RyGN2G3khI/P8VUR47kro3M+FuiLoRjUwy7HteJx/7zlfBCTCjQPtOS+upY5peFAS
bb+Y6kPZC5iLVJj8TlZHSjOKeB266pyHlMncNaM1fpm3QH9Z25pUmq23gy8il9QElnxv/7sg/gL4
yY27jl4A5LChNTWTRVk7CaxgVtAzr4piNUQk81nUQEk13Lteticcgo+KmVQMTJh5X2ltWfdC7wfq
kGVvEx/lIOcn/omv90dxxN6s0KzsRMNFUcIkEZCed5Oh/l48lTBWPZi1uWNVYplmsyl7bfOpw6+s
czwSJE+S3L5bOcWnXarde/FEVMQvzg+vWYv1GM6dXDbP+qAm21K7qc+isg0EkBg9F/jQ+zphX+Ak
6l8iShnHGoMtyIhLVu4MSzT8C0Dw70YVx72J5/ejX+DXOpjVg0vyn9hCqBk6A/NdITf3ocPogRMo
aZBgRzxPL7+PrFvnG/7H0OzlsBSXLEB4mRMmXCkPmB86WyRTEk1uxjVqgvQLu+OlH7P0+0FZ+F9G
uavvhZyL+Y96GNFhppBSRKE0HITouJmmZbtBBxp8bIkTh3oladVd6nzBj+niZbT5V31m27cC1wwz
jRFdCqhaeZOQooA+ull3yRIvC9o86oikj25B5zV0jTUQvRZrIo0PCgaYdMpuMpa2ub96coXf4GJA
/ORkQLkNRamWd1y8QyX3RBDWhrZTOm6bntw6iGvlWSAzqzkldlsn//AgMNBagq3kQUsImfxp3e3F
XSfMGot/so/X8bhqTIUSkhrX1jxHCFEuFIBvaK+9mag2jETlebUkVrgLUb3K/A9xu3OdUolufiij
ZGYkzatuI3Fcgrhc01Le8eP2ljVm+JxWXvohrWfp6xapTUnIozGZSsMqUuEdywLgL9UXEJ8TPIDU
sCW8/OkdEq1BAADtEm/Lt4eWw2THEkcaeCxYn5Am7Fqfqu4zFF04R4XdZvnkNqSwY+aUWia31Tkb
DTosYE2Gra3uY1kI3zXhp+1boDwz+U4lGcOVl/aGtJs2Dd5RDMpWGQKHTPZAY8DoG9GlQ4pvfx2Z
M8mnv823eV6tMrEU7RiEUxcM9haAhS1klQKCyLpcrDOxrMCBP6q2MFXDVrDBBlMf4u++ljZTrq6k
kaABnG/LczE67K2WVKP2sycIMjEq1hoU9ZJ0NV5U0j7rYJMYihxKbttvmrG9FTSl6ePHGKlggCZb
8SaxcYjoXuWTkoYx4TSLjNXJ0aNkV0EP8wrRkubZqDQQBy/LK9DGOLv3MS2qKwmDKpAeU73PwWYe
wOuF52g1XqKBgyQEnSDO5N8QwSVrAlEI9J+yDzONBowp4mL9ueNoCK0FpVPRu25u23yt09uS9eXK
QuGDGgNDRB4eKDF6JD+4/xtGmuFgmrdxVTYxBn9B3NZtA9LPN6S02gtDi0ZZz6sUo5qobY9xu2m7
syiD5QtbwoiAYSByqfWAzedSQ8yCsFa16yWil3REazoUEWNhFGIWsZ3D8/vls/yvtmiaFTO+q6eo
DlyzMcXgMX25OEosAHslHnoMTtZ2JGhAbNH+QDXSrnAfPdv2wNU9cbNu2nkKuLF/kAm57KUl6O/z
EhmtHqlubr3dvvqmL5mbR+aB5YghOS0HEmNb6dJ8Vtv62UjIDz5mpTs//d+Zkq6trL386MMk6KSr
qb/hc4nY0mbwe1DGEw1ZjybqTIEdDlH2LNeq1DfsI5oORDy8KYFk8yp7gmcH/cR+XBLopd29VXjw
d0GcIbQRX+rcZwFGMyZ0JYiaMQ3Qh/tG9kqoCqdwQLpqjEhioqfOFxtn3BWnAz/t5+3L3F27wxBD
4wbqvU+kDjHIAY0r1JhusMOgO2HUZ19bIWRG79hfXH+lw+0VKaWPFRKulV6/LsBaUfpen8B5/IBe
++NTaftNzZimGBEdoQQd+5OGcd99cPheZ0umVx/ygtwNcUN2tx9byK4dqhHwCYRxEOFK0ATx61B6
DQQtFXYdMOaclpE5Ew0X8xlAUxw04BBCEK8LMBdvH3UISlaMPgDzAJ2pvb0boU6Fb2CwZXYfpduE
Xo/TOSI1bXF7EQB0obH+OpYNHmjku631B4uUGuPxjr/VLoPx5Cw0Vim2OlkVv/bMNi36UheIjnlC
gCXQGXC86p6+HXzqB4Y6EyoYYIGAjTJXeyu4/Foj97bMoxFJ1sh9Z2gUvhkDEk46CFm/j75sTb+6
nUiXDRp4hm/uLUfwGhW3RD4EBeihU2QBN3RgPqI+UI2kkIFj3naPgg9WPuKEseT2IhJ+DnwZmdwY
IeoNrmu/5kRiJj70N13GXoSi8mCCOf66YoCFItcZvyLr5+KRpYdtMX5Jb2fgRBnTHf1ydrSn1BiA
jtkJh1a7q3WfImhlRgyvqzxzjjuU8pi8BuMWVbLAYAE4WluydBjTw3YmZJbwlgHM7Tbvr09R3xJ3
L462S+hkKfz6kVP/QOwG/bdJ2RiBZPpgApoYw4xNan7RtAwTLcG5o2o83yM5p84kXmpfgrx9S1+m
VB5Ld6fLlKhiFQMYKZQ2skSODvyYS5RyCl/+nRet8HIXJUsXILAbym8tqv/gfG9/Us7tczepueKJ
FQZdDHWRO3PWGqV4aZux2UczecJYSwm6jawZLscTrhkBPaQZ+x0vPvYLLvXXk7cdR5NXvbHtT8/g
lB0ONqA/MWhcFa8PWoxlDkuwM6O7NRR+pylBr43xLAuN8Nd5NRPztBXPwf6UjD5VWEWi8Abf1aoh
wp7ojyaLQ3h5+oyKxPFf1cuWaxwj+mV0zW/Q4oJNd8glNy+m/3mUy48fQ5L4nzAkIf0Ut3IsQw1P
qXQr/OoXloYdBGmi1wLvUuzFC8GF2Xd279qRViQtEaqDYZWzx0HquXOv0ld6x6j7IXzZYYUmBiti
4SRza+0xryTGo+Y7dA4Z/h9Dc98LORfLAUKbFPQ2SbReJfW7CnAcxI5O4H3f41OZykMYHMBLtLNY
x+6xg4kfV9NK6aIiyrZXvCM3T6V90zUbcZMhZ+wyMHovNOaLXWrFjWpBi15EJmjmGI5kjNuCGVqi
qt6NK+oBG8yot9s22LC8+c217gffS4OmkFURoUZzv4bcIsvPwOLFVrGEggNPk5AKhlebooXePrKl
whEFsCqoQDXfORxm1TWf6iUhwb3m3Rja1rw8BbdOaqK/yYO26cvvc1oWTAcK6zZXZgF4eyBA9BHU
m6ATTUIcTPLgLXrxx10i26tYmi/+G+LTpDHfFzPh/IryauWVWS4PPQ63SLQHANwH+rcpjMJfwzcm
lOInuvptQaEiKV5fe9GikmiGAhGfXS2Oii84CPFRlXboyj75lahLevhkx4hH67qcxUVU9eeq1rvO
FTH7YuPggI5q6ZKKjehafzHJpyFnGKfToWv6wS3z0K8N7mn7/rsdyb2WAyEwDT7bEVcpb1KfMxHg
xfQRoH+2ldl0K0potKSrLCWvTryHMeV9HhofVXn7LRR6Q80VLulPsJt3KfG77UWzsOXRVlAbZIDP
edZimi7Z3Rb7ShizghEPwQa9pBMQCxEokTVQAawojT1s7H+tYBITmqIPu4gP5/IgbVbi1bBWorh2
dsFmmxvbZPTyHO4caqgjaOgKyFETJXWkQN9RJKIR/vQgq7+qEDq2QGU6PAI9dBUGmWN318QAqBKj
OR6jwH+kq2YL4je60Vgd/dx488PfExTfDzQoG5X0MqbeW1v/5eBg2Nke/zGhwuTH3TRvYrbKMc3w
K7vQGfmRVSvlxMdmpS9DBpRg8GP4FYsj+o4yMZSWRKgbnyg5+h4Xgy7nhadLeMg6b2C4YYCL7tQ6
1VZ5qxrRsekSuUqDrmNN90DoKV6B2AhPUW1L41DFJbVpKzSoyhi3F4KXeThs6TwGUe6wMJzoIj5e
nr9KZl21WvtKAIo5tiPFhI/LM49MFYd1Dw1Y5RaXsfM8mVil+rKNRVZ2F+CQv0WXgu4q/0ixGwcA
Usw3oUbsZsszhSbDhgva2UvVrzK7lQ9V4ovWByrfDjQhzlIDkEmKRJC1YNq35zcZev7e+RFSrFL4
+Z2pO/VNFUbmqBWT1nTtvWNGRdaSGY22npTYycEPoXJAaG2wNpFkvOoE4sAYv4Q4Wmzcx2vLCp4f
2FAs7I8OcZLZJ97fBoew7MX9cz4UR8blqBasbYNd2mEYEG0arvuRSGM7qXwxZ4gXYBc/NJbOqj58
Wi37MF1EUA2MzbYbwydSG/JtQCqu2dDWa6zFoyD2XR87RQ5bFXYltRjrV1p5tEXCBhFUyrjulVh1
BFS/inHuIsbBV3ci+9xqKgtQHtyNFuVPS8wOdsnSmzuTtVxPCbJbAnPAtOM0y9HCuBXhPS6eFIPG
vCnhv2eO3eHUWsldf7HBCoxnPzmhl4tvsE/avCd39VhdJmwGLbdkT78zBct9eZqnZ5cS7kfQITZ4
sFo/C7GgQKdEzDEhPasHS16j++d4JYPLunS2WVrBxwt+kCfDNgFtzlai8P0RMG3o9BsgHpWOR3jg
kpssEmisAwT+K8NWTY4a4iRhoxs6vJ6KIMxnd5HODFnGpWxjpXf8kCjA9wKMYKMDMdGU+HDFkXaE
9B61jz0ZCvmvRWUFOeF5d3hFZpm82BKziwUo0haKawQVA9CtkxCs4m1E5TpJaZJAqbNS20UliSjN
8Pf61vESeiTAHayrkTEoAz/4HNkdm8rTwSjkz1uXjMKUpoLy5/IsD6PubH33p+V1KD/tw8ocEjxe
ho5u8Phk0XIyooRyeWa/pWp9EomSOyBDq69O5Q+NRHeG8OKbyM6XjbHNgkAL/9/s7hDUVwIHXnzC
HFw1tHnX2PReFqEFASNFYi+pfMS5F9kCDzYQeEwW4YiIPk4nKrD9Y3DtyvFfndlqI2ykMRMrEDR2
ff0+ZIz+HSSULih2vvp6ArZPS1/ecSF8nUvO93eTNXjSGQi3NgSxmrCNKJPty9IIAB6uleVsiPas
B8rW2brbXeUBNQB1VNZXXqytzHUFNkvM6BckjoMN2HGEAhRpJWTuoLjXbM2Y3cAG8/hh717D0QYs
rUJYarNraV5+hFp7eTY9z9NqRLv4J6d0MFgpyKnccU6EFzgIztIfR0n9c0g/3AsHJrORsN3WRN0H
Zk40REfZP8fSvz2V37tZRxTz66mskHvERFNm5swGknLl1iQS8bAz0H1eFzgGr9CDuAAyvPhK78Wl
71oZy2Db6oA9xymawrF9sh1FhEL/rBJbQRliTEhgtlPsPHVEUZTEP5Y2pj2160FX4Nm1gSlBIOYU
9TQd6xGOh5DJA9BXKIzqejtM6/gXbnqVi69cujUxDRbtYIbJZOzp1l4OyS5fglzyrJGYw2l9XefQ
KxV/wgV0zloyZrDIxU0Cpavc5+QFhwheb9T2xvHOgbTaT7utRUofjykgKFgExXVA1CkbdEWVWnmi
eZM0SoR+EXjnUYmR2ETaBxCn7zbVf31iyWrCtG9M8Fq8Zp9b1ppGtXima85JtwcpAoMvpGNFMXfE
rl2AyUuopi9Ben0441pFNL0DmbvC0rmYM0qxoFobw6CdnECJgD2kdCIYJu5QEKjywnJYaYTftPV5
7KC+LqSTrsSJCvqtNMUDJ4PpeUxPssxOWQ6T8E618QTJLfRuXK+tjafwoa0wrFCS0PP0w8+2yeT2
5hdOwgCNs9Z9cv5G0q4aZxabTGvrMn7fSRZZch2jJS8TKrF8gc2JR5/FZVu8XpvTTnOd1Qu2FHW2
ZTNwgYbZBgehUfgPLWm4Z3cF0ObCc+cD+YQlM3HR/I/2kYYzBTZKMbrDuIyMjEMoLpA7MnYl8YaF
V5lxuf19P0AzFYzXu/rCy3HA1Np/CTaRlmZ5ohhiYBm2uh/irwZFhJfy5n7MCOX29kWYqfEg4V9s
kKxfkpROeN7eqX/u3bClGQdaK1NmJUaDPuzOayKOtjgjWaIEbtXLDhFNZeo1niMriSP6Wf6bmGCT
l94XD5NPXEber0jjU6/Sas8iPjkuryHGSSbpUmB34ZHjE6co+gYzQxrWmyr17iAu+vcKeqjsPJm/
C9g5C9kxLWZLq/R0rd3hu5cbFl49gI91dBCILtkanuMfzyFm3fFdqhwtFfoOUO4C9JnILPnTM14/
qcNYKbGcRfZf3aUgSqWumFIshhT55yxozpWpzqzer+2M2JABhd41Nt4zLS9rk+iAiZb+sjF6UOCc
+AH4B8tBwarTcgSvGg7V5eyRaNI00iJjW9tNNFHP2T6azHcFxiFF6CaDnktiDmZcrjFAVhnVVDt5
uasUm4dkz8fcKVtXxlFc2zYK3s/yPP2iINHTAoZ/fonZnx6zUyBubq0mO0vcQ+6UTONzYX43ZlxT
z4n3t3e3urLpULeJVto2USP1HMqsQXRzGk0csnkOedXgX/9Klcgt7vwo6oqQqL7eAfjncpB9WIpG
JkzJif2Y1pzsJGLV7IGStvKTi56CWu8ziobf0As8qJ3ZMDLI7JOtiYzY2K48yCS4KOmNdvjA6+Dc
Q7JZUarXCyyaV1L52v3ay5p9pciQeLgIb4xBkSYFZOm3lg/7VCcQuwWoVC7DHaI0/R1zucpC4qhF
eedOuk6yEMV8uyFcyecJuY3v5oZhvNgrh0AFPTLnXTv+D0yAJcpJN6qMfMblvD90TPPo0tCHeLzB
oHihOIWbiSl72DI7513m/7ixohnaFdL3YJ5iXxrWken11okaI/Vl6BXJl7xnHidfiBZEXHISsKz4
Xbabh3BtadXuLofuSUdSz1gvDHhwArwyeyYZzj2xeerfFz7cV2SHBdB5L9V/GLdG9GWc17ENqnyC
NUAHI1lHW+a//UAnVEnR81+Es3J/nR7Vvzj4d1j6eaiKD0MDG2D+QjQpxnwOUFSRSm/G6zLCX4L6
vE+4tfsSgZc/PVvbhR/HiUW7t80Gpnlh5Scdwqp2/5GXm73qr1fl0XQ45oAx6MadVZyWCPDCuhCb
jTG1WEjzAYu4GvXcwdipUUCpGEUHqkucZg3kDlVxXycmnSej/JV1hfmQSgN2ruLmhXyPje6c7OEr
wRtCCrgwpG5LxAFTEEfGz18jfIXEsS49QrV5nHUg+HB02og0yeoTXlCrGJfc3k09hY8v7lI1X41Q
eZHFZUqW5sewm2bFzfrjrLv+QE1h7D6Fx7MPf+N4yzMqTNYaLELDq6gWhe8gAv9xAanUSJAe9fFq
0Rq+mI0ASL5YWZQzgUj6MsifX9N4/WRCAecHh+QHanlOQBow64W7BBRTeuphln+iR38GXvlGCeIk
i8JXFTffMHwXp+4hSL3sAGiHrEezO22GvCCXMcUesPdIC07w6/15CiheFCKA8mUeD8iwwsZ0BbfI
RkL1fA2ossjM4jDRTeZLwGNwdgTERtn1X03QCzVlCmTAApajDkmcxxx0wrZ+OaZWxRI8glQXuSxq
hQZFXdwCrByBTROjHnUC7jAzdnKEuMrxptwDnPtItr7Aet4RAU1Qe7O2V7qUfsf+y46rEabH1hQZ
R7e1D9Rs0pPfc/5tPnVxhH8Yo74o71ps0+JlAlKjW4zMhXd3dPv6q0YVcaqL9nft2iL1Pq8yxE8u
Fcj8lBgYZ5AfE7OhvQ6Ha5FT608DPD/1SWXB6GnFFBUc/AMBu8fJotmWSZe3yjaQT9dgemeUOkuX
PIgItiUPyfRgLYSAAY9TbKjhzUf2o2IZluPUKRn+Mm+AEAx7dlCt5ZHCfSy8olW508AZXZPwWOI9
Uu6/CEBudQPXy8gihv8dh89nVYge/iCQqbeDzXN9yMcTMUV8lfycSC6VSxkbdFkPM5VTrY21hg9+
O2kBYWpDUCPmsvt+K8pwd/pd2eWD/kDZVsIbiepJn+y5VPp28ZThpMDYthhmyU+AWFw08JDpvs6i
gpXvQ0FR5/tP1MYZUu+KBjGbjtAuJj83c1GAeL+tj74fu8T/C84ptb0kn7H7McPw5zu4GVu/j2xI
z/qOZPqMtsRfssZ0m26HFNJYIiUFxhf2i4XcqaldTHuZOBmzZ6s1p6AuZ4gtJaIxSihJWW6nnnNx
cxQebYJmghHckgf6f+h3gX1JnpOpgL7prcFn3uH+Q9PC7Vi4qnSSo4zDtcaoE7F6AdvbQzipYFCX
OenxlXLwN7xaZFjLOvccNR3y3UjFgv3vyx0BmaRSjwbVOH2q4SMeK0Gcj8WEEJWephx0qxvNk7W6
HI1ihnSBLfVkxdsJahhcyaNM//wgtKh7jcaWQMqc/RWLBKYsMPfnKLQu4WF5rsBmwdiXHurtlqFp
6qMeJIRdeyukmH9Sr+hyWLzB+X2GgYZ6gH6C0qjCxtNEJCd1/gKTdQ4z0pSodeuVJnfhPcM4+wRY
rcpQskUvuXaTB+kjE2WIgu/TsAkWOCmtVSyVNA5V4cgABbXIl4YsOUOrrSUl0gSHkx+qXI1j828W
dyJsETqVlxI0ugfQbFitavMpoLaX51SWFaSJA2ElQ1jTx4KYYRvWcY50pPBWm7UGAf1u6R5h/Vn/
Yf8eo7gRBpFCixV3danSbeHHmLQWLYUYB2xOeV2+vUbNzW7Qsg4YQYi9QIeqhMPffVoFe6rHTO0W
/0+Zzq2aXL+7lgKyZSFY6iwM1zdwEJrhnNTPGZiIlAozRJiI66vNwLiesLeM0Z9sV7AXS6YKbzkk
/czupL55vj1PDU2h/uY3q3+CBAhGyDgh2arQAhAvxpDmR70binUnvztZNDu4JFkt42GgkdwYmFmj
tcrP/IyA01D3cPIezYMPrCHcmXwfNUs26ItOu4uhsiuLykJHPtTwfELbxD7BNXv5+5LmBRZ0jnTp
x2++yxoYO5WYmbuzqymTfk1MrQengAWYkPlb6wV9Lx33aF974aq7hZMzaiFqk+UwVut4bOfDrpso
i8r+rkIvgs9vEESbgAvrPbZV76ZNheT+XlXzOMmn3qUd3T8EE9MjS86Kr/6v4kx/7h3wJ/drREa6
IhQc+jg8AIj1HmOGA+XxKhHyua0SSEbzxsuHf/NOubKXg5RFlcvl4LrTd6NgD3+DL1vmVWvt9cVy
PLSYt6VGXrLTI+R8GT96DjEMBzbFQXtVYeIHg8fg1hyTZ/FpzVsES0/7PmIjMA0p2om5DmnHhVYL
YDcbznCSpzPetJ2La69xl6wpmHloolF3Y4qE/q1zA6nRse+Aq3ai7RZTlIDbwaWlPfSIpCMdnn7p
A1Mr/aPi1dSCPyZe+QvQK2ufFdASMJh90tabr+kX1TwV37o7yA7KcyCJUHbY2TGEUcsbCi/GPVG9
lNwvWRoe4p9LvVZ3RXdEbD1PoxcMjfxIFvwHx1ueekTHTm8qd95ai8jWp9dLpGR1LLpzDZvVt2Mc
/MNZGz8Mc1i+xJzdmkf/7EZzyjBOR7ns11kEWbM1wVB00On9V7buo1C5nzZP93FeffEkBPbszVkB
Be9Yqgm9YoF94sZLKipL1h+Pmxz4FfiFhdoycPcvoB8uWyIMZve8/HbHR0grXrtcMslVau9VL8kx
4DUHX0VGh7UTH/9ALVXq/AF2JVXUOxsQMxXbyODA3QONrQ31/vEpVXIGfMaZVtz+TMwF89Rkm84S
XawAONG7WpK/uN2GY6VmGl6awaq8iBLAEiUVsgCE+kZKm6v6J59YcM/9P8F5h9P1SV5NTPO/QrvI
5hvMivr426RWjCsaLmxXrOkxCFK9kTNCEeq3CGlpwK41dkZDtLFqsEKaBDcfU4p4eV1ZxYyb4cKV
9ajIK4rFtleEdKej0cU8i2rig28BqGxFpLio6TV9+C99gxgQF3Bvg/4c5Bp3VrFcSVupFiWdZzUt
iMjGTrEeWJzUZWhQG8Xwo0qOcsGJM2VqVLM+F3gZsz9N2lG2Ptgz+GVXjMVufrBuLHPBJZPBRibC
JXU9l87dQ9eo3LN5IgBrmGicyCePxAWC3wvYVSvDY6H4RFReLGXMIdPCd7i50lvCiq/B+QDMnxQi
2u+GvSvTUFBW5Sf9sRzDW19P0RfqFn7SzZnIxhX8/xl+gMVgyeVh8ydCCr93260PHdKbwAsDbz7C
YQGDKIVP8o9cR10YQntQU3EXVIx9n5ikgQnPZIyQqJZd09Zu1eD6AD3ICMi6+fWF0dHAjh1myxgs
bQ0BTo/j2uk93nNP5yBImQwc3yh3t92d8XdesKKfrHEOCuR6jUe1lUcrOlao4Y96/IYlMUAmvIJ5
B4LoQ6iI1MU+NP5Ccy2VNgcaBAcBWqsWJ/X1cPxNWCokj2YG1FZoCsgKHQyspsY78JgpS/azgKEI
NdPg0EF/9d0/vq5I+qCROGpmuXHHtN51tToDOhf6P4w/EvIgtnaub41e7/lyEhn3hM9X+jpQATbf
XshonKhhylkeST1KGNSqDXJ6WJlnNaqR+dvM6eBW0eAzR+dvpakIUfy/Vrj2DHkwgMEqlnw3uQCB
UVkXULDa4VsQHoVFk6kiucDTMmfJeM1MLpD64SxEGFjmb8+nJYIN9ASGo069LFcqgTv0v7xd/Asr
Q9go9HvItT9E1+sh2AkjMx/twTRTHUKryNsprjt2AzePZxwhNvm3EYWZyB6csclg/uk4MB9z05WJ
q/eKA5OIIxMud/qxCBPMKjakinBQCPMXBVnqgndWXrjD4Pz+22fmHm2QLZG2Rk8R40G7xE0/LnEv
nwxM2vyxqKFbIwB/HDKKH/99oPd8CzLQpM1TXqpA7/0Lwv3odJmSTrfbLZ9OxIZV9+RnOC4SzNBv
K15HO1J/ldIcG/UHVKH18+0pTz+oBpJS0PKYBT63U8zwKrruOHL6jtVoW2LBFAomZNZJeI7a7rz6
jFpJZ72p3Xj40+JFtDc5WMBtrC6CTgBGdqb6oX4kFbctvRg5acOhMa8PhsyN41cfHss7uYoDPW1h
6m4aZm0U4rqHMxWru+Htm0T565DY62sTHnFsbvdJIni5nIkLtty4NeamLUw9u05nTo29WhrsnI1w
g7gCBYoUlG+BMcRGDOFyF1XGeO83Wx09b9HJ103LIkyQ5GQh77IosqXGzpeoGsFKb454Rni/HWtz
uXmcZSzctaTS01xkWNAlg0Et65kyvEJ63yAVboEU3UMVQPz4bcGr9MjCcNmhXeVaxqUszZ3NAKdT
F24RpKUzosbe8Ld5zG4Gv/fGjZYKQhOlMRFZIoNvIqBvE0JNQWuaKRSv0g770Skqzm0NERtJQw43
87rWNtJpKjinXH25oagqO+YXw9TUHphl2RyEEcrYACJ82pyf5TnH4jWm85uNlnQZ2GmY4leB2IAJ
t/sguhkwZ/Ophz80bdmhGOonB80/Gb5ZQtf0iq3+w/DuuPABzs1/WEo/B/T1FjSq5927J7jrdlwv
TRHsNVw5/DqwAbY6qmn92O3x2qZwqgNwHZrOyh0eTuoddclzDjlRgeWBrt3XPlrrv55UVOue97+y
C/aLq1jyofoErVss4BvR1ygV8MLlaRIod7v7PRVYvnRiuUPvW4XOLm9aoQn7SlDAerMr5UFNFpaK
kcvuqogk0krC17YVjCuCp6dNqqGq18iAEdoCGaQOwy/o8jxzUrvB1cKtpVP5hgiHu6afl3PED/5p
jeVksCNmnUKCiLHv6DslqHF2R/1yJskG2cSJHjKNXPvFITB1AX51F1glzSuq07Etlyexjj3pWdSI
EkX1GtxGnDmmULchb9BlJ2WdQJMmsaquYkCOopbUumSeg4nZDFakyf/JG7F58uuwp5pGeWf5+Y6Q
TN/OC/lNyt2k3NiyfulbFP0uGCJjJg5B+srC8B0wopXkn7/DzNN+ABvOjJQEnxPT4O4/q7+E2urk
8Yss9jwpERu10leGwqEJ164AjhcLn6RWzBqS0Onx7IYi8OzNtuliTT1WoqZDF8npp62wy6lod2g3
xjTY0bf9VVKQVM1d31Cs+X2rOfT+qGOJvWYSuBx1SMwcvKGSDix0bSxmSfmQtUCWzffB1SAPbvU9
3gNCWU5iN74wc1Ho1dxs9Ggcoc5TpPadK+RPByXaNbCKUBKknMShZC27lOsou/kIJDF0LF1Q/UVf
zEthixz9BiVP07WRwR/j0Wh5hDaDbejCbbTHHaAJ2wYyAyIg1zzhbUZny64QFOglfQnB64XyNQoH
xOKTS5pLpuypYg2iCVP3ZRE2i6SzNptc/BQdQbHVsokqD89dyasBpCWtOIx6q7ROBLsrzp03Lwnr
1Ivld1tBDUkJKyi0Ocv5ET0UC+sM0nqSh2Fl/eHEQu5q/eLzb+ydNK8qBjh8fPLZKvAiD2hxj5bi
4mMQfeSn2vwDNqhnyfs4GRkOn2qppyBD7ixqv6WgFDK7KsaB4JWVVM9KdA0XNiQzSEZTBG4ypK0P
AY3U6PJkf1m+vx5qXJA4x2+vySzLkbUnD9xFpW7ysik43xVDcgwD/XoJqeAIKFU+cnqprl+lWxZL
34LhEF2OMGuEqKBR1QezYaCoU5drF/CbIbLFaz0atnCFzFb6pnBhZ891luYaFhzjkoBtdlbF4W2E
Mz2JmlHq18YHz+IJqvRWe7ABKNNeSM/ObnMmfr3yU/XCe5achbJK5Nk8KI3DofctPO2RmZsOWy65
4tCkK5Hp7lzHRFAnZO3OUJRTNAhrn9916y/PNZalFQZJtMq4FEsBWxtZGtzYEBghV4QeH4ApSZbQ
pL+qj9s7nSIOCz9Jpur/EYXNhnn+qF/jAsneTaKaAHIxtrpMV2Ynr8x+RsG+zCS2nsfSQKorBFkK
KtUUzD10tODXz3S8vnn7RK9l6kyoJCOA/wRKwBZ5AoSmBvdm1ocibrQiYtrIzHdZ0Pu5yi5+BEoN
+2DN7e83KhYtnTHMA3psb9nI+M0qnthC9qHFkNuZPLkMhRYAJWsUBgtreT43NLNcpeqR/uK+Je8c
hxO+3/pwrJIl/HmpFKXIn/ngX52K90tC1vMzxBJdl3ZFknkb2VDkrG2NAuSD1L/k2mp+S7cOLD30
+a+JSTSymRIoZpj1TBcAw7ahnDuA9TzXKt/GZTwFMY7NtnV8PPKWtrCyCykvF8eoO1zyley3cFBn
tOlzOI4VeN6/AqdHFFaghKDG7t+7+iOH6YONh612EAqzvAZu2QdGhFvdyx7XqM16aGXxkklIEI/n
Tb4SLBlPu9pEQT0h2acqOh3PXq7/d9wwQAuj9i3J5Tn8EHeaqqTNXm2r1CguyqkvJToDCOUMoVVK
Eg3BXFeHAWTPz3k6oFtKTI0th4ldq1yGdILtayr5nraEi6vsYadUmp1qjpvFiWTp61PHE2nhUvFR
APQdsiO/33pmLXGnHJExxC35ZhQPOM5ITrSmmYMSsFyi0tTAXWYqaLmAMDx61wUiJ8HSoFhvJlBK
8CYRe1XCoMaBP9VTtStv6bwHF18SGZiiKajGvBEAVqvGvyjwoQpDyXBg8g5L4HRaZQ7rKlklcHOk
/pCH41UYdvzAwtxUUsrCacupARo6FjBgKdCg4OCfOLny140S0CQxAcP87SMmwm1vAWH0L/KrI6tz
mD8o6YSk9AoDknOBq8vPRyvqCaDkJZsKSvn/e5i2WjpOYP1NKusbjBwQshl6zb5gtZBLoTAEhb4g
gQw+YPYm9Tfv2uufvIPf6xluXvTtz1Akp52gDwD9XT2VIn7hpPEeP4W4kB7EByO1o4cEribbUSRw
TVweml3aKt5lq6NTuAvO7hkSOwSObtLKdLiLQ8uwvmGrjmsf2VQukJ2+va5GpYGBVr4OPQTpVsKC
ZSE2qmonhP1qpWPLMR7B7OIyBn3iHbJ+Hkr093EGcU9jx2MDNM9wxexSZcYTTp2dGvMEzOx6O/2i
VUb3ohhtwZWSiBRUN0JejWGIGtCvuLS/sSf4anjnl53U/HjGGiIZC9/Pd9B2Du5QtzFCFa0cQ4vc
xZ7o2AIkO2eAJf/wV7jRAKJwBhy8oECR9gheo+h4rLEWbumyFWWwas0lImaJ2SuTdYHIv7syN63O
PMvF5xWsPkWYnBlrifD4TdVtApmBJhr1fx5q0I7meJ5sq/2dAPEN90J8FMdVxxsveHAncki/5D3Z
6y8O5Yxzxt2kb1lmyfRSRA4XVe14+uWgcQcbzuuuRYyY/jcYsVghVY4uGpCYeZrCQt1UAQDdYaLG
oruw3ndoQwZ/2A4vF4bfmScEUbdYiH7v8FUARi39C2PHuq7eq6UmTjhuFWzXbxWuxR7KkDMTMsXv
2GHpGg1bU5z8MLv/8eQvw5TVfbaPnfrvCmA7BrLQMiAGxaR502OmnaXgFq7wLCmry96nH7iHSpcc
BO/Lae1y/lpGADTJW6dav44MnBuWr1K86JKm7x+n2J1FStTe2x7ilR1UMF5fTXANET9HDpHMXWTO
1MkSDSeuwz2pzPbGJ5q9gUkfrCnMV6cgljzaO0RXYCMKhrn2jFXmupbWnRaakH+ekJS1B4BtnQvU
lcq0bHq6JI6nD8gRhfunevRgeHku3wWPgyp08mya2zWDbWdnZjWBcd5z2WWgJ//c10UT11dRtYGI
8YLDz4R4Olit4OBShsBwQF9yg0nWe8Scjmf1CaRgTrA9V3EeqHvIim2scea5sYFBw0FOF8qQt4l/
T9I8PJwDVEc4Ixde9/LpSm5pHhsHL6DbsUeAz591HDOKsS+7Hp07Hk5TwNpVRAMcgcmV3+5EUTjd
1Hywkw0D0SevuOJLop/Cu6kYFTCMSj0XV1RQZvo7nxb8KOKoo9qiA4M2O4UVRlFD9R74fgC5zeB+
vv7t0eXXt57kb2K6jLxYxe3EDTD20o2W16vTblxObFfOYEHIsXJgWRC7eGy8Kisv+HHv8G0V/mpI
U4tATCsu0VrVwLG3Ibjny9bs15TtsXfDIhTnmraCkPVYsdw0GTmZ0mf4xHF//Q300/2H1yKZWhny
azan9A663XcCSpZOFdG9cRHKkaqG3hX6BJH6y718KhE/ZJmQ7e3DX2YSUgwkWtP7xL5lZWzv3Xfn
/KjsEN5uDo1UwdB7RFS52ezfgvibI3d8U4zT4gJtmf5+hWzh8ahaZRyZiLd9raQc69EanyuxilRl
pEnGa3KdOWO5UosveiP859Hpxr2Ui6EXiZTQJ69Fbb1x8o+U3iF5YSc/7mLVLYS07gBDVkK+YY7x
JaBaOViGaNuXwd9kWH0KDYfYCWegUCCWX+cEe/aMhauXZe87s+0V6a+DSlawBbhTa8SaIvLiEafw
dlDM+TlkKL+stDIKuYwA4NL1pfQ5SGqOpfEY9+tFtiaAhITfneXzCf3VNLiCgsRQyjzlPr0c11w2
b/q+n6N96dor4C0ANtJgMztwStqmFZaAXCeJTRX3oSt0EKiaLzJb3UDJL2Y1IhON7bivZkwNOYnY
+krcRRNhPDnrSQBsl9iv/FqJECQ7NO4D+QuTpAFWWjaCFiJxQKh58wilBJn49M1UruR7NG/8QVIC
/jPZM/C8YiVvyCFoA2l72robOZix/g/TRLUcWvrPc6NhOmtt1TRcHFzEgu1GUYWVGm+DHcSyCtlS
Mif4ozWOibN5YWGJ84yMaeGhuPLIjypHgt3yi+gfFe4B9DbcsZY8KpmNuXKTpnk4WgFek3g0r8Ib
pKWalSd1aelYEDvx3JStlAI0bW2npq07J/ZbPgPLsW+kWMMaGeMCSh1v9FI+jG8y+37HSgkTv9fZ
aS0Q90opWmE8alepuJmlN58yt/DH3i2YFyTdtPhkciEdO2Kp3RUa8zGdBQMBGoK3U5N7yKOGIHHl
jD7kV/33hv1I/KAUGN7sN1WBM6yn2xM7Q/SzwmLTWGL0Va74vmzPtA21cjCwmblzsjScP/oJ26wX
m6Em9Y1UB0AAUAjmLG6HQ8lyE3AM5GlKrp4uRdfBfcgvOnEA1BICOpi45iozASJWOm3J4YagohAi
td0524BGm9lFZkZUnAeeQjt8AlOO7ltB+E22nbYeDPo2cXtaxmnvR7wnRrJ0BZmlnOAvsXlOWSr0
l5RVJaDDFVEaMHf1AKS59LIXg2LlJ9nrXCXYittPDRZfFtiM6gOw5bMDirlGpWwAyInvGOUlGEFp
atWvRHqRnU3Vk0zWzrFBXmPYFdQcQJuq5wCyjCa0Up0DzU+aP0VGQGQsWxZRSHoF4P4t8jg6jlVC
THE4jL5CxyQmcfTRaNMnoWVuJCSHorXoWnPxPc60mYE/bv5NaMoBV+0/uzb/68FaEa1QYMlqRc9x
0h/Hnh9TgLJjXgbtbwKicy9rxEWqy0KMngPsVyh6+3YqUMCfrHfjwpPfx22jjnewujAkTdvS6NSs
lr63RrHZPtWQZ+mWc0biptq0ieBJLXT6JvmBq1AOjVAnEBaaEX9fsDm5esCmznBYwvWM7mChmcxD
3ZxUN0TjNgKuzHEZ/fBRgtGSbEK972GQBGriFSBEKp1eBMBl4OH3AoHgkoN/PdYrtIsslJmuYh+N
oRisA00BHiaPXSJGs0piV1q0uFEouiFJaqkeno6/bA0miTtjbv+dBGPs8gwV/AJ1kcKWt8dPFngF
iCcKrZcnKp2qsKS8w9uFfzaZWSogmLufxAf15h8F0tNwfCqeReXsTBgmsgSlq+Y+5eOr1Npck6fW
YczrBZm0iHgXVx7KxOj7js0EjyEm7ejEh9Hq9Zqoafj4vzf+d6Ko21bBl3C8mfc7XIFZjo++dwIw
vQCoRX/T7YkhaYFTA5x3PQCxCKzaDEFkIu8MgduzhgWsERnoTuISxvx/aZkUpFGoDTJofgMgmzad
tS2M0XG8ggEATOTkp2JGnX3AUODglE4SAKOohZndInW602eBIEu6Pdm2+YV6YQ/9ScXqx1jO7XVE
PSiqKK7NUrgwB0BCmo4hFsJLzrozjQc67Bk3/T/So/H9/8llLHt1KW/DpTGWELA0WJ2RnFRYv+qO
O3rsnxyZNfLhJoO5HqRjUcSCvV1VzF/kcUiCmbsxsBMMVzuORlh3iAgWxYSKi3xpPIPcrs7gKdqO
RbaIvDa8FgGbRiLWp2x4ZfQFzYK6xKNXfsRSK0+2JKgK+9dM4u7Cf7RKBCxXafqdEQKlp7ouuUw5
dMTXqqFwfGYSUM33+C0WOtuTrRbs+vgIN3+n42IZemEGenCFjEtXxRka5hejTCJwgBUGNHRZuffx
FaSJHKRdK1RuomiKIqxrNL/aij5Awt/uzQY5iZBMeHg++6FJNjAadJI7tXL3AqDOqJsbbv5dw4bk
D2eWd69j624jPFkmtmXRcC1MmCEFnizCXYaP5e1T4vI8waNLuvACUMKRTNn0ZtAVbUf430bT0gTP
t3IPBAocYXMUP/QYFJffjYUKShANjkGRcazH+1IyJRqGbOy+Nw0Wbha1qarvfB2SGW8jqGS703ue
eqgpvZ0qzGEvrEhD29xWo988No2ieqUz4vSovrQdmS11ey1LK7TLfSr0VSteSsN1MkuVxGyMhjV8
+UN1k/xQ3zWqT6pQTgxeCJWYDidC3MhxZCUonIo3H0fEbN5rtURuyJzSQ12WlOSqH0gGMpQ5DKDU
LjLS9D4zgklF6Ly9rxIHkrOcOzKDEBUwPsTZ0GufdW34TbJ/Iwh1TaRy3vL4UDUfH7D9Ks/uOO6F
CeS+qDQwPs//62D+YhHUZOhmHfGyNl2+caDtntd60pgwdycUjbt4hgzNLZRPrMU3+ObFGSt3Z490
sXFrh48FDxGBcB/nJwxShT1egCMR19rlfhPQQwoio+LVTC0IdkanK8NbB39ht8haGQlZzARw+G9K
S03h+tlZZmId8fD7sUF+tBGcrkp6Wro9lZ7eirrUW2wHpk00yHBUGKt44I7FPOKnuzOEKdNKh+nb
plYjnFA43Kol4SVtYj62l4yWC+75G66NYCulPMkK33uoNgHviFuE0o4mRG4AFkw5nhzoaqJ1Q0Dr
9IboMOfJ9Jp0wv45s/rbk2SYDhsYa79Lc/wrgiGuFE5zjyMoS2Dhz2TrHV5d5Tlx6+zj8C1jwWZk
NSvhSV0/qssn29eRIA0K+T62+TnFaDhiRk8B++EPu8pcXg+7xHWNTrVDcDI6cQQjzSOzNf/DJ6GV
21jqGwRETAQ0wCBpsq0Z8pz5Zx3QGKSW+uKlz8N0mG13KIsG8Cr9ND7DBjGxoB8Xji+kT04Gk8Kx
QE9lHGe7rNApp5gmdNoifMThu7cbqDAhiadZouCX2gS/s5VgpY4f3ax3aY0IMtlxD2JlLvTN+ImV
nljllDfR1AQpBoG3+VjVWJqNBcPO5j5I+lk7vKFH6EvcFrrwkuRou0yDVJkUbtND8k4kLXmpImul
bFXOKUiWeFWhA+idVGzofL0PfWS14VYi+7mVzouIH8TJxv12m/D9c+MrysdnW8XH6eNING1fmvaj
gztOPiOY8QevvIt6zMNzg76SXimIVgqwZBEp7B6zndiyUS6KL0v0kKujHoJiBhbxk33fNbD7H3/o
aQO7lgcxuSqMOmXHqeR6EXegd6t82sUSWqI4BnX7G6py7sSgZyhD16TFShUDNVogtxwRTgbtP65w
bJHMgIkZ5Ix4qGvkkWZWM8G9yoHkRBSDqmNhl3lrPTYx5lp2eZM+lC/QtOMgUaAsSbBhSKDfhdDC
hHotDP3HRqsGTLZLAgrGriYsigIcjxopBeNcLL9ge/YEoMB12n3sSTp+4Eedez6Bm9x4IYGD/nkc
fFB/yW0xMDKJtsoW4hjZAE8X/9CnWwDP1ALu4bt+E+tdx4LsSMh3lFdbieGhJ3a1gXHuhKV7o+sX
5WVqLAllpEfi1U77iXDHcUSwIC1sjDLRtP+4G/9OZDGmO0EIPt0hBXomkb2ofrPMMrFmKQjglrCF
J/s2QEl7GLOx0YqI5sWZZF+/5hstag7E+UR5SLDcoQjbmd2k/oep71vmDAaEh214+Tsi0k1HizGb
QzRFi5Rk+njTHMxVTmOKK9yr712oxqm6RYfSNXD/gIEnildCeflQkn1/4JUoAK8F3NbfxEy1fdNp
/mgENnt6D/TZBG5xAwHhfgkoBXK7/BHph4whSJRe3RkoBte7YlN9mUoVddxOW1sZeZI5eV24r6Uz
F9wIUEvf47awtBPXtH1epx9wQepXSPPTC27A6mTH1i/Rggs62cWdHQDa1LhtjCelftowAa8ecN/r
ZXZz8ZCh21n/K2WuEklyxapwAvf+NADqMqmtohnNTFueELklpQ6mfeMS0jkJM9D5fZfnipdOpN+y
BdYsSrLRr92eGrnYo/umadd6rkY8NnipkkRmg0cKvgScMzQbE39/Rb7Ily0HrrdlogctxfHVRwQ2
n5+Rezj31sE2yAYqo+80v5vRDc9eOGoOAPkD+ClnG5Uq9OcfNnEOl4D25Gu0s0b83Ep+N77+WQpF
S0IqPqUg1MAO/UPUtuPwjPpFQtSHB0NYSmINO3cU4nKbdTxAZPqudxhXtPJyavZHhqFCfZMVPdvK
SWgZ0pYndoi0cj2pfcTGfsUXK9g+qRetV85w5rJOiAVta7GW+6lyizHHI6D3nO5Lx5dpxOaWtt36
t1yGJeSw6dChPaf7nkWVRildC47sO6/5W8vjgYcjJbAycy6ucB/rmK0A+OiBBuWw58ZJSW34gGd1
zAW/rOLs1bWEuz/la51QaQPOvQgXaYsLYVflQx0oyfHfujz1VgQ/eVEXLktH1c36miGFhhaRsujA
X9sCXi2Hno02FSZFMVHNz2FX9wrRqkBcGQsSSUNzd6/ZrhjyTcDRZwvWbKsWjrzqvJBAcunKIYzf
7eGtpDSmM2dnFzRCg6ggSYy/Gm7zJCYdyB/pVGhvFPKfpAS4T4hqHQWeoRVDzpPIhI7zCtCVoYI1
73zy20Sv6Ci2fQ0voqjO4TDp9DwPSclmqnaikZDlcQ6JP2/3vnrdc/evxrbSSyl5r8e/A7xPwNNl
C42ezXsg2i9X1ikssKu/fWjyAIw0U6jQSNfS6Blt013YDhT5OAy6WQXXNtD/Njs874PmiG2vLrjH
6gJLdk3Eqt3dOZc6a9IKCQyp34sJuGAI4jl28cT70eG7NAulc8qqzgccxNNUP3Yehe+7NzOcmMJi
d9EzkjADHfjAd85xgNH1roH1qaO0seVoE+W22IRuP/RiJz3JNEZQwfqdbAL1ooY9b3Yc1xo82aHv
4UopCeiBJuBjSDBqEXJWXh11q2fZoS1Iah4QBUNSigAtJoFFBFEEEm4gM1zOGI/tHeF3J2b9UU/5
6d8CnXblSSzXDMAVtygx4zx/8Tk4KX8boqIRYDj/omuOToivxAZLy/FaxdMWJUsuhOTPfvAPQLqx
jerqvdQ3kShrfNFZflqoW15CgP9pdJRAh0PeorvjYsX6A0vzELTN4VMPugcWGMtGeiJzTQNXsMN5
4ylnpopJhjKgcZ0a8qge/nVtOzCwZbH8W8GLrrA34JSu9gRYfTXqS+lBGUqaPf5SuZwPzC4qA7E4
ex1xe8/qg5I5+Aqvl5VZi0GPWwnYWB41dtbgXPvN4qy4Vdvg6+RQBuswNa+N34oFZukuqTWSZwbT
a4vGniydRh2BcDOnX52954MoWZH7OKc1FrR10ftvbn9FT0XTMBWPzkEstNs9MVOYMT6oelovzn5L
KrRtPp8/TgAGIg8KdRO1IEFTkIQYS+33uC0n8GhId0ERmNkS8/da7Pj6rCBbDNeJeIDygxEKN/sc
45eHnu0RgnOythaL5IYRJFPzcoT7ycpenlHk053xBgjv9tvTHS74Qn+AW1cp5OCSCdEEfPF/sN3a
I/LcBir037rBBIt4oY2XmHeM8J81HEeAY1U8Mq9soYhFOIaU7yhOeNH+/VKBOZ9t6PtsxrN3KjSD
O+zgpy33HDZTOQrYWvPr5WBzxSJ2o4UUpPun0eJ1cdvni5gWuSjTylyHYyA0mEZQ0HNI0Ge8YWdY
VPtjTVlkXMj87PK7r+3k2i0h/pq7Qh7bzaipJiHsTvgcvnZ+hsdZJxpniXQWSqcJ2xkopXavZiIm
+7FPMAzIQkyBmoiMeIXAJ1cQiRss3Sw7AGwY72S7j+JjEmuyGyw92tK8itX4M2xADPbpV92pC8cW
s81/rWWgM1b3VL0iyw4hyrys3NRvWdrYZHNELxUna1C3bDZsrf+3G7Mq+HpXFVOp/DmtYg7tFcIt
7r3zjGbVbfcDRPP8ODK0goMI8ibRi77SVlFOnYJzfBOErVp/mlTvOg6R8s/SG5BoXQpOnHJION4R
zjmZFPhCECOGDURsNDLIG4vXvJIybb5Cf4i//1zRd7kNnWo4+AaOn7Zsg6DizsxCRTibXj2ecR1s
EkFAU1aWmmKPCqN1Xz6dBfd0MEkF5JpwzwipgcU+SJFrSnDOkzRdE+4+tMVml8mRYX0IKAaFbtGt
DmJCVazYmyYo8KZ89eoLVkrvccpHIFcNuDYLS/9AA6NebCnjgk5Ts+5Vl7IlqFJmhLwChgBNkhG9
EZakFPJ5KpUaP4EPw0rktNnu74QHXVOc35VGoxDdfDgajklfObGqH78q6io2Q1bL89Qgj79ALL0d
4XXjwuweaIDbcXuDRZ2JvX7LPj19wA9NCLvNF15lZ7Z4rVkRQEMGQfscgSkIaYYLKVgZTxvGZiMb
jvaB4RbrX2aqG+U7LGC8ar6cQM4yEUSnzQ04PyoPGj5kBDZtuy2Fk37GPowUyNpn5oKGA3H3M6do
/yFrHn1JqMj2iOdNnndZOsWaxxEONri+EUc8vAQiuzX8RjEFVKUHgZyPWO80mYiuBzhvndET4TdL
cITLTOfuwnhkIaBOHyDJnuHFb49w965wBmOuiacu6cAQ+kO348blT0JCFdBTLdUlm+tJ4I0s9PTA
k57Db3d5Z208Mb1sIt6yj4393sb0CulWhVtVvQOSiVr83zbLRdSVMFCJncaJDjsC4sUFHq5qfC2r
1krd+ZgqTDohxGxFBcYnoPdQjsABE+PBrOMvaxy9xguXqrNtMeBhms5w2k92/L9PHbd1uBuk3Cm5
gDLMD2jAEG+ZvNd9lK6pEYFR1lTrbpFDBMFVDMfJQq2Uo5HsqrmkYRIiwfvUi06oJLRAIsRsLWoa
4DYWxXFCkjjecao2LNAJec2PZxxzsE5tzSQw8k4y3U33jnTPzoeGUAXjncFnwT0KRvQLuenFfmdp
+ynsqGDu1KpJ3vpEqDxqxwifdjXkCyBOftT+rnh6VZNotbbHPiNYEQr2Sv8gEhBUeMvdZOVdZ5m3
d6sah6KeJC9QWlfhMSZwSXyRYkem3eE4CGFJM3U5NPNNAYZKtQ58GdB175UuqqOgdDL0XEo2i2XA
Aoe6aCJvKseJpHvr2foIpfPIyT+8GJ9/50x3ngImw9ZkycQHMxmkOx16j24MitY723kdZujLX92u
XPAht3JQ3n5RAxy0sD9vQmwufEe8FGrqyDpD5e6a7FF37XKK96F6FbBpM1VIJ3SK6Rgu7f9h7HJT
xuVYzrfCvN9z97MSZOfvgzgb9JxJLe7MHUOtkZ/Pkci9OCS5T5EeVnbdVJE4GsEP0Oyd35stZ6q1
wj9elfR5DdMXQrCZMWEydxTGtQIRwvdycfOwOcmz0i8E4Jsh86Zk7fHqsN1bvQ5Zb7au7jd0bulu
pGrySZRi6nlTP9pK1WCrAHsLI1Dt5UbqDL2TljRi6PExpa0CzvjRiLUYOlBsrnPVfLovCSHcdhVB
nOwWur8gQqYHgxqIPlTvz7X4GcxCdIkuPWxZpFOSTTghNT3Iz2BpdkwHe5cAjJKxeuKrPrOfPj4V
89QdsWEWskzfYWVViMEKyjJ/uRzdnO4Nas0SF6vNK+NQmy0WObtKj6pikm1xkZkfQzfWpn0JfU0V
3+m+PwcLkHguvQKdJ5v0xTqg+a1qaBUbb4Yr9u7dFAS6DixTHrSjbbrVMcU9ioFA5snKYIUo+XTr
7MyESwXkwYxLP355sbYzirG0vUwMjWGdZfJHMwUgbLml6kKAKLbNVp81NtNT5PolCDTFDIgeJq61
2zBSpFpH0AKGtEuSXT3xPnDJKQ2g6KzjTUcIBxh6XBr3hu4uRg34FXvmZ6QpsLl8X9bx50UYDevG
Wz+4hKurKLsfuc+0jxQKQc3hGFzfc7N00NncAMEjgGqJtAIkIi0hgsVfE8O1n2eSeUkXAYQ6NhKj
rDesOwLMXpjWWm/LSF2Gms4VyE2RNA2BqQO2jWYRuc8q/lHj59+YLprD0CHL4+90MbLjYTTySQXl
/NZrRxnr8dHAjZzsA44sgWWPCBLDwNN7JNUetzLGV8P/MdO+0m8V/tT0LD/4Gp3RfZqJKnz1P8/9
7ZhYcEKRbsHRLYEsa6sk6OPlEQGA9H+eKbENG63xToQPfBPAlxPAihdTpUuzLyWeSg4EF9N6AA0m
y4H2RlNr15QVJdwZWIR0vOher/N2s+3SrVSkX6Wye4jc74RFog4IsE5KG2VhTRdZuUbDbkW2hZPb
OsRSjcWSO+WJlxF/L1hqDCr5hIfsJwYw1d2l0hVLLDfi6qYv83gJpMO8zGQ7RrxShhvz3xe1DqMh
Ui5kVuigD9MYnUy/I05jT1tP+EcQE7TSPRllzktGVhPjIoastJZs6KKkots/qp2lZh9xJjY28SB5
0yUPLQxW7IAd7B33J+g4GbIAPAWEjl+A7D8yQsgjh5CsEC7bYtYuRx+BxJWnYAlPJ5IU94cB3z4Q
3gMvzlxbbiljg/6jUF3B8J/DH9N9UrLqhtofNfuSHUtt0dfEEmQOXe3MUxaCdtiU9qEnLJJ7ODKz
Ua4OOCTbIIY2nr7XbNUC5mCEJGVZLMSRBJSQAHTKfEiu5bxi5lWLFNRNdbqxXU4VhlcPcrIiB0zx
3soe+OzIyiHn948ZQdaSouE+zVJx9opJ7OMX3wN2uxrMkcyw8HJouOSlXGoQPvqMP3XfuHtzZLwr
RXKEAvr0sraW2Ns+J1ylxMiMJq02OGagOjkvHk3Snvylwfq0djJhuoXf3sKCw4LaaVn3v3EsxeJz
uLWazpr8bpUq2OkCBbw38FUfh7v8hktwzW8/FIESAaNULpDn4aegYI2YZAQ/7f3akLkwZI2cNR2q
T1EjjNMHvZGnKsEye9RlEfdlK77FRgtZpS6eRh/30wCxhdFd5tX/SwnZLL73DWTod74zZD3Rx3eq
mGRQN+hLF9CssEkNAPS/4LsgDhjaH/eTcm7oZbCpFWzm4mS+pYFvobob8eTeTYETO3LX3w0RZOQY
OXGFkVmMmw8DBX9ggQgyLu3G6kT0I7qe4dCg58GRuz+XXjcTUeeonvXEzyLqq0pmueZyX1kDqXrG
kE6Zj1AwO9DS8FrCFhfBy34wT5BOO4l4RycEJhwQ/1aw48R8yq8fm19Ba0QtPI3tw0Tw5XZzmacU
HIA7RP4+2p6cD1cMVl8FecdA02scPWqENtJPtjuq9yKpUlMKzLQ0rBM0wSiKtui4OelvEjziyyS7
P17S8gfjbSuDK5SAbhtNQVfbhUvP4Wp2GFUVjeFbSR4bUfh6i6rbmSzd6DoE98vIROYl44LfCckP
nq4OYjvR5F82P9tnnTiArvBGlnHlzLcb5K0IDXCfRaxItrY2o8RFCl0HfieGbQFAcTwAQkNQw03S
CzCG52sZOApr2Gmwz1qnvSVm7myFNddy15VMf8yFRe5P24sa7ursh3C3eAZs+Cri341Bwdc9Bl4l
ZF+SIxAh5GJ5etynk2ttMKoWojYmvyeM6AeFWpFVLTaKsjBuULOWddjKswAfXZjF2hAPhUymubQc
mJwFt4RDd6vQpnaZygsuQDRY1AE5cdvswokfG8jUMEx8o9+XxgL4ppzx3nq2uwPV3HJE4BXDBePv
YDMJbbCVy+Dp3G4piNfaKv4+1hJh648o7mQ+51cKufox57YWPiA4G8s2nYmSPHAqYFFc+JPH70LV
yBHPyHuQwmsqnqOSHSjDcytwbLbjwz6HMnh+bQssoMupIt/SGaaQxkh7CmIPpFKq3uTJjwt0cKBw
BYQUlIDysgQpirdJvFEeg6uYnznsySe893qRn4Z//bejg6KFNnztpRCLXuLtv8hQJirPSZBKHIlo
0s8gD0P/zUVP43TEg0g+W6ZYOBSNK8Z1vn0qglp+mtIn/iC9OQBOkPxgo6zXcrJzB5T67jXXC71D
Y+hnWbKj9qIOTZXK+g3HBUipkTsGNQ4QRYY9SLHaFWsQMN2kDpWJ0FiBbLiPDDUMP4QXUov2zv8Y
AaEWYvCDLRhPmbbs+JZAjziCir7RWGwT2GfSZkRKVcRazBa+Q4wuFxUVB171CZZk78SHutjvwJ0J
zMjA96+hnqS7nlqixtOt/+/7cGSqtoEeKRDnepRNO4E4JsclqAPUGZHTrALPIr0V8F2xPvD/EqiK
11JQKO5W30Z3ZooJJ37mTpRMRmWTaG0Sg3pTSgJm4cvvJzw/X69JldBvKKH5PlfqarCvH0DZrrx+
VixCaTwwKEy0ygRVP75GW1DdF6pzpVsnSxZ4wC4YV/0tXgY2QV5SXID00dnCsYZk30qWtY424R3g
rlDR4X5+8oGRyprZIky6gb4sldAup2sWeniCylVHNHVrEBpRqbGBLnYgunllrYzEWVtZHAJ+r12D
nZRftpT2DHB9GsI19cd3rTTkbqyRXyN8QN7t+w+ywBSCeZxKQS6qZwYLtMPRWxXSlHS3RvFUKuFu
yhDtBYsRNpqah6EQP8G0bdrEhbUYRHtMVuu7nN2I+9WmpiuTrEBxCYJRru90BkfZUYH7v2kLUwVI
3eIgQNGexEnBbrCR7O2dcLra76WR9i7BX6NqFLiiShsmbHxitr0lyqUYm1dflDZznUGD5oRJMCKl
LYplAnrmYJERw+jIOVXysjqVCS90L9NPwnzs3Sjo913iBQf6/RUs7hkHNLso4ZXOucENPg8WON7q
7NRIDq6KDunPvlES8oxnDlrkuF90bv8ODhgJRqgDMw0VgaT2zGx6LHVmOljfuOFaPVbKkDelDIRV
Re5yeRApCfrDyE839/x7UquwyDswb/1vMvCJbER6ue9kQ9sZWtwM/6OD5IjpO2Btfw864u8drxye
7O2MfnuWCE3svDsA/V6mnUyBawDmKhfigzsIkh7pi494jtIPMTO+TLyK695CEXAu8DVWeYYBhv1T
rSnoDn9GqnRWrcGp0woTN39AP4lGdlfzf1FpiDEQMgp2RGOmcT4zwQ0hEXzqwdJded7TrQeL0m6B
3V7fjEi2HB6OfHNKllWVfqqtq8xS7kNn3fq9MrP85zOjmWcVDD8T54fR7GUfSEJtlIXGiQdkd298
Swk0/HFWBeWUoDlB90SMBi6ZTJygtlQqWItT/wC0CW+EpCD+Ed6jVH1Xpp8izElFABusWKqI0wtW
ujU6JkQPW5nTQ4HODoyKsuFkCSH12bUdzscgiR+/ZAGglpUpeyIpG5wkJjqCindhMjDrnai7pEUc
Lw8iqwbsEhDpstw4SG9tDL99WhcZq3P8QY4Hnpkgh2zTGeNHjnKLCD11CMe4WCSQWWSQsyF4XfZH
/C8f+hCLCStHJmsm//MQJRK9FDlcz75e1IO0LdAzfcZcCvJxQwYEOpLQ4+kY9oxNFfoVKMUjSZVw
5VJDlcnF9dx8jc3OtNjreLe8D8pwMyRjm4w0+mfaILkz1zuVa4oyWbpu9AD/lJpzPjEulj01Hutu
iH+B5nPyYMXP9hkFX9Fn621j2A+nDPOZRvMCeOEWH79ScniwODN2FNoCCnFb/HyShU7lpNC5BitB
6Y0DUTVYyArAqc/oJfiRueq8i8BhhN25QnO9dOXw3LdaK02beBogJ2mUMF9++FSCl7ZsiQeXuy6j
SglYUbCYRYg21MdeC6g4sPs0Q2GUW5J6wOIOUGtZmh67lLsp2tOmZbHS6V5yDZZ77dHxmlTbWz5s
wIvdOFfFalqjQv4qDEqgGfe/tn4dVI8L+o3JS5necOKzLYOHSLZLzcaFXkxMkQqgoB8pnQbH9wAK
2Olo1OdBpdupd9X8RQWt388uveFA9t3CiWLMYU+w8szTSZYhlMLBhRGpc67pueV6fbXxCU81Zyem
zgCB6w9pdTYTMCLNg+psK2QT8kGWSAe4t/UVbGOw7UjKEoC1fdlJAAGiKtQurniwIPVDIViddcF/
Pn8kTLuPxBE1zycKS5zIbIjpCEY++zvotliEZt/Tgoe56kd6eOqx5rN0U8eNs33lOeW6vBcV/Hnp
v5nagiQEVlqQUSBuC3fioiSxvh9P2kHJSgGEP68uJPD1FN8m36xhDZATcc26omt76efRXFS42TfT
OaZDf6kxtmjNs7tPO/O741IVpg+JcATLx+UFAfxEspq2BBly+jlSm3NI+bjTOj5Yol5fboo8o+jf
JFupMjB2PtWB/KT3NTz6l2Q8CBCJ82BHUqiiU+6jfEJpF9kzciFBTbAtw4eWoKVVkokzCgy8n/af
hqHxSTzbtHKePgpQm9NdOYT0yVGbOOuWQDi5qumATnGNDuEnrjnBI7wFIwAxzu6ZARwScS4buWPQ
sc5sXM5mQuXEa0H7sOED2tYH/xKvlmc/STNk66Vn7A6WVvflzWa6eznHNjELDCLxCRdsBAWoqDTb
Xx7Ksl+vZUR0is7cX3fSbyQ5wnCHgp3DPPEFZfVy676Gq/dKqw3VDvQuz6i5r8hM8kIvZtBUVkaH
+Ex7Cmz6LFGQSqd4oSWAEbr4N9t4FNUbnWI7b7FMnsOUvhP/ZrPQxp+WRfh+ucMoe4FLyaxrKmed
G05XAilAtc7AEZLbKo21+IaHNje/SK/YkpI1Uu1eIVL0d9ijEVJWkiy+jm/SGgoNpyZhxX4DG4rb
njS4oI1X9D1W9qhCsWJ3MK3t237a1+UQF2otnUxPe+x70AUzLcV+pRROvPkIy4d+34iORhd8e1Z5
T/AVWBjs7u9zCfqQw5jhm9EBBXjjE1NI/4B3MVK6ycdqnvg0BiK27zUgNZCss3t68Q/81ANW0MaT
eACuEhQeD+kpW1UoqMfN2eTntybiShXFLnk5MCJo3MZvLg+QYrjvfg30oq5xiagZ+AdrNJSBSJW/
0ED16W0DsaTCZaFdYkJKiw+HDEZb5Ob5TkImdXERrnXSitJyb75q4JQswx/hpRPWrgVztTL9cM4g
rQUd+fXSTdov+5eggVasfE8wKoTiowy8JLKTSJkhj6WaDSGX1f+X/OXngdhy/v9S6PN5Ad0xed6e
MW7ZEcJtrMViLAQsn0Tpcv0J7HxrnMTRAXYXYRim63u4JTJrbjKzZi7km/YHsY6gK1B8QCOwPq7E
Vd1MJskyNYk6JI5ZN5HHlFS/NVAHZZ9qdiCC+Po0PlPEEpQPDeXRF2USzFy+TITd7LHCoEJhGgct
rO9PwWVsBbYrY7eEkO3Y95CrHhpUrfGicXAttpkwmxxmuW8XqtpPZ3rjmlKx9Ss4LBLLEZeVSZrm
jfGNNsm4cZ21K/jh5QCxdN89K7Mn2ZPPvnU/yfI+HyIB4wXuRxBwl0375kTC4izSpq/xGyaNCvtf
2vFOwlLaP8n1Ft5a7D6K83tUzeDq3RBXJXy050LmokdEakNc6u/JYY3M1tIFmUWsWmp8gQC/q7pA
KD5lgDDdqO3gQ4nA6Iy4bZzd3k0yS+qDTyG8RiATEUsLcYjUUfY7c02o/m9YatkenCHyIRE0vxb0
z7ztSzIeV29Jxe4ohW1f2Nmx6LOofFHbLwx9Y2nSYWaO+IgwaK1jnv8Y0kVyhbYClxn0rk0nFO3m
qMB0cD8f4S/oqoYVmDrZkBiyLU6EKeHat+qoUn7851A/f3k5n/YEyjg1oLTqVxH7HL5H0L53uabJ
Gllq+0FYbyXrpBWPA/9Y+j7FE1j0/30ZZntkQS4H5Oqnz65QKIoly/NcKYJM9MQxL4yJl6CQkBbO
4Gc4RtTTrCrKEwZOqmW2DI5lxiCdwAsJRJ4xeRz1msc2DUrPHCVMCrY5lerawGXouJ52FH8P8hyj
FhKDMmKvNm/C31vLkKfN3g5XjlGjD/r4HMexmIsn5VeyhSpYNNDG2wpb2f2u4XQ7z8VxBPtrrejl
7+GHjRIcrIm0rO1CqLgcr3ms+4+x58ycsR61rYySpQ+KfkZbdsBCRCWZkN63uEOKnxSPRooGcNad
nHjtcNs+xGLsopa3pUXo4udW8o8ou/Pj5i5h6z2IBZygzDmn+L8x9x6u96gqHw9PuH4BlUzS+Lje
UFqI9dIIQLmvr5gcx6XygQhtJX32Z5L1/xunWuL1wKsydciwaISAI+2CldpM6m+KYzaQ2gL+eq7u
3Xm8GmhzPQExYTFdX6FZOu4IAL5HWB7Z6LO17SrBx+ZVXYEJNiv0J7jjUuqSgcGD4R93LdEl6ABG
OB1PfB3qgWtC6wBCTrEVVEiTiUEwTSYMcddfHl0Sg7lNw0I5dxzTnjHXJiKROwAAC7ND5qp0GAt4
hrY/bIGVnclcIuWFsBwUyBZfUT+mrpy022LgmnnU1PFbB1AO8g8bu/YTxVGUitu1gD0QFJM+xm44
CxPn8xsEl2Yebubm1/rHBGesq00qtLP1j/0x35RM16DxQ3LeMPQffwggmnEKAmGaWh6Cy0uq4RTQ
iSl8xOxzhZECVVuP7KhG7THvz+ma8MozWbKgK8XhiUKptmjFP0hbBegEJoThRjlIIgILMq/5W23o
GZmdeHj+A938TxRqihwv/aZyU088z1oqDy7ARIPublFPU7d0yH1rvJbQDAVd67yMFKlWCLmdPo+2
kS4DwRAdDFVyxTac6iGUppDK/WKuDbb3JmqVHA1v2l/NRVY5YlH+UE2EjtxeaQr7UbXolvN3ypPj
1Og8XXYQknMBQOkrHrVYfEH0CqxaZpaoLUqymFcox821rvH+SHyRc9WEQ7gxH3HoYnvXsCmGkkyu
2zVs4qZIKI0SSo9DpOGtkXO5KFvQOJ4hrWskRJS3FmbZhSEZ08KyPcthiCF20aOwTUMVB9jqOiZg
q1FR/Gp22/5NlVgl0U382GjVLBc13DBBdiJGGu4aWg8OdpT+/BqAZOFEiB9sY4VzWOdCb97+s2Rs
KAlZH1UwBSsM5TSZ5FCbnX1rzgwo2zxsASZpK/EbNUpaWgiFWNImvqMveZCD52i4jDV5pFp+P9ts
keaNkNMY7XMkfDsD1Awuz+aw1hqCwpLOj4EWLNYePOyEtuYvkbSW6SARFy6zbiF/aULyUmfjzMww
6v/SlHAfoTLhx4L0k79RV6cB891Bm/u+fCc8cumDUwz9k/e7j7WISI4Ozg3VJHBQmni56CoF5P6U
C28KS5RURl4ODXBqOqNlNLMdPgAZjPthCMY9arX2epmamJV8sFUmQ2gWE1Za6fTqa6zOvYD9ybdW
80W2qLV7MdS0yFA5DCesN8Q0m4rHHpwjira+Fw0Bfpop8qNC50eYetbVwkHDk8FgCYYrCz0fAhQE
uRIAMr0cR+HrrJKLW45sy9VTIMt8cWu0gjM3i/Gkx7QoRXRKcrf1clxs4XZhHfmCOx/KqnQ/Jlvi
qOF6tkZTcAx7cgzjQfeQAM60uHQohn4t7W1MSdA+TxAApzc+pxDlwaiiJyOemshBc5maxLw46lY+
aWOMczZij5+Tm0k+3SrwDdOrXoQmAsR5RsJe7IBRm10J4Vt7ArBDtMpfIpt3pZcMyJfvXzSLyA6a
UWWsYHUyFGW4Z5R+eqP28JjELs5+NksebtkpzYbAL4VTwY7uyh6/h+0tWN0w0SMrw1Ir9gC8rQZt
09yclZwqW3ctZest1+bv0GOXjP09xTe9WaGasVJm7ybV53LBXd3ObtyzS3T7op6qf7YT5+IBl2uy
A8Un19dgY7cTVRAb+nEwebFYjJh9tpWsMfM9xcvITrUq8JRY2KkyHQGeDJiXA0eoRXKerf6aEsII
wbtE6Qi45pK3N2wrkreQjExjx2RW0ceD11YVOe/hOooZD057dfA0VsBo2QWB+cAgfpeYVt/jS+U5
jAEOoL+ZRBCy+jJhjKx7bS5uzv0ycgwTKkRpVoI62aCIV1+AI4mKtWEFp5QnMUCqlZlOmamVURZr
Zp6f0R86N2bIPh8VGwHHNlXl/F0ID1cb4ciB21pW0WjAb7GFyltxb/impJ6G3v8poqzwFUXojvmV
76s5EspeMTMoNUhNMHMqn8GD/70DV8NjgEOl3QoRUY9xscsi6xC3zdAYUlz/Ynrv79DfmbahcxTV
0QvbylQd7XBaKo6qEt/AorNb2i3Q0J43E07ILDYL3KgQ006lUWhjDbml4+rPEpd0HEF8u6FJI4VI
VWpz9Jb9WIKhhjFndFfjGcId7Bi6BsOrJHfMJ4GqWEHwLA2CClciQfkO8+7mT6cIU8yGL1hjduWR
3Rn2Ml/1zBq8VUIkstyQUvGKowS9/PM+RITyQtiPFtUF/oMNhKkSldKEcUXsk1eIqxSgFmtbneQk
gukgTFjm6ZnEec/Ariqn77nD59iJJu75Go5nGN4d8jE7Q3/7EIrPIan9fA393ASdd9lEKuEe8tZl
39qbLxGT3BbGqZj4038VmAcAKFWR4aQOMi+RatLm5IxeRS3x2czFHuBSZ3BJmEMiQXYoWhjQ3ROj
G9dnMzx1AqlPEqD/ke83WQovFj2YItkdFKHcLbFc1L5tn8SxXkOaaxqgroo6hY35zkbhIV55L1GU
rVnzW9kN9V8Xw2cW0DwSslAYCFgVNoNvNeeseFlMJsz9f8xbfRLhcFUUkdR9q5pdw9OR1RiqRu3o
wY13Vvh0FpQ4jfkj0Jz+xW7vEyTgMfJPB50J4sWFidg1mAXyYkwGCto9rExyWymD3sANrBZcXH8b
jx4MNcVmsR+u9Ai90WmfsLEHvE1tRpi+Yf3aj8JIC8zT8Q+hlJmcLZaphnz0Wgj0ZOjQfhkWXTBX
bLYC++Yn401nsOHVMEJKSMxgZAQe2Jt7koYcFQT1tDzzX4lNNXl2KAEOIc1//IYDo7Ao/odRll7d
UhQ9hTEBjsfIaYq+rx1U6klXBuLxz+RLPuAw+Bfq42IFfpvyvGrbCQQZglNWbNFn9BzT4ewZSzox
YEvm/kKLWLef96aT2bvHN4gpOyN5kJzfVFXKSgsuau9PUTadPEmi6MwSYegsaVpuyITnEgaToaUq
Cwigf3I8ACgELQ2KCOGuaCe14tGkIfm0I1uZ2RR6n9zCb0N/tqhf/MxnS1Y9f4pweB4IfcWqjdOy
UxxFuHso+GFfxekEeSGQ7nEs9WyOlrFFX4eumxLRnCOR9mOFPdKAKf9WJpDBwL3wrSI3cTCO5M5L
k1QM6GPV9KFvnKxB1ONp5knYct2HonhdbMnhv+2b3kiD0Vdl6blUDM1hEnpN9BcrKj9knYOdSEiv
FNWT2A5b4Qs6q0s2mROGstOkAYggL0YLR0wxmaMG6oOrojLqj9zD3b3hQx85ZDJ19eyNUffMV6ql
GnS/0wIAkC/pPKXoJ67DQH0afSCn2TNp3UYAalBXLE8ATy/8iVRpJV2FdKlEPlquLB+NaZ35Grcg
CUgdwCcYeRpCP/KFD2rRtcereMFoHZcrXYatskFC2hha8mo/ysdZ2khh6BvR7LLZrE87+f+ZT8fx
mbmT///TP48NsYsmrIg5/h0Hl1xTXAQtoA1QVO9cn/YIPpXFqbcCRc82c2lDa5nwAAfwA+hSe0vE
8F0SMY1FMNEFq8on6qPtAYTtZ0rEVgs3q7tx89kDIYWzER6mxjeWHXOOSN5rB+pmBCXzzlUqDRfz
Oc9nwFXTcnYXaJksJEpdQaVkOOHLAGhG8OEP6qSgeNKit73LRCn0rtkuw12TQh4iRemuuqsnnHlv
kMr7Mmzcsh4MFXldwYQgxR1MNX4cQ6rKjSXyVhIBt021NOW2+dWhqW0MZ13bqlHBITdRXzgHBhI3
LPkvoDQBf//e2r6BRq6G9pBfd7caivNLfQbpbdbbHS0YkMMpyps7EjBpgezXQ9rj0DQ0XpCDXzS/
pPartg3NWzWErr5dSwtZLfAqxDfDpx7GEK4SdJvnpd32v53lk+IeI4EEMLnerJETcARXYvgLoCy8
TjSda2ciVyvXkMiFBc2xe2NccfN3ksodrgZ2AMG43J1zz3wdNs9C4KbBC5JFNB6VpRhzEtle+5WT
pj7tJbPHBXsM6Q2trhqpA/I8Mll9gszCcKlgMS9OrOSw++YFixsAZXBoqQ7BcaB68ZFDnoFkKVpB
Ry/m0R4lvEU7u01Su/hootQ7MxPebJn/krlu0KrKdTsBfYW2fZlaKS0wbtmXLXGEVollNm3oBmm4
orqi1FcwYEhbWKAiGZDOlxhgX98QPryVsT5epHYi3FgCQaNQCvxSNp0W0jyZtR7kfjaikZkK3Ev/
8irb4e6sBm51TbXskXJ8IBbEosuk2VO2qFJu7X8zMWmNlRpm7qWrJSlIEBnJN9UoX8XU0Lqfuk+D
+BNVp2BqwGzkKxV6Mmo0Llq3NOLdq8ErYc9YdPk1sgU9xlU5sDIFmcGHpkPhdsCifMPX46+l3Aao
l9ahUnYCkt4X8zBptBXTnt6juoZMPTDZEpZo5Zr4VYSL0JU6PcPBjnwJ9pLeG/sR3omwTvNJNGFC
LcKjFYlUy7RmP1dPAEvDUVqczbqQquSR8DgJ9fhReRIaxOya2GT1ykr0PWpvYXdIokdXo4Nk5NHT
u/C1xKA92LpaOFyMBnk0UlHXnMDQo4h5DRwhNy27veV2/jsKayOnLSMzJ70lKpfEKr/BmHhf0UVE
nKtn/L/5H2J3P+lYs9GLTX+Z8/o7/TcHyvLzH96QpzU2kwzeOnpi46xQ+wnYmXG49PbGVGrQDHDw
EpdaO4lBItRYT6FgPSL0iFgdN+N0zaQ6YN5LP0i2EbNZGRJBxqdVuTETGhBlORaLuj+QARRmbuD5
ebQe/2PCAyGnt08+DNcHFUGPr77qXrUiI0PzEAvkYLG2gm5mrcN3OE1x7Rv1gxX/qENXZhV2EcML
A5zl5GXCu92UW4FQjPBcfxa3b6Wj0qevOec8Nej1EWL8e/fWyNt41PGzF8WMuzyowli/7/RpbteN
wtC4U+4DJmxxj8rgNZMUr96+Vb1ni8uxM5UMWxj+lHb74LKFZVekY53afKXp7M5WBQ82+tbJVuSq
x1KVI9qhNZbSBAqZpPlEXQNFAsUAk7fciqhoxLcDr16lF2tMtauutpalajuqMtMrSfFldTwzY5xr
pSyKZ/YOTO4V2+GWN5qmtJb6BbsG2G/l2kaBANHNiOYBWJsBxfjyJaWj+jVsJSQvcfzZeQTvaiJB
mu+CDNhTdEMuP11l6Y2jSuNmiiKFX1LbBbu/uhXfbogw/ushFtBA24hYYtMpKjc2JNURk0HNWyFC
kOBaaftRGCIUajaoyPS0FpZiMhecWettKj90/JVpRJ9yYAoGnsD9+Dbb7M3YvT4iwoSExFhNE2vu
H8mMqYqTdiiP738RCDz1HhCZThGAQQkbVuZP+tBUyN9oDsRpVic5JW9/wzNtKEPfMSIxFPJzz8P7
nBGy+Ms2ZYV3GzrQVPHZwZs6jxvuHoOh0k2sPwXF07/13ECD5WfslRIk/PSK6lnX9JSYFQUUa2et
uRPa3ei5v2BYsVv+vaKxyJfLEXMOA/jJqFufpLPeiZeXJTKFrs83oHi/QK41xh8Ol74ghehZ3yCT
c8qRvDZWXFCIw7ZAyP1o5n47tFPqv2TMkxzd+JgyDYyHFC0w3iBoVw9GoRx53mMU9WxZpKUCSnMs
xlAJfpZ/Oz3Lwdi0a2a8EozjUF8PJxJ9ZAQyb0mPBQ2zczzCEXZvP2p81GFZrxd2kjt3jzebg1+o
u0bHEs1+jt+A2BQG2bJVROxX++sL27p1arvSrkJxUf2ko3zSnMnxvwVe4UOVO+CoAOnStAweC/T/
6SwJwPd6eIbOyozWsxbVNwp24XWERcsKWt4KfkhgmxdfHSsF/YGXyy93zOXHPUZp7kzEYcjJ8+V8
/bBrYN7HMCk+EGkC/NkaM2RzYXCaSWQ7mLzmfv1R/6A5Gwevg/jDXQwfw62O/iVDkdKFPMbHsK+s
OSQqZdS1pW9h4v/uYC9NlH/4u3K2mY1SPdJv6ecpm4BokVwr3cMd6/k5EL7PuZIcWJHN/Log6Uyc
v0d6m5BDMGJpLlIOXNJlKJZHK48EkkYjfZ8S/zPMeBBJDC1b27UPzkM5synkd7zLIYSO/kNGyLZd
nBrGwgZ6k25nNLyB9PdVPWYKnFv4EhH0jxZOOtQ3JT5u/UuEj7woU8ATUKNKm68lD2no0ajCiqxG
C6OZ4tG86UtKXgJf5vFJ0ySoJb6OarYyXBIpDI/fQGr0MgxrGKsOz1BEWX/SCMcUcRDvQrJakyFr
cvabVOoxuT6WpoztSUawx20ijYtu/GhgIEGtEJWRxtLNq/1gZExO9J73z/sVDLZmFKFvQ9Og21OX
TJCTHkzis0pZWSXKxHfmwTKJeJumTVwGISZdkov+MS8P0xW/pVI48j78a0/9DRTR+NjQgTEXPUfp
MwkG328fGq6IAqAIKUIoEQ9+ssvER2SYiwSAEmS8aQyeKAgYH+th8q1fyNp1nZdjMfy/EsxQe0mT
++EgTvU9UMGt3yvvSNkJ3jmhcIqMAI1jmhaJdcYFMGSLG8kpKII82yOXWd3j1bdb7mb+q84iQcr3
8DXgATqWSnQhCiARX53aJy/jB1FxiaZxVZoLWaAT1jCu/NTKzzk4cEjAL00rcunT46ZBsdZidCnY
6C2RerdR739Ro7ZgR62UaV/5YZq39HY3V6Ghf0JDEALVfp1E03MZ4UnKrwmb3GH8GdSM5LUiY4qN
LXFDyRvjK5OV7oJYJt3vm5IIfcuMcLw16N8CGpL6B20ta/iQp0ruDarFxFhDmN7mKEHSCSsp9vGR
fWjwFksR2NqueZ48IZWENzFXqWVkc9Y/mJRJfINbLIgOdqDA3L52Fx7unoq+RjFpupgsz+qEyLjl
WmU3LjzpoB7Czk4TgArtcw+JfkrDvZRwe3LURqLHzNq8HuZsL51QLYFNDXt9IKlKsMULozft/qTe
JzvCsRgC3J35R4iw0d11kdVASkYumYxADpKzaUc6i/k0wjsyB5qgu+x92g/3jrHzyAptYROTpXgU
TxtyAnjawLl993Hp4rY1akvCmWmnD2iXej5g204fvRVJT/6r0/uEZr+1goJQ5C9CyXJPcqcjqVeH
2yKAv5P9ice35oAuf4hRKjhoilFb3lyKhiMUQwlbtGtDD3K/2w+vOa/OIBN25k0fNiOcbgPiM8XD
AvEYVRXVP4N7rAUuzS33YXF3HhpaKVrcxvwC38FvdEp4YmwfFEnpy2WjxwTZX+DCgnOH8BL8SuUI
WMWL0BNPTa+Uw9uZ4hWx2B9TSj+cBaRZK2N9e+6E9sLGBms+u8E7/bPVZiHRnuDFqXPuhH6arCug
3uZicuueEqXzt301jF5OG9s8zL/HtnsUGNPyRmiJMkIb5Nx4ZgktSGoYHuA18+3NQC8IuADDC3vh
20drvDmAJNiW846dsiRKOjDJrYQiliAtzh040zl3YHZNHcnp8uVcdq2hL5/L+3/UXCMpsSUV2iiZ
CMiBLOaGR6gyZ+7+Ujn1Jg5a9tthKvveAXpH4dhXOTkgqXhetGJO3ShCCZPdun1D5qBJN5OmMLSb
/l7DlMEIFicay9/YzC5XamCywCSlwfUb8F6n+mUYtKSTEbLmAtsPtOyZrGVrCnzrEwCBquONb1HZ
B/5D5kPEnJ5emIod0oZ5Ep/apWS2Zgw0QLYcx2HyUEuNH/45ZedMqUlkWeLPibYWeTHGf+KoU+Ym
wS1aZNHMpvO3E6bnjiQFVXL2ZLvvS8xnPxd/XiPhIJC+now2pEe0hdnLiEjEAg9cse/OKx61IptY
KJkEWr9Hvh3L3tDBq/HdwlvgnGi4gx9CfwouSBmjF3UDuzS4XEybHuKdPYGUBrxaJ3ShY7p5eXYQ
PQZXo4D3Pm0lTyZgN/wQYxIwZI4jOFyIzuLqrKmdwQ1CJZAXVsH5VxRsxa6FcqAxbw0Eqq1m4GXf
CPXZ2R4M0MfFmazBYznTVq5lOu/Q9yslk0S6IndVkMFd3nxfcc6byjoD/CrxfqATQNf5VnHaHMbk
PebywqqJuAMvFRLfgV4yebNoinr4WSJCj0Ig22iR3tqz+mOy9xEb+1fcjpRhRcGLjOoJzaQUBNcU
tJaAQATcSyrV/PzvCpc2jC/efQgcr3JNXbyRstz7DoeeJrT7COml5OuXibhZH2gdQdRqOaiUUMOd
k59InllaIfun2fWPfYbtGdfCpCoW5OiiKgJTXRhAwfvKLKU9B8VoQ7DDPtdCkgsTN+FusWvJagug
IstaT1WmwSJfpQ7nCbKroGn2+EA2NPswbAIHuL8+pmiNTsknOm4l8MiI91u49r7fP3yYBSzZD/V+
mtshucRLgiAyxiZiqvWY1DIf27iGFGV0dIH9vZcHHrQHYrogH9Hr2oKu5eXcHdKgOKZ2srKO6bLi
yB+Tc9Fzsi6AUFF+23tphisLBxMkrrMarkymTALBpYdRmnX7ZJAsMeffCm8wn26RRakFtl2Qrqsh
5tEJWaLTCQGBimV4DNYnMuztCXbfOdCJ5NlqNqt0qurmwYWWPnV9BjasvwUXBJM79apDCBnTLSOD
UAXwdUXMJuFadc7c/KHxgO4Sz5LSIfaFE6xdnLgakvek5LUmVor4X9BpWyyZ5dwv5Ipu5DqKY/vM
cekS0009ash9oiYVHjwOkjC6khmOJdIIFVj71nmowtyBA/DqdcMx35JraZHggcaS75pD2CJ2d4Wr
12eezfJlhuiWNH0j9r9pedU4UvGYCoQoIL0kCrjIm5Tc5HPov15KsMo9oQPWBRyPDZ+jnmWbWdWL
o9j2GkDskDkVNLfFgcPk0YfoGswCirh1TsVqAkPr9MVE2QeFCE8gDZjSdYyRyeKyFhSzUR2GaNaB
kUGXgFTyDLH+4XExKIoxJf/9Zcijs3HwVDWuZoZLN9BB9HKnI60F/tyzQlGGh56i4enUni2eSuSZ
t2HW3aLKTioG0TrX9fof2LPY0rVm66tPj05vOWhj4g1vdD88rI2EG3DIawZPOLUZg7r7WJkb4qBU
vbTfNAxGHo+GKly0UU1yJlV5dtmj+w2iv7xsDYeLwMzG6NymTdW3T+Ko9/nEWhmQ1R8Qn6thHUyb
s2JFKQbpHBRcc/kh8KJk01jdnh28D8KoNO3CEIKbsFPwOgnpdgsAQkV2H6HDACsQ/F5xEDfSM3x5
FeSFKP59N//DBmmoimo/IoDCoVfwg3NZI9PzPgWaY0tycRahZ9f2yHk5WdGovK4inPpq/p29slRS
L5fojWfXBx4QVvVw31Tj9O5+6hsjzmmhS7g01SS+rlfZrmsSIWZAa4kmrD7+yC6VMuExfa6Wsp+g
ImJtAHvQHdKq8LrKRENoOsvUBQM6YmoT8QKiH9c/8NtmB22E2YVgYzQ2CUkllPeHIrDk3isgZWWf
A+V8Ogs5uPXF8+sUGqgN5OyA+9gWKE7rvMEfqJHvLHzFi+v9JWllTuOgAYJvHdrSUXM9ggrJ2NxR
SFDcymNHPQhTvQ2r0K1oV7yQNbGKBo+j8q8JdXrnMQZqWDFDJbENVfdFzCWMzE70h/HKhTJMYm5W
yewL+Gvx63YGcG9IC2g+6waj41M/DN4XL7f1mhAz8gPkV2x9ENA0RQoiQs8xiyyKX/e50eGf8RAs
HSa27HbLfuBw6L7JC+7+HOupnDQqRwgsBF2dyovl0/+vz773uHEerVQvB2myTC/JyyLgkld46Xq9
l8dnqQYuBhAa6sm4hTocNYT2v+3J1hggMx6Tjqmmx5k8CyU9pXa+ePHGCxu6oRfSvteHP7NM87zc
k5zCCJo4b8e4uyaPk36wSS0LtodjMmZUdnexi/IEn4syUcHDuHAY3rGeEDsiO0hmSSob31Bzfxdk
ANWBYbLbXapYUfkWw7Xh4cXjc1Uq/FcWpf2LdhEOPLE/P+XE0ibNC42yYmhJWi1bdlsQALijMZQV
eKXUHHXnY6OeHtizLF7b0LTbllyuIwVy3STFfiY9dT9No1k3GBq8gqSx0/BhtSKUKW+RzNueqOZ2
K5uwmcKoxklxPyqsU4NsQ2rxIpFrSRZiLOOcGXv/Xsyd9nG4Eg7f+SMuHIpQCt2+/+5AW3dj4tmG
svovB4BaiY3E88FoK16pqJ4K7YAwp3q9WIrk5WBhgMYMtVByikaw8i2Hf8InvzdrNJACuGD4QClm
zbNFHFc+nXXkX5Rt74Cd9j0MFlBI/phSFiGzzMRsowuV9JwAjG5lbDfFIdCM68+meSywBsd7ITCM
PDzDZFfL3s7fiPLZ8wEbtnKqwxaXi34YvXCVOdrUUtrh3VCNA8w6bqvMmw7S7ZfXr6ebdQtlLUJ1
tQls4/EJvzGQ4+mxEniydYYLIrnwQp9ZzuYuyeXcRCgjFMNL38vZQqykYxcOIqvYjTKL4fj9WdFd
XcYvGRTe24vflSUprX7eutBchQqJ84ZOZO4D+ssZMjvylHf+In/0vOqruiwQj1/jsfWYZ0GTtAWq
h6wLKalla5bPH+8HmsXRVYl/JvpwJOuaKo1CiE1La8t+hhCC4svW655cv33w5WltMwGfS0hpfDBB
3KSRZrbAr2YmyTT7RVuLLE2KyznX5mgk6jkExISYvaU3nvQlLHfliYjlXRJ99fFumnkOnJHKVK36
Y1WzFHfM9ILQzn793w1jw7eMILDmO5GfwBZLUP/EstvUnLXsud8VCQXJgVRv/6QNM42+Ytc7gYwL
/NhasVdF7Sq2X1TWhlgc4FxQ5ajfCUPhX29gUB60C7Re0USt4D4CdVGjo2Ccpx1T6Q4EjzN2cXAr
tQ1JHY0QUAfIseWTCza1CEijbxFfnN3PqTdUbM3gVEtWFGO5NN4obywNw7aYB+FoDnCZ3HjZWjtE
VmFBfb/K1o+gu7+JN02QQ4NdHlFZoZjEiMUU3VzJ7LctunzmhVrGfliRJyGllJrDEUcVtTX4UlZ1
q4CZ6lf1DWJTzP7oGTYnKJyXCDXBN3iueVykjdoFsDT2BeObYTz1O5UqmoYtwOpjEN4vWQUFP9vR
uqtnmr3jUmsvE17Lgvkz5mD6VMJxjZhJRJlr0xAwbWsa2ivEnYelrlnHwZ+gWC2saquNPnDmkD7f
kdjps4hebMvAB+OPU4y2ex7N5mGFXWL4BsBZbRWSxSMXflQ3Y6NTEdxPKAIiYsUj1CY+4wuSOwAL
6CWghapKL6JdNKxrKdafbqR6LexIYo29JchI5RKR/Q3m+ug5FY/HLm3loZV3l3xC++3GutWCiHCQ
3E6YfGP12akc7gJLlAmPrk/Nu0AmMcRIPJQTiyl8W2OVy31ouNy91ATJ3OfX6goNpBdqSfPlzs/J
90n5hSAIQ3pYHDld05VLgvJVUwIMR26wUteMjaapaADsAmRIla07oPEUSHxL7wr+bJoR/+IuSXCQ
y/LFQK6FOqaW507ovTRcIBsNhAT9VDWl9iz/hyxGtoSrrJ4uJVq0Qzg8r9VL+83lGy9xRkf2PzX+
5w0dnmN5xMRwHMuy43M6T62V+sPm/H6eP4FlQ6WlthHFFNAB3c3Bv9I78FYBPMGQPicoPg05Ia5z
3oV4rG6TbjP7nluDFonSXrLHcSyuyQMdMQ/MI1yY7nlgFDpBK5q6RInByF2oRQJAZ0YOwJUbTf7D
IwIPG69hRd2sJeibnBuq2S2CCaC544iMPclG88fcNTvpNzVEHZmcfKvmk2S9DM0GHn3tzsh9+vVE
w686Jtqhw1bbD3AD86t/YrJyRYf1uuHcUgUjcpLBfqk9dRWsNrtNSiSnclBO7CAQFvd9cOTEcjWO
qw4WoaezA5QREM9HylvURP2fZRHWl0mKUa1kjBuANsSGLWIStFLKDbK+V6iU4ACRVIKphzIFf4A7
1CtiLGC8e17YZr4p4hgAIsmOtFh+zXxXFk0hljXgKHrrgks4z/dB+cPEw3g+W1PWxoWA7puVzekP
ZgVSjuq9/TDnkv4ko6w4JHdBJZyEhDJftVsM0bPedS/ULOILlGx56FovtkACSjCvejokDYgAFjFx
YYmsUxllgAndGV1HkE8NQQykiTCg/xgb4GfSh3HuKpVh36kUnqcZgMdgUeYOeyK5YnoxI9S4+vFm
eBFe6JVxC9qw4Oj1qp/8GpNIChg4N5pRU40rFjyxBeRVwxycWPHjZcUVqzTKc5h32E22bEL93ksQ
qG1d3IlzcxIVfBzuLsWs3+U17VlUOZXMr9+rxfx1TBJUSv2NPWHSZQFka1RsXOZ8KV8F5B7Ucdz1
LD8bz/g+W/UmpRcOcns83juTh91igIzcA4peyYFvv7z6L0SM4d3o7v1kXNNCYr1N5xzOUoxbUpyG
qEx1A+acpSTMAUAsIyW5ts23nl+Jt3Po3WJQELZhYyZMx482bOfW2uzCs2z1ZDN3fQk6GzRCDm+y
fttOwBGvSqTg7x8jYydZHbAC1HWXKhBuz3bLFWPSEQCzJdcrDc3RidvZ49GJuQPvGKfRtLRuBCu9
9MqNp2QrAgqgi9iVhxJBcK/GKf7KQzC4dvsVlfiSK/W/FrmSVB77RExZ0HEeQU446gbE0yAow479
IFtf7jnQtFpCWsbISetQZua/WxGc9hcYNHBArmkK47pBMF1C+E5CvGPGJt8nVf+Hqm3N4iIIuody
Uy4u17szQ2sD4coZbEITUKdd7RMTBqXAyXzjVV7yAdNtBZKLXUEfZOtriZN0DUlXGD7FNMXMYGTr
fAqOaJusXetMs+we+jHZn4I4E90X4FL6hXqKd/bqIe5RdSFGJlXHWQjp2BkZ89/QZZS0FIzaVFJQ
a1k31y0R26mp610UbvPEkHelXSWIAIVeBi6t96ybBMETn06AGe/DVHiJXS+4TNIg+4agsuzHlqZA
r9l/VVlDoAoN5f74mnhM/3rGFC3N0gbus+OlK+gRXTyJr/bn+FIuVMZqZGxr65pEoqPzkT9/1oOW
Ah+jNqufbzPnt5BOdxufibVkkdZ+E57zocOOC1Xf3V2FzE6F/cQuXzFFH+vni7qvVIDlPKlp0rCr
GclL/3kDXj7ZOIb9LvzJKLldyotrtUS4Tyn18JpQdD2Ejvk1cTZyegiEnWo3h4SZTZkkU/An3pDB
idwjhLMx34BpIPu3C1+M034SGiSSovfubt5ytWOVrqaEvGdUzF5R6uX6oH4dhjGRhjFcq1JnjYT2
j4LYaBbSQTPKEEnyfj0bvbnfslvl+nAG/MnXlC3jdjBjzdmRRphj/nb82q/2GRACme/qkSiyAh5g
dTjnu7QWoGlvPrQIXRPkiJWNXUIcsCPtyZdk+RAdO3hsu580D+VxdbIAHuGGRSznfqEdHqU9xtV1
1vIfMZrRNeJEVHZcsfuefJZN6uR1WWJnRRS/ROEYhGIPFZrAYvW3P65uwwlcmkoEzg8j3ilQKAz1
qQPyorm345goz6xkv/+BcgDIy9cu7PNWG5Rt2xIBlqNdFAs59FO4PLtTa5OfpVEc+Giz3rs1FDOd
FqKq5LSHQq7J5akBliRqBxblvn1nFIExgnsnQPrnpaoC6Ba9lVLfj280YvT4FWsEpwWqpfnK59An
rG8maJPuk5PZoPvO4fA8yvMbY/3djelxUEEHF9Fxu9+2SRtFHdTRyW485rg15hvEjr818oTrBr/Y
MOPqX5vJTCK/7TiKErOoD/ADuQsFc0q27F9D/EionVLHCePRimJlNTbHDJP/SYN2yIUC3uMfkJmu
+23yR9j9yjkKdNgDPbffSl/iRKWixMYqVc14wk9WHIwYeHy1Yd0QLn+fYxpUyncTsaezYuSt4kLa
8+fAR3ynQa703/LY+ovRE60P/q9jtndTBMAmJnc+G7EbLlySVLNQUw5YRyzls8oeyBc0aU6Xhaur
n5lxPlXuFOjMViCmfCatmjrqw8uZwzaf+Am1KShI4nKt4pAvZz17BZCj9XJgcRsguudNxOHeqek5
EWtY20L9zp9/mNJ35cKGKEXPVgqGACno/hUHR/p6R84HZnDfJS+LGqbMAbVbkSJQnMLJ2/fTO8Zy
5UCyi8ua8JU3FjHWqNvHDIqAo03UFJXvjbDmNG0rY5nQziz0KtE94ZgW8ygnB9JiXLNVAFwDfrXQ
jP9V3M/9Pyuk/jcI7iz2sZAnQXXANtsH+o1D4eCptPLFDk9zQJhWI1k6uNDDtDLheO2yndTxBVpA
FCcnQu6P09lPeDFQ24k0QpdwdcXqm4rpyAdx0JV07hq6u1+YOSR8xXhfVLsJcdgDNeqZXC9B/dq0
q5BPKLioRPVsdAkZxPFK+Z1TMKjLDBKksY3+mJEbDLH8L66oavurOOfWto1yOyCqKs0xLArOVYUO
x7KbS8vUitsfxWwl4yNrYYS/mnJdvbE6NebDQwZNYntLYBLXPxvNQImIcj49O29c480LLYP42BYj
vUeYds7TWvP6slX8JQC3rhv9NDWwCtXyQJL5YaqyAyZIwf1YgWLaMKQslXTpDmtqOqSpkC74v8AU
YcOHzZD/wh0H+6huT/5iU35L8vsCk5RdPnlElrc+OYAmB9fMKFvUzqLY8KuA5AalZ5c+ZTPvurcl
U2RprwolXrJaSImA/leXqbWFjUIdw5o4+GQ3ScJNYUKCeXyFHDWWXwC4OCEqxDnGs9ZZNqGgi924
nbBeaerR1pYV1sdk7tpBGlNVARo32gIl5xRF+qZ6HJFQqNQHHT8Vqlm9BzbzpdtpM5J/gpEPjoz1
2GJn2xgaVthWRI7jlCyWUEjS8cw4DRMxM3qXME/KiYGmxBWz+CS3xrPrH5pfYrXDviBryb+1hmpv
4zl7X2Obx/nYexsmJ4BIoO4SqAORhhvYrL/WOoCQTy2l3oV5zujGZeewRX8u/V75VIabsiqqjVxW
PmqN8PUeCorjUKnJa6XOc4SDHiQRWtFM0qVfVzTTsrpHVPIa72F1tYKhC3irRZc3qJqPaJCDOz50
8Y3cc3W1j/a7bRiMufy/3ha0hU0EsgnQrIdZQF5cqrLwlN1irxpnyzfN6cgO1KgzDqK+ZKi6TAFv
9abJ3mBrOvqcUJAM+tjCpQEpe/qOBX+w/VxMqx+/ZqPtGvlN9SZAtwjOt9sv4B3PFGBWZR/wWa5v
rsvnPtzmnW/nDXnANGC2Q1sRkk9AObK8CiNb1wMicEJfxmNlChCmOdDrNt6TRvMEksZG+6BWQp1l
e9VIq2wwF1odzMje4PGnclTFpdWfxurqusAMRCRXCABE/jf3naMX0ls+tpivQ4xvoh7eex5Ope6W
pPwBX/5x38FwiTQpe5q6LlcCfZfUGNeoqYPb6odBUpkIpG6KUNIXsI51DL3fAIw7LMb8697LRITL
CIDjcTpcxjggnfknXqP8nWLqih9RnJROhLFGyIO6z7qPabamXP3bbnaF0dJty0fuiePvYwPT4Tas
yODy68IebCv14nE1Ii8Crnr9wzaAmvCm8EQKq1DuxnGZ5X8Otaxv4UR79VHrXYDOIogC6BC7XpWT
NeSF5zKBNAyDbcL1JYeO9X0higTqiRn6vZ0V78hCGfH3yikIks3BYRa1iaLF5ScnJzEd1KR9xN4D
d86WmrKw+K5uGsYiZcCBybVVgStLdjyEb/fiJCPtwniFSvN9MbFZf7KvwjdaYohfIjTLwqA2iVlR
vhUIZVMSzeHU3w82zgLjqR/J0u47ZjJ+hX59mmNc/+H6rJRwQIZJns3sEcmKSpAmIzFGRaFwfjIb
xBxdX9MYKLeHrBQ1WPJkZTbk/oPvgHNdADzOHpMtQx92+KkrsC5y6cq3K3qN0Erkdik+bv7m6W4N
3IxjrBiNqPYZZonLOHgvqv3uhvcWlSNN3cBiYFgZg9Q1MPdX0vj7vs3ZFvN87kQeQbgy5l9zOaco
G5jHheg1hiUEPVySmnZ4QKxT1+vJknPf44ZGmhSosnzuMB3W1fAAp7Rm8Kd6Si6OgaHQjqAB0lqV
eVpTA6OC1g96eYlrRhLfSVIpGmVrMnEDRR2VsGPp6PKL0+GPPm+TGf02YY+0iztZ5ctlBIvLhjvD
ZjEZT8Qpaauu4vuUGdvCcHD+QXKmaA79XWFDl4SULaQ36zCa9gOlEDNZ7tW9Sa2gkguQCHq/EIzM
SfhAs8PTDMHju5plbKdf+DmM3Il3LftVPziPuGK2nsz+SmoLvUj/41hkOiE+YLUjDrj632lWW8Lq
84mvuwpiqM14ygFDWVuMArNkRptEgi53amrtxGgbIGDhoXbKrLdfKcmsCdyHQzVxqZoEYh8U50vQ
Aw35ZZT6tbJwIQNyECS7SPhNnyvRejpqAIKZzcMTt0FHSW159Jp26YzFXB703Ji1e1NLoa38cpXI
JH7yJ0DUomslQqDEs22ZaggmvhWHvfr9g+tasqr3ZR9AJikaQQM6WRsXXsmx7zcGC/PaL/CQVyfH
ZhzYsEeG+ToTuEVV0mLRKa99N9wh2abaJL54l+S9dZ44EHTodS7sCSjQgUCZ39rkTV7KvyMh3+bb
2w58ItllHhA6zI5JWLqtToVOINp+YbME3M5YILQo4f2XLScT8YBvsTE8pvxXCF/Tr+iqeN6XW3dg
575Bsw+IjdjVGcDX8HS628yWL5wshDSGy0aw4G+eJh+XssIm2It915rSddecO5I2HwrxUy8DgKRX
QeNipG+yjniTIoHfvdoZDSeeNvhvIzCpoKw7ZcDQQoLXHwriXrIOGoxXBLwrTTN5GkXHV034IoW3
BSo1M5h9sRyZ+kbg7O0RJGzo6OdkTn6wYIs/tXXDGkkPj0wmJmzwWxZ40c+Xqc4rFLwRjuYZ0O1Z
dXLzXdmua3sUItRGNF+q1UiIY4SW6gSylxzqd8UsDDgefIsQ8h/dw/60AfIgNKgF0BPgnRZlNYZg
25ZeFd2qXMp4RIQzEyZoJdvBjqCs9GIjE75tIz5lxIKOJ2WRgvDWjAywZmvbIx2Ey37QFIBPX7eP
E5dOAN6wMsZlTGZn+efv3D3vf/MKsnLMM2CPtAfylr0NBbjwV3EjDNLANPZv+p+7yC9qjZN1Jz7i
IfCsJbPvjNOCt3FwvjJo9l40aGqnyI6ObkUDSPiiMfzQkrM+WXRrfkrif302hLRJuraImJt1/ebK
jOedioBwmulniTFrK39S7OWedeCqGVDq9kQNffSyKhzN9VKpSm6z9BAvEoeCmLHeegki/XJ6xWbn
Q3kVTehquMCWUXhyL+yAhwNKTYWp4J6njcsJdKEbo4bGAB1PVwhPQPQHLeCbJS7DlV72okvTp2wl
2SKHS4KIICczLVEJbsSmy4ElguAsL4kn0t6xNDg2uawlSVZ8HFcSniFk1L+gZ34RCBDH5vtVFxqO
G20nZQzrw4+lxSeosNfg9zvRdsV9OHpSAwx0lyocJ11S+mzIvorbX5v+BRbBLW/+4TD7TzWC6cX1
5KeQaQt6GqMkpLg9/vWjnOYdxXltKU8I0IN6QbvDtDA/9D1u4yF5+qSbzzGwbIthENbgUr89ouvI
7KdV2ue6Kpr3IEXM/ohDOYy/3K4Iz6Iz9I6nZFFF2g7p9b09xABZ2wHyi/QoAIa1rHBmxKAjpEn4
W48rNrO71Ey/4bDlY1Wsw1QGcHQz+z+VnyifRfnEmcsypfQvJtvv4wL187cHhGrZYD4sVm6aPmKr
sPaSOSnYHN2+2LhV5lBrNUyQjWzG53MMOIrFT7BDNsSRWvIyZwpeJrrwa672J9g8NTJVI9rS/YW3
fEOk3ZuwnHGD5vdPvgBdWPwU8UcmZ+AO24XF0ZB1sUM9BSTybKLhR7XS/sqnQ3zO8ZrVUKYgmBoJ
q8hL9kbx/mMUdkFxo73YsSS9MQle4I3tFlENSXl1wOZLkwPs+1Y0cstZ+7RiTTy0hFnmogeERcIp
7Wiou0ow5tBM4RbiokEzzBar1ZUYEf7Gt+4uA7fryQz6mmH5siOLcAdpNV0nSIgQ1Q9VvzfdJQ4k
jZgNGigtm9bRfIHZK5CcF7d/x5RxZgiDAZ2m9odjrVMZU/uTlo27sAoqXYZuZW+uEbt4cfT76kk7
1ba1HXeeyXoQjQFWBZCwYiZfGHl4XpPxz0f/8OWhKSOtVTs8Ztpz4guODKlHm7d26QgWfzjaI71t
tuNm8LLlJ3lmBsspcYQj7zrTQA03NnKClcuJ/9piKcV4d7314QkIFbX9GElyqLW8xfxwlFMUXrDQ
tDOKt+epPO0+BjQCkcESBnBkY6Ao6sIN9XBll2UY2CFn+6ytFUIPdGCXGnxICKMW06rLBBDs6kHB
TGMaJduDkrMuN+5c7fQ+Jcf/7nkEUp8hw0aU2bm7yvO6oEGjVOJkc8WHzPTHqQhnfu5XMDoAN//w
7MVyZr6LD3+mptgxfc9nKr1q63gH7syra/SjslKV51VaJ2KmdgX+PMS/vR7jmS1kETpgzDyLkdYo
JbjFZcKCCbBShclL9yCu1XSkBjSQHEUGjuuu0zm7P9RhF1TZ1JGPw2JVSYZmwyTr76t8VPftsCSz
MUcRdWraMOFo6Jp+wMm69601cVQjIhtaDlvH0mRY91yU8QOwC4Ps0xZ8OwGuSgvLl7E0S0lqjBOJ
XETDsOWRiZx8vVniopZKW1gIy/j9tm8WX3cdVddEA1kH0jawJMXT1k4cG4W8YxXXNWG5JWtKOPgX
2mMDHfhWJS7GQ8J1T21kOKIVMch7Te3Z+ea0FGWQrDZYSZlTxg/i1dx7mtB4UPNlxQ7A1njxB1YI
ychblztsm4sSSHeav5rmwqcrgn1iiEWtEKDrR/Hykdvz6kHQSL5eB4JrcNK+jJ4GFOIxvPGDawJt
9vMsKEZ1LCjbWu/8Pd3Ch+1T3c2YudfpHkIzZMBG0l7ahiIFYQHkQoUKOYcXFw2LLPC7FoxlJKQw
UNkrMrry7Abm8sSlMJ18pzewIYRLGwgtLIPFRbmELbEc6JZEEe8pORRDF6sDcJJOc6WrAjb6eq/a
Biuklph9TCWfhyxj8pHreB2CkcSBbl39FtJd3XVhaC7olson/qmF0aPobuBHo2KR8xwseOuB1V87
a5b/Odz9cHMniuiCqoGkgCc3ZhcsIyFKhUaapBBdTZE0nt1s5/iExD/agGctctDkhhBE4TJnDlds
clan8m+l5+cpUFNsiOLwTUdB/Jzd8wZMhU/Z1omAmdpXWyBFjICzuqPDh2d8PDw4foCvR0ydowNa
gpbG/RNvj7AaIXupXlY1cWgYBlO2Xw7HV56Y2v2K/2uletNyQjTNK8V3cGSGJH1hYJQjPecWIAAZ
XYiDv/3/LfRsxp6Hcf+Bl96nDsjwoBUkEwMQc+rDt9w6whPGprJg84VJkE/cpbYxC+cMjraRWvor
jutlkp07peerrvt51NYr10K2DiNYwdHLnJlEpi5L//Op41SjZpKeKl5EMw7fsvbF0obO77sKmWj4
m3xy2K9eCzEChWCl0qzC4U8TumDr0GYdiZf3rXfmUn3GfcB6ct8EqC3A5PdqcKDlPAD7wBQvz/Br
zxyyw0oD8bCBoYaT02+uKcX3BJOHdWiGuSzsjaXr8o4u++53p3LJ8RRK8vnKxAdQcgJL30iv9JRW
Y2RNsc6soGqaYgiMC8Sj9yWhomYO1eVgZ9H+jzcmRZ619BIDmKVJ5JeajYpWwYfe0d4hpX912Hlc
FZtGIJbbq4M0XPPX6bDWljv6e4Xrh2Eemdqro9kzqQJtdmtSdA493dmv/0WgxFjVSB4ayotpIkrj
GPWvGmFHngV0iQfaxcfLOPb8kGioFX1hRDzGsR/DX2vMK5gcSqy7wVElvc1yLoZ/ELx/4ATEfA+8
VFS2+lZBw6nLR/+RlmW6Bi9FwsKl7eJZEDeLYU4xdtexMJ6htyfxecgFj79q5SgLqTQxOjGcfA8v
3CkRbS1UgnpVpGMYWmvaIW7AzYse1yMniF3mP7LreSAbXd1yZpWOU4oVumPt1WNVm0IN97CyK68u
/Y7QuWkDjAUU++WdNcBZASYuVs1Pc8dqGIQytHTVB2zuKbnBOkWHNV923wtsR5ESJxIcAvbymdXk
Gw2LQQ2caqBJX8z5iLiF8vCutHguiXeNdPjtfTPXU7zXupHbjYDFEL6KBc+At/d7THr5JmIPObxS
feG4Lxci6hGhEge0xcN5KYgKXMUNkVu0JNI3oJtFR2f1Q1erTwj86h4fO1TqS2iWnx9NatiUifdj
84/mOOtlujRIWFaczJ00bOYbKMDs92s3LRHGzDW0FwPiOo21kyqC5reicIDKq0Zz3Lmza1t9v4ti
zS5vGLd636B8tym+z3BACJrjC57JbJA5B9tpm1Q+pmjRJp8eNl921cfztkjRD0WrSvV3dS6U7uZ+
VrQVVzDAokKphQjU4qag8VPmIFjNPrLQstcNHo6flZTnM8GRZu6IKfFmUQW0vXqTU27x1d0iBEFa
6JF16BQS1z+giXDzHwTll+574Bo2FKvx4+cCM9eKIBZSsCYsWsLm+AAE4SigLTX1RJGP+A/xcuLo
JTai4wpxDuPj0QRsLEIf4B1VilNb0D7dVvRPi7O4cgsMgyKOoMx42VzmwpKfIIMKAOO1g+WSaFHU
0Iy5hNLgfwmPrdsbQ64kfZE1cTBUzahRETzTjsjNhVmWxoueMN2mC95/nXNhbq3/wUGlMwChmzL8
v0FE3b/Mp77nIRlwuCjrKU6QuJZ0F8xyrQTjfqGXqO2Z1YsjsQpTwrMY3vUrhb6uKnoDmVqNkrBp
7FPrI80TyiQSBjF7vjgN4qMz14Gr1csM5eA4BNzJ8b67+eWgDE2TCc+Ybi/ufgASSZQJHbnb/Y1X
JL5gNVhY7EUPA6n2kvVY26eQK0uy7vwpNk/2bvLNd90ln49eX5nGC7Axer2hwoCtoYjngAwGuhWd
Rv2KPYybEEISWBJ6j3qaqB7wgCMN7dT6hpAjfjUoHKRZxGTTaHUMSV4CcwbuKNLaHaSf4NgVjXqK
CLKNtZS9yhdM14D8/f5lak/V9WZvhVLtrOXwD9FR7kYLwPvQ1HcJioErkN6AECZce2w0Gmcjhllu
5ru1j7xj6pa0WydlvqdY52QkRaG5vJMt4L/a9aXzNMuXGKN92RYRNMw71q7LWB539UQyXIeT6X5Z
fghguIkRKKaKloXwKzxp4bxzFYjf0iqkgOInU33rN5UBSvzBUPo5cGAsuXoHFm1PN4NrWyET0oUN
0KU/GwfP7g/8bW4uhVAKEnRLHqBK1bWSEcFC5pmVTodCL3p3USPfaLDR5Yd24k/HwaoAgGMaLazm
xJqBWm5Id1CCa77HyURc+a87mabI3l1ephsa1gQs+l+Wd+kiKsA0l0eJy997gSUb6Em8GL3306AT
XBLktC9nLZCsYlvbW+NvH8jG0lLqcUTvgd+5rFGh8JZU/3E3mgJ2CR4VlV71CeN/KfS+LWmKnNdx
4SkV9wCd5lW89e8XWmKLiSsiUmHt2GkxTMbSej/W0yDXU539xbiSY7ztQ7ZFixDNAQUh44ya1izb
gRsOhliIyLbHzzkC4VPThtnwBmBKgxxt3ol2md1ioCewLDkDSbsofKaxHkwOCb9zy+fnUNNTy/ud
MuHxwzDHmv+6NXcTvxjq7/x77exUAaXqGEGIPN0gel/xc8tl2RXthZwTZEpdgLfM42fHuc0W6j8A
l+8YuRL5WSCz891YTgpf7cORdGh5dOEoC038IJpJXtz8qmbemFaRUcU709YWn7gcYnVX4OZg9wQE
Af85olg+GhaZfszA41CCr37ppvbj4rVsM+GSU+mIm+Ax20BwvxcPWiX2wC1xExHROk3OTI0xVkPF
Nq+q0yREX+ZmZtD1mnJ57OAbMiQfPCZMVeVwjQbKPz8uIUa2HNY3mu39wfQ2jag+MHZazU8Q5mkt
O91MV8CnjdD2AJL5VGei+Q7G5rxv4kW6s9Pnxv2EJ+TVMAcrHWCdv2ckPFJMJ0cf7vzMA2TFEEJE
DMyilYYGcJAnsUg5abTEFcNbPxR8oADoXXcKOiXF3hmE67/50ZUMg+VRo4rUuOieqwo6Hi+S5D4/
+YgKwC6q2g/2VuVxG74hpm/oHdHRKz3YcHq3fA4Y1Qm/WKwiuEv9PsOAhNuv0vTdJBR4qlRFvBqK
qeKBCCDhdYf2dUxqwjjMtNME5L4HkMMLxSnk/zMXN0oCzYGrrFx3T1dxU9IC+4bC8LlJxE1iqy1U
pCyTkXXiZhsxkA82si/RyURxJc55yGyGAwXBOA9kJAI8HatFdoGm/pK2sp1usiCDKeciiNpPTatX
Q/oCsYqiEPSUqsEyA0LfqF02Os+DOPNSroSXLKti+cocVbxbd/oFqLQzZYPKqtrVVIicBr0g4Bbr
rK6/hAtoTCGsxeHD420jhPxY7zgyJXzhk23tjioyiPOqnHwf3obKK8zT03jS9Cg230lvhCGkn+CQ
c98+bG5p6oqUkDU9NIsYgjDbo8kUx9stNfdMGbuUTsWXf0vC/SVgIqOxYMsuLmc+wMoj7PC5PO7m
mA/68it+SEcd6mDoelIQT054wLzxCdhl59zJITKbf8j60hnAeCH6BC0VSlDNo3EYrAJ+s3iivr2W
5xQL1HfcVjwbq7KOkicP6aYSU3wNxf5nQozMbI1UWnyY466GWYZXIca7zQij0VUYuG0xZDae22vr
cQUZ5xgpAiBscD9YDNOsAecnzSw0SdLQ+8UqlgmKaWXQ5C5yf8HGaW4oaOUc/9UAf9IfASwaw8vJ
UNLgwLqGvk/GIzA3++XIfoYDHfQyaeIwvfZTKueWIcA6HURxjUPhTsmugVZFmzUgHAcp3ZHH4AGP
CPfdoM/ZQt1QXF23OZhSH2rsMdTWWwwYDzzoUMKFaUpDs5ZYkO4QNXNY+1xFuDkEP5cJV07HBsCd
STnMBvGyDiXqg5gZ+qU/UMeGpt4Ey1G5Sa5fLjeMsEAspFHBe1rsBKpXuCYFZGHF5oykJKFNnodq
+ksQAlYolzQSu0V59wqx3KcvHXiwmyLr34vzeFyjj9wOGcH9o0tSP4ADy70SRP5ncX7i27spmLos
XVB6q7vaUEatQLMQp9t6OBo6u0d9mAkl8ijlpk+FyHYg0g97Zd3MJ+xX9JAdQ+HlMZF+oQhb13fu
S1ASC5DZdiCahzmFt8iDu7qs4869f/swVyq0pYO50WWmeJKkuaLO/JmG/Paa1GQVybH0KZl5TRNj
WHdqNcJhaJ/v0sa/LCHU8+gJaN992COiEBg0Snezxk0dLjZPoADQeYd0jyx/saS2kBu1G/hhzHtl
+PQnR9CSyCJuZw+B2UgrSbmQzc5uwSvPmcGNGkVPi1FdCGeQ7Hj6xFZ7Xcc6mGH23zpBjpgqO9rQ
cqpx8W356zlv5FbBL+GNIkvts9jv8hsbYxbr5jMBqUGLI6X/29oSfG4/9ew5ghEXdXrMDYGCYvuB
tOURaRr0kZcNuP+il6uAGIoEKXHHqwM99ALaJuF8QTfjJ1jyc/sy76KIqZ75p994AIgpipGSWuUx
3TZdIS+rNX4jI8Lk+iJ1sMoK0iP5d+p+vu1CD9Sv/ZqYZPPYg34NoVjnRU6T8tPvnmHRvFVFzJE/
/I5/1Lk5KKEYvz/QMzhdIPrSlZuADwbFkOYLqedK0WElcivv42UPK0sm3pwHFCoXHeoO3HDsG49E
nbzOhcEnyQq1HPhW0fq7OEeCVNB6/U91qTZDLlKUPwGqtUg2IE0Ix9qbGtU5NdknPHlaQS8xQ9ka
DPcYb5eRPXHwDN+FcnVM3IsHSyhoaymT5nYc0Nv+sj1dXNGUyUlhHfK2YXbKDdS4n7LtX3Z8YjnI
lT2LRk1Ms73DhY4NL2fuIUCKqtm+CoXvC24jPpL0l8yggRuUXOTd9ZkjwhqlVT758S+abNpTOxCZ
Z1+/1PD5XqBBbR3eLeV54vJWXVgMDcyj0k39VF6x5nVPFJvpQ2mU0FRN52+MxvFk3HFG5agwgkgO
U2t9+U8BgMYAZ009B52E0NaF0bUXzSrDM/RQ4sQndk/uuOg5o8wDBkveExLjw1FhNKyQBg+GeVq2
Vryu/nN9bZ1FI2sUFJN6lGSsykHncc03iX1OO7Ycs9odxF593tU0LzDEoGQQ5Z80EJLrFhXhniWl
Ip6aghIcxNBO0ia3jiZStMaESut96YsoIpCGJa79SK/4/ST3wzZcEkpSFC9MU85770+6gn/KSCuB
vu24TH8jSIiD2hZLYbf7koPF/1NsRGJRWmrpZ7d8Vuluuo32ATYRikXTOXtMInrEIGgMPvHBWliD
jsrTEN6ramFQwIjbGMff8VRhI8YNzrh9ZZxplXaIU72yuufo6Al9WXKgNE/Jb5lDXUayNgcB+vGe
Y7vUGZWnhy98zLti+0PoVSKcM6U9NnbUtzolxGW83H7LiP36jW/eaGQVWbbTerTwuqJC1ip2rOir
VXCbWegjzl7f9CTX/j+GegRpI7fF9rgNS9RJ1/Cj4KKdNS1m9/02bb4Wmk5Z9Cs2X9o9L393bp0X
c9D3dipPulezuul3LeSAaCAVsHRebBq1vqbHIcxrkEtqOTKhiAYdJSHyjMmjCEJlbluhhV7aFcA7
sVv7NvwhyDg/1HXVon8P2Gkbt1TDTcr2T7rYaFZX9h9TZF3IX+cCkbee/B8WUR532VaSWZb+Csjj
LmDbHakJcc53+qiMgUu7DONrdc2n5nyzMK9iEMmiPVUZi9LfW9fpo3kz66vCTPehFoPSrMQKJMmJ
fco9S1t8wWHzFyZJWbfbSEnuhoAxrO5YnDCauyuZLxiJgo1u4rr1jsVlBEAZE4zQuxl4zsMkkfxt
k6DYzCmr1W/3cgt4VkC5eodsbwUG35VvH/+a/WS8kgclbe9PJXnRFsndb2Sb35ecFLiWwi6HX/9/
yrU1JrOU0N1smB72QF2ARGnzY40+8MYLp4do8XbSscsL91ATJBsyc6w5G6CBf+KTGbWypeC9pcdi
oWFnotvWJpydxmfRKUyL6C/OVPmb+MrzU6HuUdnQvunEPHEaeuWiIUZYVYf/Hm/HVu77rOKQIY7u
iFbXKhizI60Uy4dIRLDIylnylqKBq27R42aS3wrhbFrIHQXqfAuO/aorYGb7OCJhUTwEjSKdZ/9P
ZkSMQB23A4s8Z/gTdkno9hPwNylEu8wx92f5bfAec190SN/AEExepCdsbzzWCJCwszfTLirc2TSD
j+o3NSkmAEJgHc8QkbW9bFNlKEFqrjEteCwJ/+992WbojGwZXr7QrURtLj72V5sp+bxZWgxg2bNf
T96/IO4Oh1nchSbluC3YyuZQXjxS+qk2+XjxSheTYzuZOiY9QuwLZy6mjKVw3WAbuw06oapQbadW
jifpobPDSl5RA63WzfAJ4+O+FQQ2vUivG2hkI9UutkixCU9VQwjzhcd8F8sgsp1FRvjFwIV1CjNv
1KzCdRwvhvOKU/UeaBPpotk7MvDNf5bo3X+WrQ7pZajsRb9P22TM51qP+oJLBO/Mhjds0D9fFbO/
1dFwOjE5ZxqdtbKc5ACXZqqGLDtnbOr2R0xg783GitMJMJXSXPPckUuM9cAnv2H+QYW2w+IiDs0s
5GQ4/tLgrE4ltqiB/sdatAo0R+njusqbkrzsXuLl5P46DZtbd+cVIG/8c9R1vfTMMjkUM5NFxO6L
vMVNefn87z2bVGfMnlV/C1CGyo2Q+V8WdO3ZOUUjeYhOr+xMHJKO9GwZO7SZbLsPYTP8ZCiP24F0
zNqFI+uV6tKCtypLICsmeGsngEb1NoVnju4XGNki8MmtIWvsBUfbWedpYnrVdAbp8atnc/JVRTSN
S+PowwPHRjEEv0PwZkr1Y2olbePg6ftNYwR3KZv2kJzCdA7JwMkbbyNAGdDQ4i/gP2nTSGD+l3GQ
SMYw3uACdpkExFOlapQdOeZdzqVEEvpG1PdIjAolxteAHuL0DIlmRRxL/rCwVC3Uyssq23wvcOnX
RpRa+UhtEq7PVQPW1ilCCRw+RSt+vs2gJavKITon/Uu0ABaVAcBDR/hPDW/C2pGuQVQ1rZiLNB6K
v3m84YKVg+D/Z6O40lxaHQu7bfoS06zgbnxJpUrbymEATUdMD5oW/pbnGxudjEgA0RAgIc/xVobv
6SQHg+UKGPTjE0/rQ9Cwm2f7Wa3Hzs0rsKw8JL5LVqxYo+yD6yb2V4efrCVUyi8XEj+Uzi4C5NmZ
KPGFe2pCikEK716oGSQnbxpzDB0pnFWqbXxgM+rs4WhPfoEcUlis0fPl7Dmi6EKx9WMrLVCQT6yR
HT/asH3IeTz8flIqfa1d7DK3KL6cqeLRQt8lf1B9hXijRC2Krp1+piHANlukpmDoutWeEYlhi/fc
R8B7A/CdnCQMOL0W/R+z7Hr2f+QqgeTLShWCb3FKwww4vwSik/+R6Ccg+ajH+4JONtQSay/iFCh0
Q6Xo2cK9nuNyGbrDNmGORZPQ5DjEIoKMG5wKQyaRZxTcu0yUruhITemGFboNP8AUotW8eEDKNL9e
sMN1K6fNHZRno+1csxiwSUxM58DHyWlISGG2ORYCnR+8Bxwcnp2crSEAwuWWVk8MzJ0hsFBmYNxr
jXdNatoQj5dQSTZIO0yAny5zX22LXHLtRSUAl6tqj4Foe5+LOyRhi/09/nIoFnzFQIywqp8ginff
Vs+8krVqTu/RvVF9NNHx0v1BoHhCi4O3zCTDwkMPyQH7DNtkeWv3VSqwL2p6DGSnyguvE8Ssl6WP
qCIm3B6xwrRw1W5+ythczdROH4bZStEkC8UVsttm7JEHXfEpeDpKOb3tzMCiScPXNxuK53tSV4Qw
BXJ9sVZnWMh4rNw3SGIJuNoO6GnTxKHCDlHT/htODDf6aJan4wObUwwcPf3+NpEPxcragRMA4Spq
r8lKQaX2zksooxlV6uUHHszbsPs36fI+ppTQZih5PbwGtrmRWMTBzN+KY/Qgz00w7+ERCoWgcW73
qFqtHZ6ek2ol/QUiluLowLyUIEiAaUF6+mmoG/KYKJX+tCSmc/jW83mwIEOICxebit+uUUchkvz4
9ZhTaVF0JXHmmuPyMLJO94W06XOjTjRKEvFb7vH98k+igbFLXZ9Wx4+ZZr70bytHRbfbpWZnId90
t6qIPV5R82GYb/wqyVShUqhaAS8gboahHOH4TmSLalOM0e4CNepaW7ghZBt6XK4X9dT4LM/OA4Rt
aGgKNaVSFGVNmyHzbDgr3w850iqbNj1UTboUZSRoXdsmC0I1VIRFKmW2VaSp+jwCA3RukcpgLTAh
aXn4Xei/3VKikBfyfZJ8Sy05hVL0bLRYgnMoyqL86j/z9Y6AzpkzDaDxCbb9L83INVQniR3ogZjx
Mak31z7qEojUsHpedkSIPm/8bHjffUeQy9zsdzYio2XN0PYQXAWuKzpeSRPDYFL2pJh6dKs8Pg9n
rCpkAxLz75SjYRtId2JqDKZA+vMJ0kINa4aXkxwYC8OjXQrt7owyzmf9Cclauqhy630yp81Z6GFX
w1eqxy3jWUxTSFzOxRoBejvfgGoqrY4pEyPc3a5FoFZceMNi1r0DT6nF56C8osw7IrwWTgOsYvvu
FuHQ68/2X5SP0TabY6vBfOI7MNKBFJGK+p3NOZ3/9DjlIlkGo5gDATxZYA0flexqZUZGMGqWL6bM
C1o65HSJ/JTIXOcmtsEwYjxs/+ht1dW0CvhcJXNV8l4XniqINZwUwxvc3tGQDjkUvAgx1m8U7Gyd
jPwNocKW3MghautgZtBdqWGKR1BF1WpyYVTR1zD8W6ha6UwlLq8vjKYq2gSpfbVgD79hFNKmOJ7I
mHxq3NgUQwqnFKVLIwNuSQDhvGoauNvbs7lGrzU2Z6sw6s6JgcXjXGlNm++xUvcNanOeFoKlGCAz
0MQkW3O14z+nVKUJ6loJMFuwJA/7BEPVL970Nhwwsj5A7Bh1JEMgJdRETfkjiZRnABpsm71DciCl
MLiHxDwKHLlSFL1rn8kasGsrUXthTLgKXew1Ona3k2tr2sFYm/6jNWy0zBanF1zVhRR80zz6kKvL
eHdOFXFfuqljVLApnaAS+7OqT5YeVviQXvwErLbQLJ5AvXtvqYrHwhMfgbtt+0ZldmFnl4vbcBEV
2tdQX6lDLPyHh89WRNtqAtgyQzlA+mbsXpu2VDxFVgJSgiRZjNVRPFkt6tYvmWwQcqya7XqAdwqK
w3EXFrYWi1DYbEzfnbXwwitOnr2emGEIiuT3ToPXWv9dAbZ4mVAOgxRYlbzw+e+P0dJWvqXjNHkV
brEGucwKvkzyzQUA8s45L/v1t8aEWB9qSHQOYMgDgSUh2NCn4G+PnGsn5qBhbN6BPSsPpifGBGBp
pot2DInPaVIvIsi3ZDEGzvBj6dF3Vlt8u4oNYsyoka7mezFsglYaNPSpRcSygJ12ofgsth7+MsLy
zvdNP5if0AhBlSHuzZdRORVVbOHoJUU5zjqeNtTA9jk5fYxofYRyANrCtkEvFyjzlxCMn2q35/1B
VUCGx/lei+58ZO3nDI19cXqtCqr4mM52Dl0SEeMB4TSrR+r5Eu2KdZ87a42jFBxU+TMpk90gYW/v
BujuaOqMsgij0DtQcKPvc55TwP5QETJYoUFKshY2V3MwBykAhfHCeeROXLb/IE2PzfSY2OtOBXeZ
vdEXHBDIjT9RUUDxPBx7etLGUZEZ9lOMolcHInxCgqbfqvHy9RheTzKkjSX7eG42p6aZ23HiVRrq
KKH6hzvaWWzlt1ijSXq6IyIHn2Zd/1htlyoRhsdwj27PniFws/LJU5M8bnc+DxLGCzpADgEAKww8
m+Dbrr4/ipTXc9yGln5TRFoNC2CxqMSCddb/F1YpGEULa7QVcIC72NQTfnoaFrKaPE+F8ubv5GHA
BIUhdvOpzr1VhA+fu7xbkdQ7R7xdjsmAzuEJVvUn9KbUp2ETTxwzcabTxScVRgtisDykMUr7XgN0
ig0S5/6M3I8p6tK1HPVRSEDFVJ3ffKGIxQ23n/WIAB61eU3QQBok2DQwycvmrtTpZgZ7lmggHbhO
8dZVhDhZIP3g6akolTMiMka8YW17BEwT46Zci2shrj96oReqN1PZjo2rwR4R7EcjiwrXHSnnnlWS
/OsJ3sHzF7u+KQbrX5tbhmcwI7ReCbU9Fcf41Pxp+ls1UrfeznlKZwBo9hRuSKodInW2Iy6j53/v
/ri9+UnQa0t9+BldecWimAqYKwXbBh3LT4q0y7ZbUC2bkOjsCkPbViWjiaxVhGAm3CkCaouttjY/
9FRe6dP/g6pWMnls1EabZO/QyXY+Qpvnwkh+7vZVBVwom0SBmNMyxM3lGZPW/9PdjUqb1H4fJImp
7fVAFQQ9buHUaws99CJcM+2H3ZYG9v80WZnSuEYLjpeP/U4E7uYktJanx1yl3PsAyUt4SukbP6uX
eWbRJyJqL4I+4FNSznPwIAA1eHA3PZCYMDfC6aycfXuCx3PIp/qcXSDHZ34rKoonqZH0e8cXHFon
I1TGcsoBZuEZ00FsNj8c39WPcmAL86ZVQeNRQxEkQUMrTaY9JrUig8WPbpMxut4zIr9yNHDXAOgk
DMWwkYRfV7zrJUyr8wn3HatAGUBg1KWz/3tGVzWWmhINiBCqx9UqArVB3lSwXyCjq8onPAGFVVt2
oiy/EW1KDaQHsL58kSTsqSUxm5CvqerjAEPeyif2MH1tA6XdNnycE8saKP1Z1OBmcCgBQ7Ggffxb
PnuqBeB3ZfgVdiRq0qjymonznC8hd33il3FAN1xAp7/ehG4VP/+pWdZ80/ghkILdQNHVXrH8Gckv
60jeTnIvbKgO8HoS9TDh8QeznnNXNYSyJgsYhpPTnJvvenPEjOevbS8m4+3xnKV8hCHgH79ATlp7
KISXVRACs2VapJZ6SNhVl8WZKKJRvAHR41L6TDQwHnlg9YbqiPT7aaB1A10gz9J9f0hX4clZyCqx
gI/BiypMEGoUeY9qfjDxtyt6G83zDaRR+wSufD6e4wVQn9BLqOjELfv6AsflWVfGwsy1IocKqod8
1DvMy7aAKCVR6xzgjSTLljGlQ5rc+w9SAormDM5NLpgLsHryg2GX4xphN2vmaZeIiW5Krndd6o0m
Ghr0NPFveIbg7Asq68KIEXs+bqYW+FMYiKNYNFbaM7B7GhCRYIp+JrffrDmdAgFtzb2ZJzwkzD1D
VhPVXRN5v8zg5ODZ9i6nt1nkMYNem6b771DMiEFLocPr9K/0C+44+zDang+FvE8jZKHaTF+kjPkS
wQdPeHmPSq01tsSuiZ7tSeoj7egU8F8qUZOpBpk0bdK3LvmaE8zFaPYGxqqZ0ERF/GeY80Iyonxn
sz56vZFS+CZ9Sb1iv2K+AWzuiOi9P9I2Kg68mqViwFZVNFgZ3C5m4ozSovr8XFFIwNJNFZYMy/wC
azsH/iSCDgvwygaBTCL5STLMDnKiufC5r1xUJ6XZc+Eyqb68ahT+q0AZRZuFg7i1DdXyHUsML+cy
IqGSDCrjPncjXB2ONOcdsawx4s+uTdffKVfaNus7Ba1wKrdAoX79g7OFSl0ckQrxLE/KviY3FBHX
YrFofNW8bv7mkpm4FDeJVaYDRcBCZP1BgD1ELet1r0XI+hvmIhkOm9YFSrsGkaS6+G953hslcVh4
YGz2zfV7wBusAFoCQeowfcJGZOE4dRzciQTOuWssPld6O7caEthUlUUnI+Bxnzpr/o2tiiSvFoot
SJKhSDiAkhOgDSJEmvnISpxZMRFKBOmiaQu8WdtLNNEUhx83jjJ0/FF5u1osjDvI6tPWrKjHOu+n
XRW/Xr9rmgAJQtYnZaiJ7Zx3Y3rUcDCuSCfoDtZDTrJ5SDix9N9qOWBw/xCFR2QurndNts3Q9jBU
3UUJK3a3U5Hh+I8KAvJkveKs33a+eMP9BRy3nO3FXTpQ3t+YneifXkhSq1iVIr+UovtIe3/4hyin
w8Sx1O60/AqCLNnA723Sh3sDevr7Dmi14D8tP+0tiInZiRcb7X4W69jNlxyIszk/ozF1uBYXAFnJ
lileuvrQZ6MySgN3Ha+wz4DR+4GLweeFOEvn1mrqNJNP86wFzni6E1ohSei0xODLTVi7yJSD3wuk
1RnWwwWoMWzM0qodXgGPcE3TSOVBSdPk9aFSJgAnPmPBajE3uKvs9spINuhSdjB1/ado95d49838
cY6Gzp/k6IFbQzTzv6KFChSmyAHBN1/b8Qj9al0Xni7Zsov2sUcLIdWrey0nDcsF5JGdp6hDdF3O
t4MS42ig5kD90vK7A7bs6onWCsZcrFq6BJP7/6YH1PzHj0ZW4RfP9BYmf4Lf4U/hi+TEw5XgKt2/
+Ms/wFh3XE9loYuB5xuWn6BGQw0MOo0M1t2OtXZ4p6IJol2ygGe1GK3vsqq0trg45wzb9Y3rQS8A
mv9s1oTX+lYsaxQQp4Ub5J9ArgGYp3twkHJ1+EkUgnq7f1M+v2K9T0cSaE8RI7ibgpa2cMGRAH2W
EgoAeaHN2c9I21OZID1+m+UYsK98DZnqn2yLEnouKdu/bcBVfkH/dwEKOF6kZnTcvI2i6v4b62D1
8BoAT/kj+tejcA+JWzFrRq7ACP8EAQk6ERBkyi0Z4BtIL60YlhXaplLfF4UCUXI+VAwnaJiTKYqP
+TnG14XVn+PImoynAYnz9H8dioSwJ8TB2XSRLlSnk5UG2DFMAN+HGvAQf+82iJNPExG7ZWyN3stv
LBxMnDBx4DFAI93vjovsVO+WI7uC5FvLGAPiqkDd8L4Q5sCw/CRKtiqUqzdgh9WoS9rChq2drDQ+
XV7dmVmwL/Dl5TXsNYcdBLI4ZZ4ZUeYVjwrDcOyrvcET1QDl+GFjSl9L/DIboKpbLd/48ouCYeQQ
mKYH3bGT/TKWztg3YMsl0rSu/k6z/95NUfWeCETP8a32kZmWhuv9kTYFGxtvUeXLRLAErv7jFG3M
GVs2meWKDvLfWmxSEVrrc5hEp59hcgP/XmjppLBjkggPVh0YGbddGjgXxasPclmXpM6GAeFJz9FM
J9CG+YkSY00aNUgER5/K0PkAxBQTt+L6X26ub0pwosRsnzV3Mg7bjmD1WN7BJ9efWkrN9aRoJB04
W+sR7OxRHTtSA1z5bskwtYJgbGmDiPY+VweBKSfebA9nJWyJSoa2rPJvCb9WgqbdK9skCxoNco0n
3ugwbBChBJIcYbTjcsy03N+SwETLn+siW2sszPaINGbGZgBxrTbMwCQGlSZBKuwxZ8xihFn5VzSF
ePchYiuhBcBg9B0jrYuHfKUn82lulpo6IhctUEethB+xKO6mHwJgooJvZlxG0qvP2MiN9EdCWrPr
8GRRmMy9u/JZBr38+oJkVLj53pHn3rYX1q5fDnP5auVnuyHkBfxS140ovz8/pOO7Mftit8ZZH/Gc
XZ0AixLgz3O/uF+Lc5GW9Vu/fdPl2l7/WuJRM8I2JgGyVImr2IMyCnhMxc1cxbVtR+IIJtFCHA+W
UGjTYdXtZjb/Kw+98eX59mH7/Bk9op5qngTjUZHNDQ0zcmTG9t0OB/8r7307EvxIhnrCXublK+Jp
ajWRilaEBMOCtc3A+PyhqZHg4udqRVu1HIRCCMgNbiL8GKWvcRho972ZMtUFabyY86mFTBFpcpBA
LiQ+PRncEnWy1D0AXjC9oC8L0vrozsD7gDGc21Hkg2qiTVe2wy1DfUToYSw5FquyyyzoNIjWaq6T
WZTBdy0UXU65rLLJu7/a1fWM/lMxPXIT8oXZWfFRvrtPDe3cp8rDbD+HTKIhe/Zqz/jv4jb7JH9W
vpQYA8VCydNp0RrHHH8/QLtogVzAverNll5ALeakpWo3uehIJbBoJL7O4/7XR6Gc6qQh4ozAfqy8
66FsOuT/JzQuwhc8aXSK2IA9O6fm6RQ4BhTqhtqbxf9173wQ4+WGKFRFb7/iuMbMoQO5UMIvn+V2
ZOYVqFx0lI60I4l3WkDyynB6ZzdjXDgvLytXBv/4pQ7R4RKFEWws4Lg8wLB6XVQxUUcah8ZNxHkk
v5Ni2GGdgExoKAi+AuLYSwchd+k/Eeux1Bj5BA7Qo7aHl9/m6+26F+VFJtFWO0AqtHYhTg5Pz1Eu
0EpSOSbnNgZskByvFrT7kiJgzYqVv32BNUccucfrLvcVYm2A2Qfdic5G0FTb+DQxM7JZ27MpiY9e
0z1lACe47KgtXeeJDmq+3X7dohmPG+NWiXaM3vJNcp5uxCYv9G6sMj7iMApSKIurVF19mSG1MRV+
gmnxEkDb2wlvTcDUyWBe4otg+R30XreXfRcZWXvpYx9EyB8PIVQRqC8A81rUyspPEkyBYAbVROm0
yoV9oIwJEQIaHNfuYihTjkqNuJFVyblZdhawMgSj6y3Ca1RnWziW8RwG4tlxPjyryKBSK/UaA70C
x02ZvZsDFe/83J9v7hx3THw7LZJBZC5rVuJgIqGqMlRzdbAEsf1fpqPMmIaGlT2dDNaTPx8+C/V2
oLgSTmnM1p6mG62s3QtiBlMLPs5zkMGVD9NLtmSE1gkXWRsdsoSJe63q2sGA8D+7Gc4+kjP5R5dc
lytyefFlzUw43eBxgW5J+hS2u013lQ3eHhBK3E4nkHHanwTYhomW5fjNdC0f5tk9VCNzarmWxItV
uYEJQkHo+gs6mPaq9fSNubZiw72Z5fyPbeL/WNcibbL98OByd9N41pbnAD6cHDTLFeo5BofDdTbQ
SIb6FT+hpZzbAQKc7jyfKNK3nNyc1DU0Gu+syc8aMQjYbdcz9pvzhWWVJ7YDH7hI2DYD1TF1I0fi
HayLJRQ82ZHX7RcfSAwjwvZGWJmnhh6kesjJ03IqXsatlqXCLzddm94aYSJbUrF3oRfw57PhtKxs
QQeSsRSAW6kQeuJ2Ju5DDlqb8QFbYltUwKc1mCxjRDyPNjOcWllvx1etS6jKrcWpYZ8ucFc23u+R
bDJhbFE8Rw3j8ZrvN2xyvH5LyRWgi/rrLMXVEwnZomgg50QWopuB3DBCBVBCAMFErVcLEt0HE3xZ
zBcCwI7eZLwACbfANj1Yxx/4SmkW5k4ZP9Nia+8f7vmjYG1AdrMKkNVgEdH5W1hOClkbIufDt+ZS
kysSHKS6AWrm3RwEJXhbifrFMgVlK7dJFBhWXRJ//NJ4eT4wn6Mypzwc98gfbKZrj3VZDBFQnsz2
kT3wB7YFsTh5jDlppwLEYeYeclG8kthxyJIOWNy8JzvT5mzk6GsVeVS1+azz9jzgas6WogW6oJXN
CFJZiiIA+uzIzpSC7DjGV9aWtCXH+esclEhwR/AAgjNuTQFf0Dc1T21tcwU56dl/zkJ8t9lw6qox
mK9Hrlm9nhFos7MvNRDTaP/E50BzPTCR+hMViOuKkYXN8Pr/7KyxnebTUQjxUcjHoPNCon4Vp2dT
LTGJsCCh4FWYmY1XUrfCSMCKWowVHuMsSAOK5q77whtAVOFti4NP7c3Pn5gcn0ePR8dRPfNuodFZ
YE03+UtlMsum/+PlSoLmK42OhyU5ub9bLXMPUg5hw3KVawMfLSTRSMfF3RzJkDBv51Hn/oqujDtQ
aYPz5iPIDHs/DvpCkHIqFyLNbnL+E8gul71wSJ/SMaU4EZfZoBl9TUaQp4Ds36HUEu71x2hio4XN
TZ0hO+S0cET0fGAJChZksSDMX03S0IrL/lLWszeJxdNjBuCCB70WTbKKtMf/0beT8GM7liaNWyom
mTy+MHBThJ0GBlI4eUNtruR0Ty8jT02O0GBF97WWQjPd/s2L6Ss1OAh+KUgPZLwZ61smM1923Ehq
IH/cY7D6FsPYmbkFRrYmxAxpRR4uIQIQ8fYtfaSHI/eRFAk3j/7uPArz1MbArEc0WbjbQFccffIq
WxBQM86sh772eUCNOfrRudi9stOK4fX409q5uEa5iaO4NYsyp7p5VXXIZou5GUR85e7Mr5JLWF/9
OxYWFDdrHCsX9ZHkuL4R+JWz286Fiv2TCNnQPsjw0zSCcytB9CKiuy8fO/vwKo92BnfeF4E3ai2O
TxejXe73NnyteAomovv1Csg5vSEsE3xvmATWH2uhwabe7GftmXsDeXUAedWuy7qiIR3gMCgF19Sd
ELRUbQmmqkKZN3XgMef4ie0D+l5S1OVNqZxX4oUUWvsJ4Ce/ZKbWXWy+Z5naQnK+ybeTPLYmFj28
lphvuFOubmoFyKC+Dqax6j1faBZkXDYKfBaRsqt7SO6cdr427qVApEPy+yctiKzjFkfvRYYYgrdO
VnxZsF5NQIfVPhbd6wj2oOJM6Gr1Kk4XmoX/GKJNNXvvAfgMUf4gM9eKHth5zJyV5ni1Bf+mn8SZ
A0ZMe3W+jnH9efXhmLWRPZ7fH5MHPxFOAve0fN2p4CNyKobRl79vAOUldJbxc6bMaTEfo0sRDcAs
mD6zpQrT/uN50qBclz81G3/t7NhtGsx7KLPNGDuuvtuKoZ3odPkhmzx8JypfzryTo4eVWXWfGbJk
G43mdTYmPBhNYgM13JmTk+nMRQk6oe6e+gspMWwZazyxPTPdx6SmqqPrluTpicIuPB06IfZS2Unx
4DBP3Xy2FSwTD2t3aHbAUEU8Dh/R5QAtQHH3stQhOEzcDTd84MvNOAN6PeRI/I9t2uqL5pFmJyKz
1bOo+K/RthAewEjWsyb/NLSUc24d7EDy/OsUnTqyPWFxBpIbiYlgOYaH/MFCFNU34QKl+ahqg/Ha
VlT0RB3UD4xeaE4hljQW3nPQSLlhXCNK6DZ1Jb9JNzaehy7fOWMv6kjMNukyZij0F5gLqqdiujiS
v76XnGcgvpQzb0vvFwbNVtDZwk8gvyLGzZlLJiq+Ak3CG9xUYIogCiqdlfDpGbaKOYjkDAQpzVhg
TnVCtbQm3rqxXEJH2wy6jvgImJNUFJVVWNn5D9/h2kOQ+1gSvNTmJVTv6TrHOK0hAKECUtLK1Qk9
B7RIdYC6hMD0dlPN6RQW0XaGCeBaHZeVakyvPTbauCaJ/zGtQ0IqqgR+C9Km6FM6jiKyi7ywiIVg
4hPjHm+jO2Stcg8QaBxwLBRx8FDYQI//ilHHx8UMTGa+f0Tdinqsknn6MEw3a3keRhx73hX6bUKL
v0CwBWXB3rHbcf8ymnCK4jbntTCzxBX25leEOl+7JxgwSgb5bjHIe/NrgXDCQIr7RKyr5elg7L9K
M7rXxTwTF7G7VQvx0lb4fVS95ijx1wbI1bE9OQe525hJ7KfqXA8USGzf2aYl3647p1ID3L5zFe6w
B7leCqmur5UXojMx9vuall92mVM8lyI5kz+SQ6pBdVoHdvUw5hZBhbh5NFvF/jh8SSXCNmqrcGK+
XAeJv04AsDXfIW5Ejt7HUWtDkYH3DO29ogd40gdQji6EY73fBXN2f0GXP/SKodnqqBFID2NDEq9l
4Aso9zNZUbrwL4jP18mBd2116oFv3+lC2OIc9D0QbiBZGYyNNe2IyAnzhtoRl9yjMSBDjucrJMye
dfKr7bj2HYZUDHdAkGas5YRUZYWqURUfUw6BYuRuSJswjVy8b4k5LK0939wWeTNohu+zm9AEyo3N
mPiuSe38C5aFVaCVsXHKyEmdUFmjMd/qOqkyjFpmFCr4/PHyAuF5LNKtTJS14trZOFB+3j+PMXz7
qRstq/g2I5cw9cZRwAtc0qQgKt9DWgAiQV89+3lol0Tb2XyhL+CXMelgpGnDl0GldJu4hJdX51za
mg8R3eB5wbz4BzuseHm0qpcSXVmQ5N88euq/unqV6Qc5/zcN/x/kR0ChnIayTewOxAgnCecTYujy
tYhlBMWYjkjhP1BfGLki2A1JSidOgv6B334rdfR7+q7NcIxVhY4k0AiXkmn7ED9emHLqzDN9JCaU
VibaynWjv6N/c5jswoXHKH0Kk7O1S3gYrBS9/mw9ZayNynlqtApN/nB1DmlO8Q6WrGGN1uGPkmAM
ZPb3FARevnxmF7oAHWtXj0SsnORDdCnB9nJ205Jm83p9cioRABB7hfk+Rf5rfR7j42+QIkNsyQGq
HCsWi8T7PuJ1xcnI/ZM8cNWHcdGmMpUAIQ6d3fdw993FpKTOVW9kJTH7pXpuTBj4tvdu2BZkRRNx
ETdLtk/adrqzN4DQhbk6j2VHgPX+d8zAIVSpK1qfWHbO1yHK60Fo1E5b4XVCCymYZZVuMFmOW/Es
Xu7H2jm+mYRE3IdSUNotWvWQB8/Tq1tWCk6ODkw6HIb6/oIRpA0KSVDiGHC8gZlr8/dO3C5Y8vNG
zk21lYW5N/qkP3DH9GwZgdjHaIBG6MBgfChcZMqN0IO2bQsSYPJQswCev0o/7d1yyJ7CbYBOuEqp
CLUZe8WKJJmGQZVKN8mguBDNVb/H1dKALjgcSSbreoMSH4qaj3no6t7vLosQtxY7EdyygaD4Kutr
UdmKZGBANpxbchIvR9x/ojsWf3AEmVzQGqpkVLCZRPIvdIefPhmAE3CUf7vrhGfksJRnqLjfgOtv
JNFcTC+XqEPbk8Klfv5CLOaHos3pmwHa+cZaTWBxqLcWWApR7avrfA2eMtWgudmUqsropUzAnkJO
rIEylA2iVlKVSywNq86Q904WQ6jBjddAbSwfBkvFuTuc1GCCTngD8FAlGVq6EzgCGL8qw6OQr9QN
XBuVTW1BSF95So+ioxarOIv2FtDVu7nod5jETJz+SdU7nHpZDihObuAjfomxrfod+J7s9RmZRlih
52P2eTc8bj6XMQLFT9bO/P0pjpC1/PWRHr5EUtVweC0GXJ2t9kDCH7KXll3kHWZnFh1MW+dfkd/p
VCbL1cLx+8vUsJZC17DjqqEz3qBo772lQjPjpAQY7uouhqtkhdo91qeOupTXVhkfC+FMD1KGtOG6
NfYzVuXo93iKEuttwHP3yxvjX2Jpso00Hm7pxKwqGAPwB0h2gsVsutKWJGHIOUrSIkd7+1xpJPxe
4ZjChl1cHQIPgHvdNxjG4WTeGT2xusKLLGcHp5dYZs+yYop24fNwX1dFW1oHmkj0Wt4KXIEPsSNf
gdXOLncN7T1FVDv+/dqaeMhnUXoJJV3eUW8xVJZS8qp+uc+facDksZhPl4zUFAOvBUccN6NvdDS2
qpE7Sq2M7XGhifenXUmImEIQMjwY1HelaWDbVaXA9bzpLTukWE9B1+7eYMrOTujKwCrnz9DtwrwU
M2rkmBZwn3ceOswcUfzmbzPjNVedVQ6KM2Htk+OKwYzjyl0nABuQOLjb6xYZFGu3nkdyMIggv4iD
3Kjkh6N5D4o2oRFfI4eVjD7riIEwY4EkEDmPhx/Td50GdrH8/KbddUUDr+9fb7UxLOUjYLIH1m9Z
rhbgIzghXWjBJcsOvl2v5mesckaiFXfmxl09g258EEesmGtVoNxb4nm/S2HQS33KGm26cwj84BMj
oHia4ih1EnAFhMIQCI8xD34kbfmQT/yU9wr+PhcDc4Gn8BAeKUIjMt6U8K+cag9J3Ad/2aokJPaU
A3DU2z63zasfWAWeOel6Vd7WEVKJsO+PKvLh2HpUYwqcfMkt3oXTi+fDZmmRjlimxo+hoDVUARxC
sJLqM5SsfrGvxdBdyEw0i7T0I75cFj5DnjXE3QyyfKVgTuAOuNu+q+cpe++iuk/FzjIw6gZlxtXu
ka0iPU/X3/2PCUZS6cwbpp0xR7dq2989Nxv+kdku97Ayn8pqHxj2bt69coqnv0Vta6vPPmisXNv+
KIirWWFcIBXLCRmUZbOBerBVETXldlYyyTza1L+NlfJy/u52gjjJHk3zhvWE/BpkycbZzSsE4LTc
cvlSzJSlfdX/efuks6ty2wQMzd3SeexOEoSwEVTr7L5ZHpBExRys5BbI2E5YPI9j23mzjzZGpozl
7wGIfYHYvARnb37W3wKB+MeADPf+AkBDHktl7+VqS1upMats6rfNTMBNEU4cVCxiBCOzt/g4riB3
Cyevl8pYsPGc+6zmMpxOXBfJ2FjO6+hb6cSZvLKzvPQ9/BTwIrpJPQmcjbubiQuCTn9ljI9DWE+Z
D8HzjMs4rkVVcPzL32hv21U2wyggu+fCGn1HoOuu/MhzORvgnmikUV9QBFfiQpYae82LCAjCfHWt
rh/OdN7THUcIoMc2LbE1cxdhy496UkvlNUN/t73TDVDQOHiB4IPqsOkmm1aytUdYTNfFwbHfPvEr
oGLhmRzUejBhpKbtRcewtY/Z6+Gk9MRcRus1xySl5rrmMFcziQKymBhXUX+QUa2K6OnEMk1ARf9N
wJUtfAIj8UhUVR6eW8xnRklBRcmfCeSs8PQU50/T3N70QhBj6OrGjvkKupeCIXRsr2ckXyaVWuQc
9sR5l85eDGv5nADC1BqXXrdAt+DzSHuTFQZiGIIFCuzqZwHzoLBMoFuJw5x/hRKbYJILs6ZRRahI
yQzGPRihPkBM2fXdU5GDYkW1fgBiduoYU7qV1Zs2kk1bhIBZOHGx1loiuXgKqt8bD4/R08Ra4h/X
6JH1wsGggNUZr0JOcTriL0p3flwR6igJxQfLRMqArsDrb7GfKPihZolDUGpPbtbLMXRV2jAbm8ZU
UkV+YOBL3uzTM2lPat0c9eiZFQ2SBEL4864PFp4ABnRYqVG6OTpk3r0gv0oWIPNjdEFzGh5KtVZY
lfqro4FYjwUsZyBImHA+nb/LsnsXCq43g0syZHO5sdZB8yBiHfl6ruoUe+yc1rcTGRH3rzulbIQG
ccf38TCshX3rxMXizUmclPwkRKPov7nb5H835taah2aKwNKZ8QPKUloPU4P/Ds4gJDoQyGTPVmQj
O7alBf3ndumU59zysnmNx/8k2mxX2hoT6qZWGfCubqmBWTOJfJdRrocpzzh06nrBmvEhu4+f808B
MTaMs3BY2aRJVi6lI1cU2aRKVR7tjvml3jRByaSa7/0pljq5DNnU8NnFaf9RWn/W4EH+eKt1sgw8
kptJNJKiwhQIJOQaqRXzYSm0of4Bme9/rKHrCeNw9V6LOILjfv+vFB1fdwCzosevWCBjYAClKpQ1
AxIXdbvBVm+4J91RWHeVfGtLqoGSqnRxmm/re9d0f3g6p3BCtFHPM7BC4Sujs7cuHmZYeSONn4EY
ZMc90pha/NWcAhoyO3l98y3ScRiOiOiasjgxeqyfnKbwParbDGDY2x6RXOUO5tepfSYFO37+jgUi
F0KWi05cs1wWzEvMyHwtyqlRK4HTPUTE/jb2EuyTCuFTkljeFle96/v6a9jbkW+u5rfh7msUp+7i
fcGiYYDksNs7DOwel0wlnxZzXJwuoFEDxt4tkhVgi8Uu1RBVuwqEl3U0ge1Ru110oX5gtzy8TI4a
RB9omVINyXY8+RpTQlckc/rigvlxpshV28VyT62rS0rJcnNOZ5aCMXzxiBYAq8LSJwmwuPvUC7+l
HjFxh1b/gqPT0wqiUuYoSAmq7c3uxCVn3eP/03DYDuwtuAvHChjbYmEGHC2Jb++JfytLbvNlEdtg
surO9DCwudADRYBJhi7f6yjd29dHohPjirAQ3YaqHajOt2T65Wa9iqR7M0hFWeXtU/wXujoGrJgP
279qPiEIvX+7qy1Ga6R8iHDhH2W5bkdiXcwO66SP6XIluJ2xlYb8dBwhBAI7MvfOrcUCBMbruSNh
dycNBZXWYC3mqrMn1ODaPV5F/J1mH98D42T+sQlcHo8ibDouyFW07IK4YU7KIwM0q8f83sSyRjrj
kS23JAwtRJzxA9W4gnDBqlU351yI+F7Kvgyba5apVC/dH+/NptrRcccqcKOuHDjhS7Lh1RL9p82d
8DWAUDAfBm4jYqLtNMgpJdv4eXgSkpFoYL2gM+XJoa124BF74znU7xqBBZHUUsis61cURU07PtOm
UA14T1NTc6QBsjKaJwPbbRq71B3xDJv01Qxq1glN+YjUsLjT7zk6DK8FIsnzdSeMugB96TvMGlsP
afSWmGXTzGzsiK4wAFiGU7YcjOIoy9flb7MR8jz9Cw4mjtkAfljJFDBZ/UZJKLr2OKlRuSTHiP0e
EtvSAJv7KIdJeshtFEHdZs2rk5ZrTCLrXoe5ZDK3xZKmaV7H9S0heTg6keiCE3ZDwpA8rsoof1H8
nHr9kbllKFgO5Q3svD65c8CqhdsA9Ao85ZYiZwwVJMRgRZ77J7NKtEmJZN2Z95db9IGZ9hcjQMq8
qO1dW+i6yaxOR2qzkr5ngim5syDF7E92NytiQ8oArPNfEOTHMmqQm89RI32vKVIXSALNP0QSXzoC
hpVO/d7EqOkEv2mfNuWOqzvFnNAUpoAbX62HasLXpokXTDtsqHs5xJDhS12k7SPTd8B/1uVJYNcR
OCUIfDeKxTAKJptq+YYdh8XlUW3SSFguRNyrUsLHehN64xcB5wbk3xlky5K1V3r8GgMHJyE9ZBUs
J+yvInC3ierVSigCRNehya06JD0kqEC/AMpRAfaZb+ht90+0bgP3jptEwB8Cztmq/k1fvOIKU4y6
Smk9Z3SZLA23lGiJCdMzmVUC8kSfKetH71hUN/h442ATkDIlrQkhTcwJQLUg4OOD84J1RVQ1jZLQ
y7o2YDz69N+VKk7J/NvpliD5BjRMZesNivFOprZ/Xc2SofTy6Ur6NqTKytCbl6nrgCvNqOQZy974
5RTkL7MUnOXyFn5nlOgUAQfsE4JCxup3kBu47uj8R6G8Rgc1jU9mnWa3e/zTt8R/EYr0W6upzK53
PhfU9Uozkf4ScwCkv7UNl8dcS7QIZBmDYIZFo67Ttj0rT2hkHIOJDvgKW+ugOulss/Nd3MAzfxdW
qaarhDqHAHpXpiyq01Jc7bYjXDWNLTEESXhzOmvsjb21CWdJaByscDC9kpDixjPdh5Kj73UyM3zQ
2xUVob3xEQMJh7mM1KlFzqnMbBJv9zjpueotmECRn0jUQ0Buhh2cs9q9TuOmaXt60GV58dC2hAyr
kitw2Cv8LkDXnBAZ9jMejHvRy/UTdwYyaiHb+dMgs931RRU2qNZuVCP+/MUeMYepQw8lAN4DPBBN
Nw1LvA90Aj4w9WGUvDSIChlsYVQQdu0qq8rWssMshqz3lyfGmbOK48gcpMqq/A0Cw1uwlm841jqL
bitcCesRjCMW9ZVhzfC7S42gg6DqTC9bh3q+I/g+Wfeug2/zilrIqENEYNS3RsyDJyiGBtosnVbt
LQaIDpPCOaP7iIlfd6U8iO/4T3hgWchxY7GzqsazObWcisnC9575ZbzpqD3SPBWffPoRNtpOjRFW
6FxNCx9ha9mMH4GWPigEjIip3TT5+rF7IKVc9BSLOYk9eK6FtSFlzAUXs1nBrz9rF3SlBFa9KZPA
YNuvYlnAAG2e5XX3+Y+aLCgoUCeHfEOd4Lit2nokxQubyMPjPlU68GySZogcM7qgIQh9AWnZAv6i
tJTO8/fmKeiAY8H/XZrs6HBxmmiUqCM3PVJRKY0vTs1t9RKtn/M+vSKV7xgGwIQbF9mzE3YMhEyU
KDfVYmxWI3k57Sx7E1SEHTnmzP3CdTIItvGbLK5ErC7uohd4QOH5jOSLStT4XnHtAHr+ieusFir7
K0zyu4s5bJJ7K/Wq31PLe+V46kKtIysStxymO5RQ/O3wOXHDLGty2kCXqcH1LjpFPIcpkFleeLsb
X+2W4oVWFpDaCUfKeiXdiXtbuWOm632ExyEjf6/Q+oUm0sLwTb0126IKSaB5u0Hj80MlWtpWabfF
8/22jv7AK3QI5HfQo0QFEYs0OaaQZTk6NX0hQwHdOS8beCrxniRxY62WQ8xf7DysqosbGbO9YQ8X
Yc+rMTA7RZ2Wpzx0qo48g6rQYkcGpSK2jrvzPvtTAMFZ6qWl94QTuiTFkS5MwVzfa0ETdzhJiMFP
z61XRoT2ObJQSzOycWkSCD9p1KQP9Ovnq37yWnkGwSOUod73CCYnBDLZ2Q06eV7/yK5ea1Pnwy0S
I0+LU6Itcvk3eIkFyWfnGgRVa9zg+azEyxF/BF17sLF4EroM1f2bLJ7cPYKfnKK9/nEaacZxH70a
tCt9jfiKydRLOlrjHCkAnBb52SyLMsaAFkAT5Qzl90t0JKBmxTgnnd5XpcbKrBzs42nj2V32ekis
KBd2rk6aZ44tIJXQ/6a4twfQRFc/if1tZNUfn5LqZoqfuBwiwhVutC6FnBjw6Ljf8IyZhKpAlaQc
Z/J0ElN4Uc2CCOTycO43WIIVpJYBLK9noTSJi0Lq0WZjgOIhC4t7Ht8Bajxbi+GlqpnfzsZIJsON
tV+iOCepLXp6hwq9ymB/WfmQgwRh2fbS93VfBeuN9Z6ucF3jqbOsTsa0XSzTXM3rYLBrEec4h4DM
AxTm3RxR6iPiap2ESOlR5pTfJYFzq6bJ0O8hhVWucST+6A7By9riq9r8DA+ZoKT9TH3o+FKxQlA8
iEO2NGcs+w/M5i7NjZ0s4eWsxmQum1071APKc4RcvlrGBtO5Z9wkUuIxg9zxUEfnTu7FLZXrXVQT
EZ9kTtML6mBBhE79YYRy0WssJz9YrZ+ukCqhyANcsj/EsyS4zhEIbbzaqWVvUIkbmpvCiSDvr+AN
7RcNHkQKTUSvE9LHtesU12leleL4K84rcWjAXzOQANGw2voT0O56lHSIfAzQtOxVuCeuxyxLY9nr
1XGbQQtOUoXXL6CJK/gV9Pk6r7wC0XDNOUVJZYKEE5DjUVfLg45AJMVifUPoqqatJXih1KsO4M3x
tnePeduErniNIixKs1Q0SwHulIwhlOAeHiMAKK1CvmDcTdMt3yCBkqUIvmpUl0ldoVAaxJp8kRSt
ixKUlOH89FFaKd42RYAwIaY4ChE+TjfCTELxGsh3UM4keH/YJ7b30gQLneTgLOafEOY4ulyeystu
GJ0Jj+pYLNYXg8/fz+lcRqZ9KOeIyPX7L8OdJg7Tsvsp4mHFEL4IvChUs+YcAp/2wGpwtsyexCrz
91i886RNJxD+FKtk3qpDuyAfYntrgMjQbuIWUkuGQi5HLMGeMnz87f9PmQG9ImbgDrXqaxnBQd6v
iE3JMdBOqXNxfOrx0anT3pUsbePo2mFE0xtd+eBVxQTj5Lpar8L7z/aSaAvv01zqntPNtIQ2RVkr
O2EI4XuVIzVlQpF80peY6kQu1XbF9WTm0wPaMRzsAP3FtMpiOySxUeCaOJ1bc/76fLCxZ/BhX7iA
yJsR7rBSENIW3ukyuVVZ5puod4RZgWnVT64YgosdCWa3ZIYSIeS5eP7LGHfCvKtbNv8t3SPLCziy
FHwC725FYa+T6ynUPQJDPBp91EAyW8chGltfvfelx3OuxIYAF6tCI29JaLhpMx6OO6CyOUjPMdH/
BkUWtk1TDHjcq7c3XF0dxaEGZZnNxd5SBRGPrwJ/BeVuWm9LJ8WSOpFzDTMHeHZXuUZIIVCHLlN0
kJj/qM0NQ1WdzQnw/HdyOr2H4P/dg3M8wHsgXDuiUkJhE4/gxCOWBWETFN37fqLWNIEswf6U8Fc/
1q8y2TE9Kuuv7mtRdCJVdhIzQuE3ST8cgE0un2qr0FkhTjWvrcVuxkHPi017/ZZzjy4yL7NGRAZ9
CL6GK8ede9g63ITpBOxdQ8ImgFk4WU7MRZTXfKoO71Xe8uxrrHngfTm2xQ078h98pKXzZ8mMx624
NUveKVelxiV5wr8AQ2ykMR+x+1ks8OgKn1gNfLAXsZeVmGiAMafx2CoMpjzF0cHptIcxZY3lesi/
QSQjYI+dErv1bcXxZXrd4VCdN6ygCClcVQy8g5BBD2jtoSjXYgDafSnVtcBPXCI7tDqT9mLMPabf
BKGtRumkMqQXFIFw70+thIBIJGBroUMUjATgg2QXy+KT75w44ajuIXx7UJL5nPGyEtxUByVRZI9I
T5hMLmLXBzrbDqzdPIIJYDCHiAXVTQux35XRWI3Y7SeWhRGi7oBwIvcJNOTF7jNc2C9OY6RcdYtK
kY0gKXgceeQX3qEZRyYJ4i/AjOo+RTk1kU2sRs9pKbY2dO1TyI/ZkOAey6xG79aC+VE/lKcZSZPv
GsBrVqefH6LnGGUYwmsSM8saELH3USN0/ASAxJQOOXGOaNsppSFASUm24jK2o5BXZJiVdlOy5Uf+
dRycnkjPeetGIRS9ofOJOzbBmm00GSnPTzZwVaQSanVg/+DCojS8zDQ2/fpikSHeKYSowcX/3ICo
/D7A+nVdYqWrbhvlLZOzVQ5BvG09q5It5eUiDX6VOuLnjHpB1c9A7entbz0+pmGymlA83leznwjz
mj6U2/roaVizjwQkCK95WVsaRPjdRAeYMw62UIuOF69Wt/UwTUnZ6GP2OxOLrrFQ/QRx2X6iNMVS
ycq+EzgtuRO78Sh1exCSkI2msnds1QxQbM4yBF7FgJuIG/Y+PD8MSvIxBn0CKVNS0S3qVbPBADrE
GcMudVPVH7ad+TNb29C0ekki+lCelxqmj2dpVm7qrADVqenudXJtg76/d3TCaYJeS/kVKIlMvTbg
ezO6oSLmdmV2DtmTVwsDbnaFcMOgj10ekmxtPUKAzCKXHYD0OgmsWol0R9UqYTHZAEG/9CgcEh4L
sXQkRe11t+cOYWZfOas9u4PWX/oVQqHgixtGsPZM9ArbjMsmxbo15xfex6qUjaItL0TIHKT0jL56
WATpjZZfuk9Hk5PQOeQhqGdri+rdOIs3TV9V4KGVI6SFvpZ45UNs1YMFQZ4NPefB0WSl7UidTPRQ
ZMpmucqkYN0qssUAHqhHA8xs+80DgacKhBGFuKDSe3WgNWqGYF6SAMaK5xKoFb6rZdRn20lLsZFM
H4yKnqc1zUDiLHyAFDdiTZwrzkpx2hRO/dLF0plijZFIemeRPRrX7FPlIP7dcbY2vQujCmEGk2rB
+RQbBe5tDniSdrlOC1faSTJm71Nb7ULxVjkXCH0BCArG1+SRahy4y3HBf8laqPGzxtDK1iUgOeJV
BDARVKanjky36+xGYSaGPOfBlmYGS4n8VQSstArFFZMwN6ZsLIlbww0Q9ZlygpMVIbmAakfHX5ro
qvTGdwMvSs0iRi+JdDXYcJrcbnqxrI3F94cCgkrng6pUQIatKfyCcMZNu6yEid4x9kEEg/u+uOw+
7ZmsSIRBFn/LDsG98UAPIHy2EgiRzEpwQNUNnLREeWKV/HiuBzJPemzYzvLxClQ9PueqG4dTQyDp
oJWdnshvLPvI4ShizIEiI+5n3UNRPErpZN2ncOqd9KwKEm1NYnVv/e1d/86GRi0b/QFeF/Z5H5+g
i0fH7ZeRXufqJhc2DFouw1s1BvJsCKKN0DepdKDI6YjlM1fnmOlq5QZj3dFGSP3yfOy2VZf6avdG
6M9hJal8WnoLhllSa0YRZL2vjCYm9K5g9QQlh9nixX27EeTZSV9qQ16ABuSVW/nXeQnum3r7JWOl
zfIwurQDUw+FZ/NTbFx17QObfq2dbwgqZDpkmumPudc8OWwavVjy4STgjdCXk43Cwa8DOpvyJQce
7eM13ZwFf51fUKQsjrFnYOPWmW1tcjaULs85NWa/Q2y/r5yrf8/vQ22zbYZAEgFWhsLboiotKjk5
dspcR/DMr11jMOaB5FAGgkp4DO/aedjSilqP68k3aNVgjCe/rArhjdKwIFlkN2xL2NblneXPZkXc
6SNJPg1gavddgVBwaT5zDSEWtOLa3rVSVb6zCrpYcsbHZsJ7SjQfRKAnMmc21QzpXEjU4uxUv5I6
9BAPCylk21pFz3SWvtnh6Dn7yuMF//KEExoUW5jdlmcQgxjCD8kkERQiR5D/kkArnbmN/qhxEK3A
NLPeUbfsO5mweaYNxq8oKW6Yc69cGftC+ecQrYgeVTWbt7axwdM2RpjKZaGfnjwr905PbOunoRBW
O8yoHChGwzEwra7GrmD7ARd66Y//HpgzjHx8O7IwX4fPjaJ3mXoTp+IVN1dCVgCrWqNMLyFurUH/
X/t+bmL/Tw4ioF7X0UrdEIHBUh/7D2U6lduDqGSK1TYNFbYI+z79bSEDOoiWo8lHSIHwr1RB2OHS
m9NZyB7KAJ3yPO0mrDPSGw9Jcjt1RhAmRpEwr3v9EctsEmQY7+KMY2UnpzL8CUWc5selFh0vKuT1
q3OMIlib2X/beYD1kio+l63trgq3JyP1e+BBGoL47qsJMqUyDOHaDAkBiTn48vItX4aZvvCGrRTm
cIEaHmZCCK9BkEAamqAbfDqlFPSpqT0wos5g8TnQEPCw0YNeZOCwLJMPBgkAZ1AOBIjjH+sAeJ7Q
O0EdmjqD400BSNr9HGtZuiUuaHz7UJD3PjPZRy7h6zYJykuXrml8cG/LfIUyop4XG7VsZ9M1PqrA
PcQua2NAuUMaCFZ0jWgN5yKBH4z++azoVyzZcllUHppX6JksuUNhh4m9mZaKkoFnyCdyoiXLOcom
5r8r/wsBnTEXEk3w/rPVlyztwPB5aS+iqM0OrzW6fU6eDg6zfDAGA/j4LAUKRtr7nTQdV4+7rFdc
lEQSn1uioLTvkOCXv7tSOxyVxWOgYcNc2l2YWi8Nj/y2kwJum6BGYf91paV3EA5g8bCnS1m9qMHY
LM21IW0kF3bDYAiqT3l3CCciNjgCccz54yuwn6j8Hvu3jiqyFSC37H8f7gmTirZGmzrXbbkws/qm
kRkMsPq06MpqG2iZIczPT0UGxN/RjaMuGRh9Efj4/8T91k9k9Dw6MrEMeauTe0rTThTVw559amaW
fs9z+xwqCbbsdZKiYdEVj0IDhJuCIcLlUUx0P8nVrVPgz6oPhYCieNEGd4iNKKY0o2r9bNCwFmRK
jvPa1DusRfllN11IlE43b3LQrLI6r2QNkuUsEP8yYW2NEtc9nM69hQkjqOtYCm7brvFWJc9pRuV+
cgIjrm+C9HFm4ASthe8cuyFe3z0feVs6XAh8Ynqz0QpCWjiuOQr27bkmDFxg/BeeOCneRDds0vll
mm0riWalwVv2aMmIei9YSVsb/TR2NrTYnZYpGJWHHsksTwkh5lEDpUN7KLl94rkzPoIX+C95U9o7
Nko017DEHY73n03QzF7E+pT7UGkteW3H/qxZvI9GYYeHzYdfRpl8H2rTPbK/7lvia66A8xvDMDo6
/1/aggDaXspeT4PrjqF5WO2kcwEci+WaGX9wtcTtE2I9XMg73EwxA2ph4f0J/4dTHVsJy66FrMgU
KeLbk62h6t9foq6zyd06yeBdIWSxMlCzlV9egKn1QoNTiF38xbajs+2uZyvMGl78047GHoQayJnP
Prm/iKe0i/vYBJW/1AI2G3Vna76bVHTQC4eXWeljdaL7IIMpuD73K7/LDnf0rm9V/hYgO3TIGJbx
ceGYCBrb5aSCtuqeF0yLRLULkksZ89nPhJVO+tFGmQ8FMsNNatCGgHGcLNk+HgAFzFG1u88/8Jc4
WgbrL50xueO5q8Xrk3C2EZKmBJm3cFqqp+lugcY09TMuDt7wye/tiEYSZuvK9p7IBNlj2CLbzEj4
bCSOatyrS+9dAjgAArw4MR/2WvzOVV+3RspLv667kLohN+0J09JtY6jTzn7l3qEm3HMH3Ifk0Dlm
zYkWPLv424RR8Uc/UNzR/Irtyu0soIa0SBDE5UAzi9Rve1s04ULb7g2pmxWsMmkDCkhBvAL+E2Bi
64ZOGtjdEN9Z5Hq3JjWHWipYCm1C2ITx7I0qKA59aFkowhua6oZmCjo8KGVCYWdEeC19T6fKSNgQ
gq8Oq6y3Co7l4KVGqn57Hy1TTtNx8yOVfCALYMKnn5kMANpFxpu3S1dTXJVTs7e63QCrSjqUbjSm
oqILk4S24ZiSELQJGGT2wZwYWMnJ+ukTDsEeM7FrlTrfofBMxpFEi+bjxcgdKFPpXGmqrmO2whix
Q3ZSgDkGSfSxOXPh2ll+gN7wgAWlhzCgHqieqjtAjygwBQoUCbi08N3lSIksTx/+HWdwcMUQWhQN
9sh1rwBUaZH5dWwMS+GtGWNlOsq0OIcVIMsMLxT4g7oarHM3S+U9Osfuu5Pk31BcdZw24SnJMDCF
4CTQiETwiYiniav4eaGPe36XEJjrlpF3Ato5rvif+uL4K31AHAocPTaGOt3uxmvjhVer774kR5Dw
K4Be7vJPv++euUuFcv/McotpPihtHmQXhFKf7n4c97WKAFllfirJ68sRMjNmaZrNzvPUrsWbiiqB
zCfSoyb03Vvkmo6zDXFPMSen8akSVVfOYAhdC+/ygQnNPujZ6/WYpRx285RL/g8N/bSbISNwhOfE
P9Ib/WtKFhzSAnPugU4x/drkLjds/VZ+2MqRknAg6phP9zpfsfEV9PLKQrcaCGEijMwrJUgqS+/t
fqWvzUrL9fau2VUkYN3a9DJqHiICw9QL5dvbzKbGMfqhAAzSB9LGyuo61cXUnjzDmGZxexG2wzdk
s5/4RrcaSZEA6vn2ARfXoGJCkwZXJyEPVCoX3hEuF6nQi7wV/yJaNTZ3gqeNo2Tc5rYJO4cDFEZ3
YeKJ/V2dkWJCpBXJbCI6Fdvifolevq0eBgt6hil4GbWedpP7Jtvc8cBCIkLpxzx69yBQpwgQITs0
JfqA2YUUsJ0mLN6R+jdPhpMyWvJqPLO+1xHSCLEVfOhzAR3HbDIfZNDQmn+BIF1myo6adFVzuHEv
h43X4U4yqWhfEn9c59PBx1O4/EzhcPcEo1i9ZhLAcoiP5ux6/QmpHSFfQlSuTQ2+vOFUGuH2Fy+H
WeibeXWrT53QueRfI6oD7n96wQqE8uruoRZRAWoNDND0f9nmdYYYu64e8Ovz5yzYOjt8EMlbdAlO
WIgN5AOiG3GXEaEzXi2NZ+Gx8wC3lIGHraWKQL3Jwawa0pJCYBbCr6Uui6jP0f8LCXl4midqAWg/
3GRG9vV0YAEHzznDoGSZhkjmwZIaz6cRqVO+2AezwR3RZ2UZT9dObJCioOeWqlswt6SWEErVKIIL
GWU8dKCYJsH3iDVr36R4VOGbYW/Olm7TduBcRlnGjZvucYgCg6SHyKH/AdH7XqtTM5lGG4RCtbLd
HLcj2SE/NzBeVzR5/DKEXNsmPbnzHR6gsZPT0Tfj1NOLXrSCShy065RxnjLXnAWItYAYMtQomCbd
xaYimVuQda8hyB1tm9cUSj8NPAYMZzPfsWLnS5ecuAxoo9Jr+e5v21r48rvZt4pxE3bbA5XEgXx5
3QnbcWyreUKWtEOAGSp7nrpV9YasZYyx9N41AsmaBCl6ebVFPf4z6LBX5rWFMGGkGlgTqnLiLVci
FB20MslUUY6VoZR0oTyNxrVIhXNOLsDpfetn6MqB9izwiC4ONhyOoD7n9osRNNikFPOumVEl7fUp
cBklMu0W3F97eE43F/EE8E7s2GKo+NZh0RoiqwmwXBLgXRudunXpj15AhZ8Apn/4b1aB3zzD7EhU
eGj+HbrOgasgURxsoUv57TR56YawEhxqUKZkrW2CilIdi1WUlDb9uNDJHYa+OVdkjChdp+ndSjXs
f2qvShNJGDvpjr9rysH+Qo589/lOIPcFJcPywX1hNCvGsk7tW1L44GVGr6A1VTYhiBqx4pyZJy9R
wQigoQGhh5KngftrJcruajSTjtiIWLNA0jFxVorf0qJtwYXpyVkSf/I3r9Mis/G2BFvb7+vKnbLl
oDyW1LrEjnEO/w+TQMf51hSX6Z99pOA6R1yNDViLz2lNulPxgtGP58AyuizcqMfjas0YNkFuKhfG
kiOSt5BAFOxOZEBqh5HJGn2I/DVXHC7ucJWNCA46QZW1kUI8OqNE7Vp2eOK/8Qm5iGeXr7qg0pUp
Fm+aWLYgLyT+A3XdBAfaQzDBqwef7Y5Sn6TQVvnA9+uj4AoJzKAyIwN1x4OCIZj0s/4Tu268LYj0
0aVv4traePzwTz3cqg5LQpNjDXoE/+jJ/3QnNHG0IHy2cWC4Rf1QIFSj7OAr73pas2vrbGkKx5TN
7Kja5k382fdVc5HRr8+qGBKLtKzdcM1kci2bcADdNWJdOQFSqr2No2qTBOefllWPVzKVCZZAEFCz
Ufh/1yJNcHp9wO+GXCP1zcPciZFwieWZ8m62N1kjXV7w284nqHC+jedQth2m5FzFgGj+zMU+RIJe
quiEynI2FRq2wwzdxjpse/sBhbx19uddsn2tTQ9R6Qdn13xicF0ztRuvzKnhe87w/U8xYX2OWHlo
XHggm49bGSZam1Ybjdoow1DEdWgyD8dnxiamVo9URmXHm5EASWaYu2pzb8II56tKEFkhJBpSLQ3E
T1o5dw3rTZk1j2ajtul9U/aau5WZUaGkBDS3qvhOzaqvzxXb2hdQlEZo7n221+IiXaoZ9vTfMw3S
OFkBK4TrcMeBzJzJwPHB4khqHNBr51hHu/2KQinNtPdR/e+UfMMW7OKYcJApFTtpERa39Km+7fje
v32I3lWloKOv2HUvyMOYWcN9A4WCSX481EQQgUegoQ7mDkj69vN6JeLE8aUuC6auqG1EncGmUzRG
WOHQXFg4CqeLiaBmDS/Kb4oxjpySnpKzJrzRngnv9gne/SU2BHAPsRqAPyC/5MqhUDwaNNBhY6eF
M9kTStMHbJiFABRyi5EtY1i/x79QJIrE55j38jVCDSiS8p2PXYszs81kfPGqw0ILXA/PecXzCB7B
YX8rUo4ILVOv3TYjrFqvdvLXECrt/+/lBTNBqqpsxiD2ot0c8sI+zo5ix5mWw10bni6D90NnhZL2
25hg4paP1WWuFEj8iqoqgJD88PcxEUQYKZKKBkTT4sTpHR8oltD3TOkVfvzhmPyV7LTy6+4R/uDr
Iy6ePzNqt1C3MsCJ3D92ofstRXOvLQlZH2wPaQDF8Rt5KOvMseVrieHuB11BoAh/JQAbWzjoGzLW
LrJvLAD27rIs8WywucobTtlpV8p3MPN8Iezq4vG1KgmnBtXNtqXHweoopxqoIqJqOQtO/T+PjqKg
cRANaBQ8Q7D9Azwy/vl5Sb+QsURfzLu3c0W9xKdzxi3RXr68JIaaAIXhGbIiWlM5FEz2yIB4VmAg
KSGl+Y2eQuLVRfy4vsiDxVhVuMZYUsw+oBXBSwQtbBtn3JMA7uPsn0/XqERlIw5axu2KoLq3unOI
O5c7Zrt4eWUPQzYioZc7BDmO8KtIbbS2O0zC9wNUNachzZIUQTLyhECn2Vddh1Kpbjl7Hdzsipoe
AzVSZm0hpCJvKevjnaGRDc+L/EJBeoiXUsSY0BQUtePk403kCnRFZhhM+jJKEwxnTL3TySIqJSqa
h6QQIKTBC9/ZiDivb80WZvL/jBTytZR+7+VAODARlcRmiRc8G6nnFo2GiudrjTT0yXAxk+ecC/Me
GhCPX8AniWQERU/BHI2iLPjEJ4hpD1DNHFycFVTnJDZ5gBaeLyB1PVnPkLqpkb4SRIODiFEyTM2v
e+E5zZAppjE2OUj1ufJLPg7zrHQdZXtj4PFnH3fq5u0sE0PYwGURTSVM2mZch/6nsZF9jswl/LvS
YpP6QDk5e5aaMPebZpi2RNwkiFsQpWjjXGwxG7K8AygRDT1ItnOGa7zzJvi7H0nWhpwhjqWyH0Mr
QwW6pDgiaFlziAFJVGfLWgUXmnR6Vf+cM3Na22YLhCsOp7OKzpc3uOgJPplD2Kps/ltlFflcz7rm
iDvMDgfo7wBA/JV4v5zu0D5ZNULuEl7LSgfnuyp85TSQWNiu82qzHm7XmuiUEIx1XlQjw15Mgi5Z
SZFuNB86XwFHfI5nWuap7yAr3cZwALn6QOJYGvKzCudXC/vPWbVa2F2cxp1BI6R4k8HVWMcuo1wg
A09OdAkC0Ejarpws8di3A8ztq1DZGniknEw79quzHMbTm/BuP1aStsyUXIRlXBOdIxN97d1cf9au
6AJVVvFmoJlj+RUdHJqIxA6AsEgF72qWmo6x2dfkxjbxglRhFlmDkwga6iZrTRj0ssELGcLtmuA6
qeL8CDoctAgwFYXbdA3N0eiffw9OExGMgz1Y7X01JezNT9Is94r33jJUvXn6ZPt2AjpMfeVRV7WN
/DZkntPS8mJgPwEgwL8HB6/eb9X7pv6vl3lcnkcDTpRwn0oM6G+mLQobgbuvSjiyIgz0IsPQu+Jl
0ixRUR+KgpihTFUzGNlQDoXghgtwEnBIyH02dCAvYwZ2TRKqkmNlNhf6XNVPu0Q221ycREStbQey
byJqIIYgcldwwXNro4t4x6llwxdMvt6N1UYL+7SwXnDG1mfIqjzywKFKzg7ytOepcVpU0t3BarJH
wQrudN2n1gUe6qgvaWeOuDqO5dzh6Q9bF//3q4hKJToFaBWMbrHEfn/Avwuun37vZdeP0trHrwK9
cXfSVP1BCC4TTsHKEpzMtjjK33Javye2DW8+ZAC/tpwO6fR6QTg+55Z+1tritUZa7oD4ORQNZnz7
gqy27nsJa7C/OFwOGSw9YtEAs9/yCnEc59TmGIVpSeHjcrG4BC2KM8HFW8SFZ/gFOoLm3OAJsP4G
cuTVf2DCbtiGMReeWIsDscEUCeQz/CtMtk5BGzi4qEx9nd+e6dPMheWOeCXDPlvfQM9QVjvcc0la
zQyBcWuGIk25JvSbaAludttfWDmyZnon7hFahGMo+1YEgkT/trNaH68oQLj+Jhwe8aqqM7XaY/3X
vNzwkvu6mP6W45YJZvV4Jypqg2TX+8yQKFYYvXLJQKjLzKI8ItNWPIMlAGf8HBqbxfn2e0TtQzoT
zeXx7DmSuJ5VpSfrOrpVNFdGoSox28DP8FVhzy9Vj8NmN0X0VpA1LkywJYFCI+p7Qkj+ndBN7ejN
Off6uhKlv/sKPzTURS4f3a4lUD+K8jWHw3JCd87P2aw7tmQnVZwOtpe6qEFY1nVtI5wH7dLr+aOV
HHtsCJzVtQDmCEdZqe6G1n1nFqlyhZXO0DrZcBhcllGtj0x6ZtAx14nDBditCT/bTsaCgAMf2rxF
LixLKrvjJqrGniiUrgvtCLlHgLF7P7u/rbPfflL36XELQgy1qnY2gqfaGo9lYVzXJ6yVG5SRm7FU
/fB+xWCObwswrI+EVh2yW1FeBDlZBz/kEzZHWke+Qplc228xMqROYkY3wKejYCtnHIw79Ln/mV6Q
GTYmILLzYGXHv4DC1mEtoZqayTQWhu19O0VSQ7BUSL1Hz0rCH2+dIFF1jg440tjN57ZWMJEOAvvm
X2JxLf6EpRmJhjTBOs3ofQyLQ3pZWWWKiej5n23XFIk0a2DiDvLh3z4YtSse/oUNNJ5d6pQVk+mw
pT6xuI0kWYt+FXVVQsG3kgjoAwkhQlxKU5emW2IjgH2eBkj6WIhqRjeWbGw8vI+ZYgYJ1r7Ot+fs
vLb49JNXh8svvJWLmafNqiqgpOes5C5iimzmYERui0to9b4xCtnie0HT5azubaTAHIK8N/m5cTpq
OJbo0KyPtl0wCyQGShP3OLbycSv4pdPMdtA3WD+EjU2X1ajULYYeMZ7VueOh2zeXXwayJiWKw6WX
nHTZabRsgVmrMHR333jYXxkjcv7ndywPAmHfvlfbmKzjo5EvkcREGTf0A64hP1uILf8SVRn0S9pn
WfHmLoDeLU2r/hiN38FutEyIt8xpaZ0hTV9o3wGibM3lSq6UwxRhlN1OBul66pukfjVzLKtZl6WD
Uu53Y/jq1c1qUvh/vL7zrC0y1t4keuwg8/CEbLp6JjKmXzWBFrNnAAPlSmtLduj7P16uoLgEYXXs
LjvEbba+YZZP/Fcw+TFx+VTGKhBdtVi8cW/KOGan6EZunK+CiEJbCy4GLFEjQGOHYWtmFvJF/HdU
+V5th0T0M8Ti/O0ZE0yid+xb2A90GnYH8kUVhPtqvghQFVmkD5wrcLkh4hAJR6Uwu3EfEobwuOr4
Wkot14XTiUNxyjaejIWrYiwc/PE9R1BmgiTlRZE/C7mLJn1WetLwEksT/N/2xOATw3Iq1I4N3911
SgpuFFgzcv9F52uwB3eiAfhdSl0fMvJiAQFL0WBQMcTCgwEXmlgKiiPBnLxuhzm2KYpkPK8zUsUw
z0e7vIdOIOOxSpxVhw39GiUlvnQYdFT0xhnWeZTKeAZNhuKWmCUoPBhEYTQ5MNR1kdJ5jK1Fx+s/
ukt7m5NsoMgCgUqis8GskvLVMOJBFGgyq1kYVkQQ9Ezyp8l5Wb3D/4CGNRvzw6V4EkBynSxZ2Chr
croe2CF1AtnINY06P/jfT8WWJBTfMeba8lYHP22falysbtbNKli7IHtQaZLVd5e7+Hw6c/o2o3MK
gFLj5LYiIULHDwQ/OjMSee3L1ZU1Rbx9Cxe5i12+MQN3T9XIFIbgD6C/gRQrxjKx6KH2ylGYL+bW
/YrsraEQoFIH80yZ8fuaXw61nNzh++GvjdGTJde/3h2Y8VbwaE4+wEP26wjkx9kqmzlzRsYq4NB5
EhIfSH1sF6WWDI5fmP48pdOoBDmZIdFwJ8k66pEBy+Mz+0QjYuSx5YvV93OwZqf2u7jD5k5pqA6X
UC8T7SFKP+JLy+MGo5HI4zCDybHac+Oka2iG/wyV1GNLPhCPfrYkWKsD89hwneCiHtmebLKsMgNp
qTeoLdypQcNCMhS+IvgyEFEajj18Tq5L66wElD4CpDgOm6rISAubVOHrX8WzoS6cAXLbhauT8ChL
yOTShvWgiVJ/vH+ij3P7spxURZw3vOkVRbrU53Wyc9tcdBRMWOowyLDNuQ3gtqzYCfDcwBJcbJ7G
DplNQ9UKaGkUtAYQmplvO/1frgoJmu7ogXfgpRvI+bExAgQxVA/C1rm0aQgXa0MKpy4GFoCZALJc
OD+7eP3pEMvFpq0qhgszgQRzSVCdubXo16mSyn3cRWmRI84xwa3EbLJFz3kD2z8soZH8Eg3PKRCO
qzkV2FICV3DU/PNWvAGsXX8xW4O02EkcnK9cNzWlHTlSUQfBJteMVpXAAuY6f5f4XRGkIQOtI8aQ
xjk3GRBrjcZ381+fXJksgzMaiGiKi6Uj/IH9QcyOJxmziIylf5Digz15c3QDsoD5Plo2I7pXzuP7
bhoJYIMTY6dv95uVP6RrAnHvn7kMrouCo4tCAqMKOGsXTnCLa4GgIsTqT3u/K8HNs793PXb3UbgI
sxZXTYG9C4ajQyLIJBDTiaWthGKZZ//hsIQFlRreFfAzHu3TAszf25KynzeTB0gWGk6GRbfRfgl0
zb6huR7UB8wN/EN8prpQfl/bg0SydrviSnUz73kXwvaD3tQHVXdobWI5HER0sF98BBTMSfiKF26O
1JXw5qNjAt5tg1ycWWVMRwJ/+2HZFEXkMrBeCYTxcb3SdO+sWt8UNvRscltSUFUkPFTQ8Mr1HDn6
l5mwP1MxKsDMdZ48XMbDm9oL4635IHIyuK9d7m0IIUobpi2HpAMh6X6wpwoL+kZ+hlgltWAWY0ce
PVPPtVbvQZpmmJNnPNeW32SOkck5QArm3ytN3EIb66VdH0L/yZV921DH+GdBT/jUSlwHPDxdJgix
CsAJF9TXz2S6l2i/BFcyZ6V2H4BRZ9htnoYXYTqV1WDeVFrvIMAQXmz+iROq2CfA7kYasUA9SXKD
Ejn1Yd7kCMgOMBe4IZsZ8AUHSlpqbB9On2BUsqrD+uUeyy++eECBCBhM527Gz/telvrLKmrSm7df
M8H3b7f83CIs/RkvOYjKarKJ9BffVay3Oin38ruAywmiXBvzxo9a/U7bwWUXgOA4PXBHq+aOHkLz
W0Rnx9wqWMDpH1LXLaDGKY4nQeiU0xMGWNnQ0L22exKr50WQe+g1tl44jp2faZxY2ESjyg92dZ1i
2unTMe0yLybyX33AHkfnLHSNDB5v8ZU19/jy639MSbqUyTJxlLtSD7BQ0mnNL8/fXe1sUmgHNu/a
4lTRXt5vgL49e0XGgNCHvAfJuuAX3RsQqE6HBuSJ7OiqVVVNL2mNpCVpWjoOjWCZNZFANHRXDmi+
wPGSj/JGaWx0UoITHXUfOHcry3eOSmoFOMzjX8ZJWuZ63vAim3vBY4a07fh4dYK2tUMjTIVTTz80
cWuTVQ70qMOxJ6vrtIiJCkqhj7ltm0CKkluhR8kzkocSgo7qMORwaafNhNa7y5UDG7aOGm5zJyAR
hJQtuYY9Hc5JC09noK1A49xCTFAQLFcKcH2hGzf6ix8QE2X7PPFswRdVnnNRakeQEJ2dTfp4K/R6
uNEldw3w2ogGl21Cd+yqt9ydyWGkM890QezNeC9lfDI8CQcspOetXXQvxK9hYeOmip8UPhgXLeQz
ROkByIsKREJIp/9KLsPD7I45jHJNZyn9W9IM3HSFn3PFSoyvg1c3Tw5WLCQoZMeQoMqK5xM8PYlP
j773ZUaGeFDYhzKRTumb3OXS8bt7lMkt2wmFH/4a2sBMJ9jZHkT8/M6h+1WzWQ7Gbd8Dw+LIYItA
+FUrqoOV+tdFqWzoQMAuDT4ZPqlt/pV8136eN7MxfbFVFxjIcS58WskxTg88VW7shCLpz5U7dH7r
9IBlFQ3X7uxUZHAPs4fa7Yju8VJu3tezrcqvLwfmYZ2t58lwK1hevNTgU5MoHi+EqtJIDom1FaSZ
7pM3iyFtrQqKiyhUdCuVllRXgqpABrijRdoMUZEklZNwogy/pk4EFKdm2VGCczxRUAPVEef3wLrE
qo6Ecl3LhWlmGbuOKTxQVZxZkOSzIf1f2nI+zVN+AH0qjE+h+waEXMaPNi7rQUwbloQSXfF3AMGY
Yv8QUeKF6J+gs+KNM67b3vMUtSdGB3mnzlwzWIqeG2NOpHEKMya0L1H7KWdJcXnTTwcP6Wi8dRx0
2sxSz4Q+BGoGCSaMwG/QQey1uqFB0QeQR0gjAT0QE1kBQQgSui+yt9sBUzdmBr9twLjxX9djcbph
9Cs7KEI6FEb0oGtMTf9yHM+0AnxoqV6/9R6OzpemhZlhKaJJxGGJNAtIxjjlKJrhvLW0kHyYo4B2
RhgYmUauZIdUwnMZEv7RRu+5DBVE9712GK7FAlbyPns/qCLk4RkCjp3rL69wwqhrdP07gVHKPIdn
fdDy4A+D8oA7s2TGpF5/WozxyW11Mb7jAXhB6DwrTzgMag16TKMkpElu25XQ9c25jTTEzwJx+Y0t
BkzNSt0LCWuJCSxpZxW/YDLnCr3O7shsuWq5OVRO5Xm5ATcD/6ofZQAarGHLn5TCGbcnySzk4qWa
LNmHrP74of9mdf66guU6OusWrUpD7+4RG5MzKddZODNGJpABqKusxhv/eUv5tO1KUi0S7cTX0x1l
3c0/AMEQnIwVBt5t81xIUraMbsDtEv+eUvpnzBoRlaNrgvWjonAMHaUaLLeHC5y7tee3RmJs2sFB
872IHIQ+cYieLukYOyx8X3CfjYfkdG17FgLee3gro53qJqQgmb8DC/cmbNCJLl0fv/0gjBoBN/nU
2M+gpztm5jzdxdQpXlmU+NWR9VK2NXEYP2iRgDt7iZSLDVnoEV2a6nUJlW1IB0GX47IxDkgZaqsL
ixJyAFgEEroB7sIE7uZZ6tom0zjdkPgChX13J7ICkeV1HvgASBKokvpHgqnHmZ6TUXjYT0URRJnV
OnzCa9DJP5u/qenGh6gJMfQ2n4/HF15UWHkAeS3aE7Cdd6Wzt71HRwvKLDqJD79uCD00b/AYjsYp
xLZ1kSQjYvCh5e/e1Csvv2DceF/ivSGWrpYzKxFY5tGdTUyw613JPK3g+9B9SkdCgXIrYJwOAhHA
MXbq6cZHah2JZHGomsxXVqi1/9Dtqa6TmY/H7z1w98m/vkGbKjRVnVM9Y6tHdUtsBaqwpGAhSXGe
PKWo6Bc4FtQ/XbO1BLWPTpc9AfxmirxwIoJ0xHKuIUFHIfcAsyw3EPqY/GPugkz07QKGY6cX7ady
yu23d00EQTr1mifut/K7CwnJ7pZ+QF8HC82rznUwN8qY7RIa5qE4CakoE7K6sOsjvSAmCEpF7E7I
IOyf0mF1j55K1Kn5fHOvaB15UO6l5HYzqKd5KIytANRRCRFCvs2KxgGYaSN5SSGz44tCSUizrjNL
0XRKIzbi595UzPFp9EIAtZ1WOa75YgaQzOrVZRAZ7/lKUKeOLyf/QCtkhUfFRSR1KRL9hVudbrJt
zB5uWWVTiYkBcRxb5nMZU+9QnJZdAPoy2OBd5eps1ULSjJe3d4LYfSLfPrDaI9qxd9ZrkKAociBT
phAbVNsAWAZ1n4+ZQZLHdU82659cOA0bmirnGdtqHxTNE1MSIHpbK0GOHpcRRMwK/JyIHG2Bkqg3
YiRnXKxhE+zgU8vBfX6TmffipPYyxYUuGzyHePBh3VrTe0WZDa0XVZ5zC1/Ec9eeNtFapd2Qcu24
7S6k3L8bAOm9cEYRXN0XBzcDs2qiwaNddLJYJ+zh6Nclv/V/tQ8ZKEECPlluVxpI7F7e32BU3aft
lro9hkNY68pXW3ZFcrclC69vt0j1R7YmMzV011FSpyh2zfH3wG4t4LzGXwMCNU/oyymexRP98FNi
JdjyIUmWdyAVRutGo95rgAJlvrDDVTPF2Mfze6Xy9lP1w+2NEwb2l0/+0FRNdOfL3EZbs/KiVTTq
4T/kR1s4D8rzN3Jqy72Iynz0XtOXEYC2AKkOLrWMzyMqUTZBF8Vpi+FdYns80E5mf2QzgMeqwg//
acFFrJKrquz422KOsWr4imH0r8aIvkaU5ARaffb75Nf8quOfKuq550a0iYDquGGNNZOMIQXPCX8Y
VSKy2VQWxf0T42Z//KSHIIjtiVBxifTt8gB5PuZxoX+2/fuOARWT6MTnGD8PDbpd62qQBM5AI9+o
Otf/kyqoDo5/iv7PFKQ61PhmrniNHyEAGnQAvebylb07ie97mLl5QIEe7TDbf6SnfTyV1mbX+0mV
iS7lRZx8kzPcNyt2kML53WSmIw+OGsFVOKmojGCRbeJDtvoWDYJgHT0gkbyOw0NUVXhisat52Ogp
YxQ3xOQq2ZuvTGf0Hd4LactPmSsGc+F2vBAdVWZGqsIxWvsUYzXv8/iLhAPuNeqMRXdFFVYlbbEd
mk9uLWAvIGlT12i5OXB18LbkmeJpsbBMExuglP5K/P0h/DUnxm6do2B29V/UIfoT9aBDQMQlsKfH
ZkXUpxoeHCT7sJRegztzkSqlGBWH4zj4yrk6O2kTxBxxELJYmNdKlxRToGH2oL+7EW2jwNrdC/hh
obsTJaJMdCIoFi87P6gk3acLNFrePxCEmfdlvE2yndnQQFJ9FPi4ZpoErc8+8vHJyudNGVjDsSim
7WuFSpWx1PiYKpW72wAcv75e2HvE2Uhp2n9URF/g2gMHg2f/mYE2OPj7hDNqifwsyeFC/ZOtD3fH
d6Om+diGvVi5hS02x/gXIVmNzW/4hQChH27P8onajtwpvhiq3E06Dpv74HeePVYMudxfq49EiUTl
6k+hzpXMoQzQOErjuYIJ8ZHl3rkMIuPvUfPqHwDizug2pN9+rSMdFYS01wfqTnABpUNr2VmwzciE
RbQh9ZASWK3eKTC5q9ibzwBPl+5ck9J5+2M7sVYL4MrruTvt3kDr2/gkmVljGQdlQDRL5Nx/JsKH
sO7mTM8olsGhyhGCl2WuwToDXqai/Dkf4A6dPZX4jGkNHLf1trPIR32q8EUZDSq4fo8+13mnOm3w
ZUI8V16HIjMo9g7WKKI9kZLdrGdFXBjHdvIlvYpVYHTrgDzDFcTwadckhvD/H3yaSTs9CTh3twAU
8/KI//sc92HG0FSDYVUnkCOaJmiAREuk8EZQzpVnc/dR2/VcCfYj2lTt/gMEpPUadHLkTIBjWL17
4dSmsE+T9Yrml9BEoaYQ+tTYTOQucOLmVrWQsOgTjCQjYpuMpxU7Lvt1EWg1D5/i94XuxU2mdraL
gAZP2PwI2rM6RosHMIOoXx1z3SNVUgUso7vLM3P+EmPP1GOnDEEcDRn2hqt6l7/6vEAaqkNJtLIV
bPyLBk/sXBuKxP0I6omW/jhU3VqHlPCATWOE1ppuinCyWkpyOSoIy7ZWeSQUfnp9uCesh3tI/IZU
XPrL+8wT+sSN/4PuHrMNVV+lmZBzM81KcyKa1JsSzdzZxYz8ttgsq1xruetVrdbl6FaQ7F5HyLgh
MYfZqg06sNf5FlCxe0d1JgcUiQKWWAy6wkVe/5dGO5njXY4EzuMmfhR85dsd9eQp2f6R+eOvbT0a
tybBuH8kMyIfxRXwIKbTOOeUax5NDFos1gUwH9wDZVJV7/iis25RSgwIpFaQIGm9O0HvaeOYg0O/
D/PRnpwcw83ltcm5AFvwyoS3JzU5HnEAb87fD9Nby5n5GRckHcGpqwjd4LI9gTmffwWGw5hE72uP
e1k5e6xh1u6n3U/5HUMAMSY9K04IYGb2wSLCQg1CSXcxR2ljiiHNN8Os4ya8/XFFYPrBHTTalIOO
TWVrXh2kg69nZmddIpGozxJ8CNPqsJ4cAFlmjNWm/yvhCk8qBYp0P3IuFsILlmHsVzjNGWDcUZdt
LYFcxe98Vlmsv8IqkcAY+gGDaUj6myBsQ54C8ExAE0o+cL2L1ND0VRzo/g7Qq6pal5tAJz26Q65T
W0EFiE3oYDS6zTt7IyIWUmz/p6goL/d8bAkAD6G7JLr8IPhORVjE3xCnO+xPiQrSc1xhC+zz8C9Y
4M3f9CFR5xKD8DXODqld6fVGSAlb/dY6MYgHfd2+VFkuUoySpO8Zt5iAWoNgqLd/3varbpC+Df9X
OI4j1DVjuC6KQI3khwDd/YnI/zPlQ4fxgUcqq3Nm2iLPGDvV3U5t5hWT2pMOF9m/kcdfaH9vadU+
aDhqA0VqDFesfBizEXMUN4w+UdFPnMPEbB5JyEmovss1GilhfHVddEAdWQDK6eJQOSchqSGhCmNH
0ta3LSwj+ES+vcaIBsSUKQLUV+xmfvqvwOJlGvZwy33Au+N85tvWNEiYLws1UcU5hXsWKha/VzXo
9SazO6C2tWx6tosb+UHODylqzEPHeGyqNPAdDm8pahNIVegB6zwzI0H/zVWa0rhnYPEuc0y1A1sL
AmHzBnDJFdZkeJRdNK/5Auf7sRrT64ta7/ZCtHgKDpJFe0vUirgl2ndxmRnWz2lmioYWgoCWu/ZT
zl9bJGE3ODu58wxetLPjkl2sQZiocB8jBOD9Oe9TlQOuXQ+Cilj875b2TWoDlfHU1bDXlPGK51qZ
svr2bBlYw2eKueH0DhW6YJhsWYj2Ro5TF3v7zCLONmO/SguFQOQuWhQs6bj3WCnapIS5LpOChAR6
gHx9ZmKfP6zqd8dMhXuqNvQABBrhJ2d9BkiHU2o487ItCaapS+PpoFtJQJ+fAtJyl8PeMsMWVu/h
jDzkstXSXGTaKmYpmLh4mczdA1DdgJ6qHoAWCKtiQtiiU3Y6Y6WzEnAb2JfWdVzfasV2fMJMAfX8
48IYY/IWzC93oWsgVdAtuhGwukoqSdjJ5dIu03oC83AjcbtqmSJTDv60I7FpWfssXoX5K/AetTaG
cZZZTROBYko9lZnuD+yq6yOWRBvq80KKCwJPt4bgCSiWQE/1C2UFwLHrWfoLN487vXrXlzniCMSk
i+0EfP3srtEK46bZTkX9dEavQ8avrGYLGiVpiLVStz46+NrnofbgccNDqGH1FB7AlmNecsXxxI02
f3Pzn/cmNu+bcLv1I/uoIUpsD5BEUt5ZjRC8PovhPvqP80iSlRdHQd1v3PbAP366lx2nw9NTCNLd
pbSDihrdGnz9Y9AreizyjIEa3BUe7O4BY69d5emXoZ528GeRp7arL8TBHwKutsioOmTfvyYw1AVe
hx2/4W7X7jepZCx8taVmNV1ca7Or5a8Xz0RMUQFpWjz7xYZs6/RZj8tFsWFda0V8YCgkMAf2MCJ9
KeJGg0xYrJ+d2fQEl9JXcARJI3HZDgs9EIBPOR+wFunr+XZ6u+KBQiXfpTIWoAZxVRht9nV9ZExC
eZQYUZTRiF5TgXOKdi6v8ZZYmJh4pk+KJxAPxVNfJGr5u/ODoY7Nr4e1sTIeSomBze14b4quGXFy
dhHz5VsOSTPNLwO0zxVGAe84szZWGxEfVMeJ6AR2WFQ+eIEaLOUoURc3oiKnkt/ekQoA/hxMcbf/
6/8OED/Imih9b+HwbqxfWxHYcMGgW6NstHfKqbHTbAqRLaeQtuxPGsCSDupBds1ptTyzL8AfTnni
h7IZg66Kv6NJpTBTcjAKGfeBwl/JqqKt+Z5ab7GP0w3FDZMdyC9sX0UgL8kySGdaHkb4a8buVk2B
GYL+Cr8b/NJmyHK32H7gBWT3zR+BjxBbDpPDJUaWh4q6G+wF5xyYUAYzOKijV9S3oetHWVQXLuGA
NYRRVNuoipcrRj3hnlKxBRHVXU28p24AeDUIFG6INqLaeopn/ISUZ8+CEeHKMd1jy87J0g3SAMQZ
NWggNiTx3q80W+yhTvhBokC9P4e3CR95BpSiAu1GQOFMbS5DK5XE81oxV232NVyPemy62xV2Ui78
FesfuBUmFt6ZhcmMwjQq2S2hNqWQsN9ztpMwPjAcRt61KU6T2iYLH5RqRK2EeFTgDRGTLqWdbMWo
F8IT9B07LrJbbAPnThehRY6qXUywvv/BFbH/hhgtNFm5f44xx117GRhHUXneHSvB2IEhP/vDVJoo
gVn14pW+3oAaxYCgsm9ajFkdULb/RpwSq3GjzZAd/nDhn/a7sz17+NvbGc0yW+0wg7RfcLq63J/s
0LpwnTu27G2MaBz0mSxejAL0CW6L+YzCMv2pGZjxY2w0bsEWMRYPVFpLA8nkJOf0z5taSyi26nqd
RXYtH7qqsvEHM05uSU6nSdFsHWkzz0ky9BpMwWeDauna6gaxtpJwaMDEHieX38LoPmqvrPUgcEmw
xvzPz4jFjmZSpXlGu62ERkbxyTBVh8FRMNUFV7K362WXQ6GHr27guN5tJ/NIGngErHbhBpq5dL2b
aH+I2NzT0dZE9VdNyozWZxIyeWc+JSAteJE9bxbOygKtRhGTl4t5rUgYxitmBDO2Of8J2uJh9NOS
4WcrzWC8ExMQlJPWxvcfHg4LsmqMSvx78UOrHHUJativNOYDBg9p94uJfVB9wzL7w4Jv1/0PqqaU
1Urf89Pjsq7zDbucMIgRStgmsv/PrXCbwPaFEwcXMKCajFSGIHpM/mH0+h0FqtfZIEvQD03QBnOd
evBlBWJjyYRVaDguBoQpKQJN72U485oHpMl/laNKlQqN+7x6BY4l+XvLa/gg9GgiwNgGU3y7MeCl
IxGtO+grA77BJ7qC0+hQ8B8E3lEtyM/6B07Vy88sXi6cqYMyZNX7TyUE2Ev6ztcnazIPWu/YNs46
f/da/n3FxJfPHliRVGtgqQiSqn1faWK69QtVIe1d2mPYPa2Weqs1FqGHzKIrBMc5doCt/HH81R1t
kdmokrWZLC7fUC3moA+VHAAvpH6IC2c+6sA4MtyULDdYAOesSoVlp7J8XEvgCDOhGCZOyLLHmquD
N/lJWGW22X1DmpvxUb7i/D3DOcIOcssu3ATkUuQ+pxxbib7ZNJy786C0hWBa2rFU9baucRjw/+rQ
jOFHJOU5qF1GXnuxZ+HbFM93xi+UO22wEQ2bzhBbOCm0KEVQCeZHaqGafeyiL6XsNKPyhPMXA3J2
eucfB7orn0N48ptSJMXa+GQ8vYxxMvqu8kPDK6T6Fviqv/2IzDnFaXbpiO20dhnclGL1XhFoxPPP
BuasMd5z9DFsRBsyeYq/xi38wHlig1mPW7gjYuvkX/yocYBN+sUbpk1tJIFh03GZV9eywDnQ029C
RUui/4ePs35M2L1LMAkEA1B5l75YToi+puDYgiS8ufucfyBGQlr2SXyfG65hzYBB4rFvQN2cxblH
znaJf+Z91c3xkC1St4c50IXNVqjgSRIFtuS0xW/uwNIhbVTywMVOULEam8KtMOSwuyqz8S7LhM2e
LOsRhJANyVLwVtBn0wTxyI7wgBK/H5gAv/l6VYO+b+ycln460ev54jtbfQHZfhl8U1Bx0ko1ygf1
4d9sHAQzhEddl7G71KaghSYObSKM+y911I9hw5RF8jdmWpRx9lB9riaxbv9U71uJlqUoNoj9GF5T
J/1CwqpdTq+buZAJf9A1SPMbpIkokZhl3GJ4xJhoX1z6ukUGi+3vMZBw3iONN4wgDUO1hQR7wl+s
34fzy7sADr2kFn+ihFIuJ6YstsCGhYjLECvElSA1NLODo9a7i0uUDv1JZNyrdGPTo/Z7UoqVk4ks
5bDirqZt/Mxz48pkSQQKBM2nhP8Tj+XINbMbMcbCHz1HJBidiAvi/42s8+l4BQFwfVPmZ0bvP3pw
/+IyihiB82cEQcRfFVr9GtJa+/clQpWehE2626/Vud3wToAO+H57b3K1SZRGwYVCW0lfTQcdOpiK
u/lsRJalCy6sdsheIQgGTZne8CfuI8N9N/bIdYVt7VpGwA8uJgKeDkHQDJFcnIX/m2nAL3+/Y22w
yeuNk6VrdYhT54nG9BLMwMX1Pu0CtdFBkHvFSKC/qyGonBQjHl8Ercmjf13gJDe35mjHkyUnPkFM
NT3XxWCw7YoHrIWKEIw9mh9XFQevFVTSyf9ihw3qdYN4qQuqiGGvFzYG6wIKJ+g6mtQBQF+tnEuN
NA5AwVWEfAb0k7EcXoXk4OWCwRFTs75PiOi6BrfZlmPe+eWU2JtwiRejwL4aQhA1bqGGSC/nlflZ
YudAuoL5qT+UNT9PlrAbgPkw6Gv2vS4YX0f+v5D0cyGSmXkUeqnubL098CZsMyewA3lM6OSQR/1x
1xa/BUc9/jQKi0hbgrnYhcrAgrzuxcoh+vTM2BBr5fhygBZweO2GJPm+HT+/LsqDpURYE6rDLcYx
IvzJg9xOmNg+w7CZjJETYCAbJSQaDIhFwAZHRq02UXoqZOpSSBnuy3yXuqYXLjyb1hGn0s0Mp0uS
QpwTkRKSlqyOBKw5xHEiCVv1E//jxT1kaKD9++uHc7V9aTSDi8Q/+BulPz6JVs8L4gZihZ9dgY7Q
nJ7NJH/al/3okxhcAtAX4s94RBVOH6soleNWw+mCGgi1kr3ik+4+zuqJRoyd1g+bwAMtyXU7adSE
68ut6z+QYI+gLLYuX2o1k1jeFLgSEjAliXUgNpOGaTfeJnI4T+MSFSdgZOBVR+JaeOHwDOEoOb1u
c5bATSrIWzXmtD4xIXGaP52grCk5m8VrHjcPsiVnclJS+sNC62n2FLFC6JcALbur1Z0O95lZXsyU
0QoFsQ4J9ssG+dy4058v1xVr3cm3X7tIm2gn/Rij5HxNlv+UvKgEBfNvkeWiNMD13q4LZGwu2FxK
eWqP39kzckpxMrnS0IgDe0iZ+GKNZ3xA0PCeP4ioZDtEToq1aq1dKdiTe+UNS9CPpR2P9jZG5k+j
VrjoLr7w7IJ1Stw16OGsZseYO2XDdhliO3dVNzeiF3zEMY6cQXb5tKUeoDLEkDQdUWYlhyvDNZYO
LiS5rKAM14jDmd2tUZcn6vs52JbkjHFxTZLr8NzfEiUaFJuKgpkvDbdVqEkSsUE0UXQETw3nYPuB
OoXrmp4cFVGd4sc39MMLZIGAGqbAKGKfr3EcluYjS5xlutaf6r71AC9FUSPt9VcVJsFHnHbS05zs
hUETsyFvtxMWApWh0R6yVHM6/CJuC+PRSNuX00AaALMAVW7abd37wB4raQP2+YgIXDI3UTXSXCyJ
zTvQyiF9WDr08D0K/HjhhJgHE0FSK8ksnqfltEmZ93SPQTqshroptp0PeDSYlKQdouhhU+Itv6pI
JqkLWL4vq3rfafKwqj3udUEKmQxHEHqg2LToRDiN2j+Kq52CoILg6NSobjp/upkIlVkaAWcp67VK
xAvtIASjRuilYRphLievTofWIe/0vU8e3qxR02aschwXba/qca+oHiPRbaNn05zMNN7hDpWnjsT/
sgMM3x3TDhdyyXt29kgtuRSvsNA8C0jYlwIiMoXaJn/KPhBMni+L0pupdDB84Z8qE9jIYjIxHzOG
GfLLNnatG0haHQhVXks+PcATVjh/+iohhJipyEQwQlSktTuQYQxjLmU7p6MbofjFXuWXZioWPXQo
TWjtd52APYT1dz/kwDY+0WtlAdPlWeGLYot5yPogiAHukDoya/24M6aO12bM9cpzQfcaTC31v0U2
I3DV4xyOM36yUf5DQiR7UJAMhRUU4Z8OTJL6O8Yf2dUK/Iz7DetmEAlOJfKunSnXFYd5AfQFc61i
m/dfE+Ec4j6pZdqFXgtFC06VQ2PhX54h07UXkChgEujpGaTuPT9C7o1eomX8r1eot5FyLie9QStV
NqLUa9J+Bw1rTZXf54K2XVdSYK+TOuflSg5w1xz6cHatbCrILvHM4KTnP1LL43IgUz6EqP1UxmlO
ZMQsVvhMYdw3I8GNXk1hOxDTxnODsU9Pvc5smq9OkW5TEopyhz1YZa1fK55gKV9826pJBQTirdBk
WsHCOznVH5faV0w1/pSy3opcHt7WMmIaAMTwWUGKK4MD2TYL7JFZ9JkcBgO/Xq9G1nOnMDZVr/mb
was1o1u1mo08Cfiigx72nMbD7TGYhxmmtEtJTKvG29maB0TY5yMgy4vy2/KrmW8g3EkOgrF7R7CI
vH2zAAJaKXhE0aPJlYHQch+fsQA0WrJht2w58M6aY6eCeSn+vwb70A4mzkKLXTk7I2QQaCwq64t4
z1K0RtcJcn71t5BfQ7KeOksiL4qQmqlwpfk07wUVT8p2sE/ds577E2XpTXKa7iviwPiuUBAeeW6E
NUOCdefdsZhebPHhYZUtgvVsMRusKVmyojdUHwZnWciUp0dFgP2CwTBTpXrZ9r8Tj5jLtEZ5jjtH
0RwMulD+kBH2eCPnmgkCu3FROdbB813SpdlqnpUwtnsabDoyKbM2XXfQgYsBqE38bNJcx3v3La0y
f5UxCFHY2guCTjJSzxoZdml+G/Y5BpIdygc3ZjaOW78E24TE47EASv4xtf//bAnxdyUzQ0hOO/dG
9M7vXTM2LDKLfw+HbIKtwVVwXrfvpA0836S9nVjVisCGJ+KA6/Ik8pq70gyrQMoRnF2C2JSpc3MO
/5fJRzcL3X6S7DUTunF8XXOu0AvDmbOXE0IOMZPY4xPT4XkI/OAa7DTCsTmc2KCyeSCsiaWp4J/X
1mZYRKI5NaaWuyoeql5P6NHrVlEQNoJlTOEtil/BVymm4RA/3HQTlpKn99CPpDM0dv9uVgtoomMD
fbRqhe2io/cc0ekPjgsjwSuOH98sZw2UPrnqx0W6138EAYHmd4vQsWbypjntaexMlHfVvCOTQJQV
kG7G/3Mucdt2HMYQWiIp08237Ert8qhXOXwx6mW8i1qUYjwyxxnwxJUxzHG0/knViGRQS+vwW8lG
cBczB9P1JtD4aLBjU5UO2R1p0ok88ZexqwNH8Omk2UMnXD6Sr53zLgXjWjX45I7wHdW+blO5KuGx
ljJxxa+fCRq3j9sJNVbs1gjNOP0CIxqkFsEJg8GDgVcOb3GogMb+3sztPiaXir8uvnNwrVMdb7G9
lzXZIvlBEyFamycQ9VhnR1Wm0RTBviKOs4G+roXloftHWoiMpBpfDAGOQHgvbmOdBgUcbbTQ7yes
bNi+0PfyDuUMMlLlVYPzipxq3+jjU9yXSTv07AK5cea2X4Jh/ZUzPLDDMy+2vXmnsW7+2VDRTYz1
dDY9m+hfQQrcHvl1lJ5W7ZQBTIC8wzHdjir/KkrJWTfbY3fPGQKCXEdbVn9pd+Kfyk4sbTorbCvr
EuLRWekWgKE0hY0zl7Y1s1ju3Bz5h++Hef7VJj92YfOlTHbClyWzH7dLD+lbQ7hBunTYViMr1o3D
dArZ0cynmJ74pACUgaApIVmOksi98jLUE+WXPwTOCqfTcahIZNCeXjWUiJGoTqxChVTbzNA6RWV+
rJ7ER81AlJiw456L8/plOynMHKUNBJ17HT2Mp2MdiFQvtttkj3T2tUxp785+E87qjYFQvSYLDlza
4dLq4R9MgXuXI8jAYVsy/MmmRB0L5sHo7bWi/m7Kr3UIYbqDD5i0q2cw0xHGEDg8YfVukcmqFfsc
18//Onp33ZStZLKWpCi6xKdqxe9qV4jMpwt2zWqMvajPdiZfzHN8S27Lr6LiSWTWp4ftsERQJJlW
F5NTnRbS4ukmS09OEO1vi5Jb4BgwIoSubPy7UDiPZiG2uzu0ZsIyoiHit59qiNf/zeq7DADIZQEg
IxnltrjFMzkaiig1ZRjlPffGtFx0uuS5ScBe5carA2FxQ1oYblYg5L3rVjM4g5TRrnkvI6C9owmz
jiC352paYGJxRix2Wc95+WaqeQWDzi230nrzwPZcQZJDYIyUyGKlnhshVhBSpl5eJUEQwXXz4lvv
lQFbbOHxwKah4/oih0KKQDfBSJx3ydkndsUSpr6g0x54oZzFednfZxlVLUOqvLCyvHJ78KlHAyC/
SsjHtfS7qCADMiCq9JQtl6Yo2T+Z0YQ1qfRFHRTvx7KPsHasP7f/yemuePwbx9Cl6+g1u+X+xrgQ
IVVax/a1zbE3xzGJcz7ETujy974mRLaorW0fGdr3tIbaH8NdC95TX1prYt/Og6fSyDMd3u7o3sue
+j6RZAiif8eLQNg2JYhhM+p041lsv2Q/i5z7bwWjHpOLJ20x2ibf0gEk8C3utmSniXKQ7NcKt2FZ
qApQlhGHf+qZWRg0Jbh5FYuUOGeUGoTezYCfIEm/QAzOdbBpIhGyNpOn918zpJY8OQ65OsldBgbq
wzzHvB78effFqDK4bSAhHdGRWy5ZlgDwg/Mu7JT/wFpGAylpuS+Ir2DRmaTVULj4+oOl4HKugAWH
KV1r8kHQPBkJZI7PPDeofw0cRLSyunXK7GCKffHPN+5GAF96fzAx5XP30yiO6jwSnORlwXHWIhtj
vlkLvR4Mmt9zB5seoUuVMI5U/umGthDDJ2oDxAevNSmiuRFXWojmvJaVFSSJKsaAu6X/B9zg9+7K
gfkbrl/kDRdR5HTfPryInfUqr/t7O9fS9z8jqMRrVR+2k+xpk1ujQEymX4ZBWtkOi6wZM7IHgrfj
zuazBEpktA1qsxeF/tXqxWMOYctBEWhxZZQFtzDJiGzYCRynAGInrBv5g01/tUzFeKbonrkrYjzr
/m/PaojbU1KF/vobNS+Dcv/yEwJmXt4+4d+nZPKGF2QaP5aVGbyGNjCgV4CiC/9cOIsHio7vPfwK
CXSYN4UDd4546VwKP41Ukl5T8U7Onpv00H0nTNWIKs3un11HOz4c/1iVYp6Qwhdf5kX8i7lXRVNn
D196QtHIryS1jCiwIdmcaOEcKf4frqhJ7/9TlV/iFfsKYTfyEKviXhVyfa9/MZhnC+d9Qco71oZy
foC9yyS2Kl21LcTHy3bPUFCs5zZqlwlPhnwIk61T+X6QgGeOl/FlYPRiZRHHIHsXennVDMTopwaV
sTFB//uSCDecyjJBavcYquDpqjSnphCEDxaUIFH+tIoxsqC1c1AbHUByTfR136lOiEBfgUqepxvn
H0MGsw+Igkk/4uAqUju8QskhJAekAYPSljXvyaicu362biVEO5ulq1Wpg38+8tP+XGljFHyX3GIY
FvyBdQp3OhqnGFv2H9VPpwXgB4O9GH/reeq3K11XeRtzBpCF8RkLD8MljSWid1buoRDs90E/YVAT
RMu/9GICDwHGSGdB+osm14H34lvVN4L1xfnju8TVf7y7fu/SQynqkhOd3pHO+oG7E2zLsYxHIPUD
t7BWyCHTqLHaAJAnvm/dAkvg/C08Uoza16WZJJYB/ymJJCpZzxQ0l3e+v0A1qjx6Xyw2eQUBPcG5
3lYefakX/I999NXlGmizZGNwb5ZSnrXjd2kTzadzK2CKekAIF7Z2RA3ZSwerqqisJghlqbLp3/vK
WswxfMfKufC+KfIz6pBypwb9XjRW2B/2eU1Y38Oi/kyEAbxiNqNYjhvyBebVT1t9eGyjaeEW85kr
eq1nBJcW1ofjFL3+wvMPI/ux4leuN5iYStGUjQDvKc92dtaIeAcQprCkruK4H+JIkXBVmyl/H0K1
Ne/kFPllLrepIV4EHnl3FbNAYlnAlq34y4Py/7f7b6P1d4QhjnXSXKSMC2tMGwO/XJV7WpEeCKB6
8pT9+ZJ9eZM8mZm18L1Pxi9N/9iFVGT6AVJxJR6WJAAXzpZBoXzxVYdDwxbpnOpglbrvBos8WusX
ckXMOFYOCAyhEgJDRFR5VT9WUF6Ld1Ur08XZvlsG8FQ98mo/D55iCEJAX3eMxsS1rMiFuNf1NMtc
MceuI8+Ob0dvFFtl44HFGu4TudQyqZQRiwF4L0kpVkql/vlhdOJEUn171ikVF4P582ao+f6nN5pA
/H3vqJlJ5RYCcXgx/4uZXHAvi5ONB5/hfyt84GcspQ8YLlT5nFbf6hpoV3p3f6+IiQj7zasuaF31
LRq+CC3zcL9eyornBefyO6kJsIN6dkqqAN78h3ukNV2gRSzsBvCjS+SvxWKsG5Tnhm24+ldAh9uZ
wwPVYdRDzRLf+VANGUY5+NwJyJ23rfziE5U9JsNRN53SJqyDdsGfXADoc2wd8PwhXnlukT47+IS+
Jp8PNl4CO0j1gvHqxFXU9L5y0PIBKLKWFthve7RtQga+AQkeCujK9ARD/tTXjzqtM4MlhbYptnDC
Mxuj6oSgVG4qHJcibZu2F2QtiL5ZGOw+SQrHMA+8/9osMCwmWtWMMHYioevvYyLW1SMDpftdwVpz
KTQcSy6SWCFDBha9iHby4o1RVQZ1vWK9swjjAz7mCQkpGQ5bxz2a4szsSCzR5GPGNrAjU5qWzlZg
oQPh5B7bSBIV9z6iT98imkRZKogYvxUyTOpYyRMrPnTdtbx2Q2LbN46OvChIYxozEPM/JxhnzXae
lO3PgwDWYi3ncv8rJdKypW7zpPiou1VG55+V8GuBe7YUcEcQqGOtHu7kyNKk8hjioJ4/1CDWp84E
LzwYPIq7lVQ0QZ0w85/8ClamPq+3rksRaX6c1D/w3dfpk3VGF7rrDxlakH8tHMForjcBfIlEClUD
9deB5/FL4rJa40Gxi+WFK/9Ir5xKeyj4EUBOfNdfZWqdgjwieVMlMav0N5CbLeROyqKLohIaNCHZ
Lgql17T7SrSVx7DyBcsOWwRXA8vfR9ErGymQLfz51OKMmvm4fdWAWmbcH7K/tFvUZZYNqNGu0EGu
Ybav/AvGv70pTl7myfnL+l19OQfN1x0jOE6KooafxbICMPZ3Xphet+lo3DLC/gvxGAPoXOpJyjmK
3AtHy+Q5bj6Y91/z93zfEFSRfGTL97Jas1E8C6b8s45IZP8DxFDuVGCDSHIHH1WomncrOxbcsRMD
Go5PUpdvtOEOeyLrFbEmEI7RrcfTUoEDaOt2EYtPXAzk6di4rxhPClE3LZLZPWy0N4nvzRtMgJJ6
I/uumNRB4+Is9UDSb1aB1+P8ukUNuTEagDZOFO1K82V2jVXjdhvhoSvRhiUfPXj/dhHH+dZXBW91
RwJAZSgL2+1ywvywqof7VUMo5VFf45dYUo98JrJwewEfn42avad7n6N+lmA/VjeE2v0Ua7jMEDcN
s8Ih62vqf35n9whcDKDYlkRZUao/P6vYC2ISWNFvRVpfL++sCxI2hCtimL1WNoDQ0wpZHlokLd95
nseJNazVW0tb7RlGViNcpzIp08SStTSEovV1Llnt08N0h0sMiaS6C/vnRa/AUKGGXHrYeqoOjDj9
Y5M9Fa71nZhPgF3BJn71fOMdmQoSx4AlxqwjgRcMIczfmGI+E3qXC6nstuLnDeU229b7rPZ1AYZk
ujmACbfUmZQ+Ci3TnbHVLJhXEOlEl9/uv8C7S5l7loMGCrcfuh4DUAEromsVEXpiODfifYEZTghd
D9Ae/XuU6JFRnvKmg9MWPH9O5/qn6YLZ4bRS1qmpVHIA6utFnhUW93E1FPJAHlUETEYgkUui1xuK
mfR57tUTklDGwnLqnCbEL3qj7QybMGGW1vh5I3YkZWV5zKKcm3VPS6lY0A+poJC4xqbQ1zJGhhcw
K2Gycj0BDwo05wFT3j6euXMjt/lMSZ72XJ/k4Boltx96lG1nHdTYyAWBjvcTdgG0CDWnfP0SXerj
u31PPmzgU9RLYno6ELeF3a6ouQGCl2WNlVk0nrdrNpN/3h42Aym/WRaF8GCUfvVcjwfN7LXlT/lF
U/rb87HLEL8UkWn+49MlrwJl1d4HiX8h946aL6vNXYYZXm6+KgNzbaup5ZRDPXHai09MPXJls8aa
1zgcncue9RRhEnjz3Xd12EjRxHenFNKNuqnSVXyIP8zssaO5mLYeA8HSWVbcHk+6AA95c9WM+xLT
4284NdKMCHDMHerLvFZUMsgyQ1ybXyfPqWJQ8sTicpq/kKgp0Kt8ATOkuj3Ank8MM82D4EC6TTdX
6odvsNLpsTpoakYUYm+bgjOywoAhyDh3626NykSdl1eunWJDX8ztxBXhhqPIzDdp8EVjooL0xtw6
mlbpm309uQtIQRufeSIPutY6YjrCGNUMGMapa/4EpQ0smZfeArl9q1rd++vdyUSCjP15C+kGTvoI
+bVQY45Lv7yoA23xqQxS8J8bNfgYkXAIplPTwLe+OczllTnvrVGQ04wOO/69pgB5WgTgDMycm+re
lyH5HT6CXPWN83PpvZULxB6TutQev02Ed476LRIN6nsPgFx3TWSx/1sI6AP+rlj8trXOuqntM4K7
6NyL6E9zEm3n8+2VzT7XMNjEhYl2pLlm3SfbgJpKJJckyf20zYxNoD/QkFmOFvRXHdDZ2Hp2Pumj
GWPPBcD7eZD4rqxQyGWWnYpKmUfhMNIOIddxxHNWoWcQIGeTXZwCN3iC8g0fA+Q1qMEeUyI9lSA2
gAXOLLlWUUQ102fo//9DchQcuuIesJKALLWToO3Z4B2LYEl+06k/uPYEQl+Tl9QTQ2QL7wt55UbS
kglNavtedstnlFYIvX9PYn88MfygHFrarch3+poBwn8nD5yWBRFMDBrywNVBoQoBxy/8ivbR7a30
t8QICzgj1D8Xal4t/dCh57ROZ4seqsnHVFlo/nMZpkPKGzR7y1Mwv/QCGc5lYGqeclqEQV15dfHN
Oo0yghcTK+BsHChZ+8WFHbcV5t8E1P+v3G7tb2mqfecQgqA6oH+4MvuwSGhN9OChkLuPdNFQcuLW
ZXTNo6Rj6cIgFobadJikscS8zUliTijKLVfzTvF6q25yy4Iac8fEzalSBCYwGBHxa1Z9/Bx/NBwq
YemLCW2g8hzXyYD/uFgC+2IWS0eiDui1+3K/mMjcRrnXRLzZmHB0jlj20mOUh04pg0iIBRZ+7sS+
tY37QfG9jYMKPxQ6bLKlQzRjfxxL9CsxOEl1mdhT3203JIs6NJfJbbZivbBXyfqp/6XRK3I9U4P+
iEqZhHniTomUiC6NL4dqO6nAcjRkRRnmhe5astM5ixwDNt8pR/GwLlJJO0yxYY7zpJraDaJj0Np7
NmjiheL4Sve05H1pBWsLLK+EetbIsdABOuHfDmG9YrVRlEGvPJa43YJ0deqQXEzVJziOQd9lIjgN
28vbcHb8n+guXagfl8kJTC1RNp8AFPKVByFV0iUgSHNHLWORrTY1ViO6io+04/YkGnvywjev1TzS
KRIh8KZGb4HSkp6o56jjjYN4ypaIId857qtAj7PXlD+YZGMOYCEFcnsiVSalnvfMHiambdrjFrxB
4mc3x+XegHQixysRGBH8nRCgkv+nxtUGQXCNvpNHrEP7Wp2V37/v3ZPNVk5TaVdTM24NdWBVZuTy
ydCukWywS0DmNykglMVJ4357DDfzFkLaDsfA/s+gUOpr0pd+RYufz20yfySETyp4YqlFKbL7gnVE
PO09rq6zU7bHFPmnF6YaEa7GgxbVGbcUzgs3LzDxc1mImPkj2apVZpXH3mSlUor8oB0S3SfCStWW
9Y4eWR6CZ1XRVU5/pIlxY5sd6zkVZ9TYbmnYwkTNcYVdHXBZDhFV/UJyi71FZP/3uBZZp3JXowzc
ll+YrLlUgipjT6sNfvBkwE8xh+AXLioOQaSD7P78pRW6TLxKMtbeTZM540tkV4EqMM23Yg63zJTz
MajIdNamRpUn2hemYdxOeJQJD9nK475kXaB4Jivv0iZUBlqPgwHEtB5yzAl359l2Bf+DOBM9R2T7
Skd5Y4kYJJbSNGap1NyEG4L/H/OFvovKKq7gFVx623RcLvFoKnZKefdDMr4PE60SVpe0J734ecz8
BZXkhfOoA2SiMrcGKqkA+2K8C6IraTkqJ3CJ5KL/9mma8owE5Zn3PWbFzAWAtthEchCJsEJ1EpyK
RuxdrfAWAbF+STp3B5uKeMv98qmlEe/6lBuijIZHfJXEuftgW07A4Ma2aoPQGAFjuBa1Bu42GSvK
XYgdHRJANn00oDfxIn3XrEi+jb/i/tv3WRhiKFYIMdl43u6Ztd5lStT8vMPVghZLzctuxFfLwbgS
1UZw8PTeTHrdS3zucUSCiV429+cITzwFCd9xW6UY+eaTaoK8+7jRZXm5MjfGfL47WLXlYvKC5yjn
tIgssa5ZV70luoluPhSeoh60pDu8+DNTpDqeg/6ipHwHtQfMy5XdX53nqcA9SQaaM5Uzm6V3ndrb
9kHZlB/48oQiF9X3XwhaGit6ivlZRvpKMpBvBRScu1T5QfQrD6K39AuO8/4zJ2dGAdMWLmy3Dlj9
hK0RoP/QgIVALBF3ScWcFtNh9zdwWck/9TXTXY2zfWFgHFmseuYwBkmFU93cRyRmdNvaaGVOcq0X
kabiqcekctLGuesiRCWYsNIOUca3bCcQjFXYtv89t2ocDcWzV0fcEXoOz0KZKAW8DLCyqZrfB6hF
aCQwhjsMcu2TXijugu5SYqC+DpFsLZWoSFE+PfigmnK95tpjfPRiuvvqWt7/D3GpdmW/wj/1ytTK
eJj7Ffa58mlMW5MxolCDuHaJXxjFHFbclg+ypkfSwVXBE7Z0wHiSa++DQGSpsTn5an7C+ByUDbrJ
gzBtpQKEkKqmb9ZFHgxyr1RLKUwbp7JHBJWIiA04x84J04RHMVxQG9kTeQdOqPN5HZdvRn6TQdY6
vZ6Q771fszkJxxNa5BVCi6T8osnvBxOOx0JHewWLqlnR28l1vplLi7B6zdW4EgSp82L135fzpc7h
7VGak42hOVChxAi8PzKv2X67k0IBWPFfT/B7ZEY+aC3mnkacM+74jbVAXCNklce5csvDrOVwch1U
ra0PIeztDR4uxODGQvDijbNRaHe6WYSEyp9K6IY9hFBuvRSITpA81BPyAtuJy6Fj45DCN+L7vV1H
ut7V0EIaXFXfCBDaklMup0p0BOZAp2Z5qiPzOrDmtaekaCAwoSfo2HKfdu+jXNuDsuFrqJ0W4R+u
Y6hqiQlMtbjxcUB8+3B5WLV7/GvlvdZ+8p2BExWdb9cpS+/7VTq0zUwJ5q0DICDuPocGXyB8pYQw
E87lcF5ZXR3V1JrhXGYVQVTN/YyAttBVjHZGojD0K2AvDCD30jPM1x8lue/mKv1+WRIXxvEHO6x/
R3K3Tv1dKGFQZ8+D1pwRdp8ffMqzYKo0InLyHpxdmKvEilXB1lg2Zf3eALryv/JtmvXbVknHrwZb
mIdRDTwhbRpjnjbPgNxnE9AxWPrJ9OjoACwQnZTD33+XanQEl2utHPwOZE3wRlNYJImla3odlfvr
V+wq+s+Bk+SctPxe6Qt8N2XmFBo24nPffzhx7lgFSw906t9IFNm1sAo6eqY8AHl8GSyN+wgtLbTi
29T2ON6Rp2uRzNzPjK4bydxrhP+ptSD6oG8toEqvXTAuZiRmfzpAgHXYUXvE2Ad+9NDjAHxjJ/Sq
ol38ZvCDIAmVUyBrwkvGmGkpn76UH8VgtRb6RqbIzq6M512qUkTrgDkkfGB3taXogWdDx1G1He4S
IzoNPzCxsmXEAMupp46C3oP0WWVXDOZG8QueIiKOk6YpL0ljZMZ3qNqx8ZoDyBI9+eZ9/zR4hzXC
H75qa3DgsNaYgebebKtfbxQ2MwMk0FQYBFwK+9UAVESnLzY+YeM9VijwsrzDFQt2aTHVc+kQMLDT
ZInNFwV7mIhjJzeUhL1GgeB/RbZ4KcJkUAc/y2o6DUpgLVA2Utfo7c19xXh2LTcRYkOwNwih3J+Z
HBRMOPlU+DZrOGqrxs+0aNAxO0mP/2EJXJhobCTbSKtQ3dvfC+2LLmu/JRV7H4BbmCOe25mhOpEJ
XGWJxOnzBLWkocHlqrSHQmCDwFEtDixf2je52eZ+a+vjnHEEr2ODAu0kWcw3gEtqsOIEJoW6L4S6
DA2SHgSh0ERxkTDbfHEcaOpHUePIbYdExSpZl8Mj41dKBLqNb9lL2K9ZvT+UUnMKFvhWwDhuwouS
HLkF2PPjOKkxGihM8EuSFYpIQaAw+RP2Ohcn0K11NSZu9nuxyApkyQK5C/oytW82fOs1Ptk+edQY
mCg1f39sBf6nUmz4QrWcK6+g2G/F4OD7z9n4e3++CnD2f6eSs9aMBpldobQ70jOFmG2tB9THT1tW
4oXiQ1+0kXm1L5UM+eY8aQanN6uWn8WZKfIRIjPmjAygmgl30zY16Scv3bzg5N/k6zcu8diSWRql
i+kZY1jU5y4JFfVXl27SdWaKAtUuTWQGh5MfGOY7A+qnppbmBoLyeQMNg76KYkOxpdu4PUmtLMiy
+f/u922pHZzSnTkWw5VY0/MoDSjrWc23dk4UGDhwysPnbBmHxOmpu+vIT9hFHUj5n381c7gZAdsI
giWE3I0mWqXDFTxdQQTiJC1efrnTtOpVU9K9Jo5xuCQ3G9trOHH4Jms0TJBx08qqrtCkU/TP4wxW
ZNF4QC5C6KbDv6LeikFAqYs4qOT301tEjPjobsl5dHmelMKKQnN/bkvTGycuFiPr+c6cU2jqyLZB
z1NzZWDY+VcZ9TRX7uF5hPl39YqJ20BZQ5FWNvCSwly0ggR1WTp0xSy776cLRnM9gGFf+ou1f5P/
sdG/MJR8d+x7ksb8lcgDJyR22pD9oDE/umnIS8hUke3lIB3cxX323m4Nrz9hio1/psNGVj/oOCJB
ebHz+HccX/1ql6W1AJDcHCbjxiRyAHP4DM0tsvzSEvh9lnca7Qvt4oZvva3jmiAbZyZjxoZxrT6j
I0B8TNWydr1MJsPAxCABHqkn+QP7JImmfWHo9DI/kSSpuUbf4p0D86yfqeBTQKA9nHrI+QaL7ZVF
sDPXwotv6Qyys0PtnoCKdWRCQE469DZkMmA8Sls40ishWW+lVfpEWlOtfQiDEm3oWugMAvo636F5
cCQZgXdHnJlGZTqbLFHNMljFunyjRU0gQgja6vcBcGBjdmpt9g5tLsdCi6nC7TJxXHoDA5zICcQi
/MsKtOobtj+M1LIpphWcTUtCfjjVVSszXzHNt1ZdU657qijbs7/2aIxB0h1j4+tkb23mfOCkJq6w
d1wCiMG7ffTxwvvGDf9gpXOLKLJ8NAvMbP0Yyd3OXg4RoMnHUhOCFW+qcTny7Keq15dc+6hQDdlB
jgMcNJiDf7/F+g01jxvzF9WN5WF4Yr86P8HkIjAAtF7Nhzbf0QqLe/QhJvrSIRY4Tisej9bBypGe
wJkzvRrSYy0nmTupLxFj9nwoxmzkmfXR1rvel3bd4VquRCn2upJVhPA8s9Y/QDkL1UhDZ7wyAMWa
FCz+JBXrtm5P3UXTWEKku5K01X0o/aTzI/CHba/yPUgtJL+BCCN9dwkYh40kE7gGTTJ6YB7u5xmq
wpSLCFcJUJhEntCAHvW6OVgkfxv7zFaJghrwsZ/D79BisYlzosxkUIbeYRdUwQZZufyCYQxSMv0D
XDQkLMBdmykw+DE5XgARxd9CkOgLTYUSMass6in5+T9V5DuGewR88hd+6KZ9D7YbvXwlVlbG80G+
rxiHd73fnl8QqYSMxeXtcyj4PZowHcR0C1iT/8QNIf8A71TxGSlpSXXDLRnUXaEpCWOUs5bXZJ2p
X018TIRcN1IRV3A3G3wV09GraUFHJ2hPaHBP6W16HVnO/gFfMbig/SQB3m5k7ITh848QHc9SfrIB
KP6tgfyCf+ar4LR/uJhaN0XLXRV5BwhOyOm8w2AdQc9fpY3YK4ujFIU1zbbEwWX59iiq5QMVj5ZX
emxgQ+gx4Tbv+qfUvdJ1m9TRgo4knXlil8psDxc7fMbH/UNZr4Dk+QC/WcOpixtruK1vkJcgptIc
+aCGHlKAPcoc2imXt+OHWZ+tTD94ewPn+sx1N0F85+DOfxnafrzDGD/kRyYXG2hsxx4xRVP3g+TE
34A60uQDYkfakMN/3Xg6GQwo2Of4DFCJkgW4oSyYHTRi87VdQybwZ9q16fndDopcV4c2nNW8S3pk
6ZJqJT50P7Ks3XO+fx5S7/mKeXcKRL9czCG4Xm5YNu8mnX2jyt5G3SXjqeyHcwiNODPYOJNHHD6r
tSvROAq7/2kGbleCcCzlvXZdpEAYpMllJvScSlCtBJmvTH2bx2c1KtfKlPUZ3C8KT+MpwjACXY5d
04ZTmK8kYTo8DqH1XJfzZ3+pSnFlQJXXVFLKfRDJjLn982pPLfUVd6XwmQt+9pVnaEeHz0lxypYc
LHqS/xCYz2wgr4hA5KE6MDxdURGjcoddxXUHOIZNhlvZjsnu6QSuD6womkgdbeV+Tf732Zt5VRhD
8EOoa0Dj5iYGmRfg1Lgk7zVavYDYmWpBOWkh8CYNGvBcraEGTffV080WlBUAOPOsT/Gmk94DtDjg
wWiXuhN0dHVURX31pKOCMOUtOfPicG+ZiMO/CvLg2cyO6iaLoHBJ/u4xjUkflJsL05fHuREwYQRH
gSPOijZfLDV2NsGT5OZB0mIZgoafahCgBd1nru50MJxqyTjlvSR0GjNEzgBfalzUinbyLw8UiPVt
41Crrmz25VDyz6oC07F9TGga62tfIiMD22nlKEo6CdJWKmLBZY1sjLjoTMiQwERSswLVYEuLqXL8
tNu32dhppTjrTKVZEqTndfEp4YEi7fO5IgzWlPChLJVeYSg2OgUJWDFJ7lZ6epTnSFhseut850VG
GxFElDE2vMfbbL6m7Tsd9PgL9+WNaIV192z4sEKl6N5f75W44UAmD7l3D6hCsekX1EDBxZVxA4Ii
tde5cFv1tlkbRdZ7M4Jx8Vb8oOAigqQb1SYKY+5mFNB8dilDVzCK3BSSXCrNwkgKfYquMamnsdpJ
GjUGkj43TY7WTK7iiKaEGD3ylOc47nCDq7Qd8U1H1Ig/OsZZbk8ggpA18Lwg/yXV59hgxnFLgC1E
u8/gsttRYbGUZcU5T9whbSrvukmCts7mLE4q8Ec+3a1HS6O1zPQCINkxfuQxwOD2qpo8vKW51M3y
2Ss94jwggREw+d0BU4US/0m/2StbPuAlEo5t/WVhIm1jT8lNH5aEhdyfXy1+wQeg59ZwDLAv07PR
/9LGQ/GPIFqQqYSJfU+sQvGkcSqR9PiISD1KFrFlppAkDR4lkdvSPrvhDICEcU1Frl8H7XwfEYeW
oHAsoxeyBniTPFCC5ZimNUimFujGYWUk1kKqis90soRIpwMaGYT8Fdw5oxFg+5ygpWKl4JqCyg1n
ypsiAGaLRxtXvHm5mgw/+qi3319fymn7UmzdN2z41T6AXJsYueM0bG2zCniEUGJEKH8KWdAxP7+e
EO9AiWme+Vggkxc85cClilLwkeZOtszSD4OavWc5IL2S3MiagqkGarKseo7Y9KJmWqiRc3pQCrpH
+AsTsacOr31rqNZfxfgQdFtR/ByvaSP/98qWQtcAKhch4x5u55G9Xp6WtGOGnMwvY6faJqkD8OqS
zUqOdQmBJZlRU3vzkxBHB13o6XUOmsj4fdBGMRtSjftR2bNqSJp2MFMXeMR21zH8Wigdy/EZX4wA
RIpVtSRc35TVJ2I7GofchQRGgJ8gHUJPb3vSn0T2lpfQ0snC9485Y2UUJTsY/1gpy0GPYHj7+nH2
wD62TxN5fvfigd+aBoogYws9ziTlQxcTOLi1q6Az6WavQ1fYkNdhlOoCRtxuydFLHxFVbFphPO/5
MEYbfPwoNfKe437ROuNXxz7DeoMPpSXLusxWdmE70JfXABlCSx5e7G2gc3+Y2w5MhKPqD7LLNCS+
teVnpnBX9K4cygfOR490zXs0sT5ZVWKH/nmEzUhRdi4Tw7x/2KV9cmRuSI8WMJPpTsxTROlhhugN
OzA7KLG6s7y/iLvFRsA9GkSGOnZ+2ZahK2SjlGVANYFKSRfmchPBxJHADk6mi86JqqozO45ykgMy
8Wpa1OIQKRh3q+XPaQuZE/prKjV0ZFIIMB/fs2wndXLq4uAj/CYQdOFwBoNkdS0xgctNmV9V/FoQ
njtGf+By0CtUdnKPrMC6mnURKvkflJfFO11BAbqE0IrCpJaXDxVpHcY/2zx58QLKnUOUgerzY0oj
C490alEzmPx2sn+QiJSbXY/tiIGa2+CNJD0PEnLOr+lvBB55RG8Uo+zpdmNwZvlkB+cE/+Sj0Te6
T6HQOUXfDWteVQBc0qb+BLakkxegto7j22uULBObABheka9/KlnQUoTurWpNobZcuFRSgu7Riuw6
X9dr0KD2sohwAH/DSJukRRIGaNXY9O2cH4AN6X476Drc3pEXS+r700ULOJW0vYTeSYGbQK7EF/m1
vCLl97NOe1ONVeigUDUEmZDXza1TqHr1dauEypoxlOoRhvFSzffpE04g42GrEcHloN1mpGTM9N+L
pIVIkmiVNg85/5H1cSOkLGjRZW8N1vtsiODdEl7z8LsiEx+VIvzJq4gmEhdkPqdJ4X6XgBZMdtr2
u/1zSC3C6n/UDPVG7nfOW9BMBSd6BP6Az2UUZA4XNg+anMxELcPDph1ZmePu738I4XrDKgLObukA
PRGaEXIr5Nr2mLSSW3O54Pjtugt5U9thTTs+HqPBtDaYtKx0qSw8pGZUwRJLapFXz34CuGE+dcwM
LUe0bSNOoBrrYss+OjcVTp3VJ4ohva94ud+B/eUzWfxahs2ejMpFckU8SZK7+bxNS8ZqKVP8whUp
6qp214TJXgzZaR/+2JHVEHbAsP46nyWGgEsPiA+1mICxOWzCnURkZFVK05q28ZiBzKQLRRak+kx3
AZNEnexsvhoswQdhI9yjw4GhiKTLsIxMEnSlY1ybFBIs5XVZfI1MRurJnVRpmNbPg0imJ+KzEDSZ
SkvjtwOdH7apDpWS7xac6XhN0RJw6xD26mZvbJDnhqOfHdiSojANdkT+oqC5ISPPz/QSHg2KanHx
B+OxmMxdI0kqFyFfx0QDk+aF3UqpnOr7563Sk69EH5MbpaKygfYky/GcoC7IJ2u0brRPHudUr41C
2ZHlygY4QPIISMjMfAJj0W/PNlibJc1zCjJREN+BtCkTdy7v3Rq+CqMT0pmQry2RuP2vUkJcddxd
LaXlO5cp+aHySjbSZZ+lftMA4gLHEaGwWyNm8EPKZVFhXz/eTmbpHxnMSlT525dt5tF56s6v5jUC
tBIEPQKa8itnd9oVmKXe9yp043QOFrSLhQFUFFzTpiM/aGU6fD3BB4qwvOdmClovaAV0UjYz+ktn
LmEqI5e+O3r4sm+fWAkHqLF3QRtKTUbGkLos6KsAMi2FmMBnh8PgFQedWemZLC8l2yKjzaRg0D6a
pMirNj0IwXqwYg3Jb6J0PeV2dGgxNwxfT53OPAE1Hx05kvk3OiVfluQUjCkgpv1nouc3fw40K/nB
PdgLeEtq0tOfwq98fWG8P6NyNMj1CzOSmOrUEAY8ioO19p8ozT3CnTQ6r8qd/3Y3pUY1sWS1F4pF
o9ZhDZZp9YSAHt1gQjV/lqTgXYF9b9n/2fOz7tqclN8VGhHEXTg1qXsIz4jAf5UgPq+nJG2+6RA3
1wzz73ymL9M+XwSwWQUckAByAUdGmWdarijN21XSKu8rDEdrVIZeKxVc2LKfXVvtZJKl7PkyU/QB
aEpFSIqANDPiEQeXMuXhwE7EwH8JilpBk7skFRwyhHYmIu9S+Fm5QsAC/DpfgwH8DQUSTcbfqzuh
kXhM+hhH5sXbgZOCDw+oZXr2hWrt+thh03tydSTiQ7GKOFLdSxbz3CqJ94Z5ee93z4NchvXVI4fY
DJc5JLJM1M7mN4DrgH9O641ZhNyAwI9zlFVDKQeOSZs6L/pGpx1TBOB4mK9xdmJ1SiSGw+IhSxW0
h9kRvT4j5ln08izpcyyC6Ko+wbBDEdmvl6sJ7HT+cM2Zyd2MmOQd0QIDsPq3k3M4HKsggjDZoVOk
nvWptwvyccWeyn9FmUfFituz58spjHLxlms3KaJi2hHRSTtvbjRfQOiMukSUQSSsKFmbzH+YffV1
6Ky2I3ucy7Py8ICr+ph7UJ3f1DzQvHYZ3hxbvT/DMjfwQWDfHAhnR02wCl6w54br0CWT8VM/V5it
hhJaPaubN3aAe54J8yuOTpJcm29A7yRac4dCXVC8cCcweWCKLWwBkZbIOAzP6TmzDGOJaig7yjke
XJmMdwlDpVH3fCRpKEzF95ITybfVlH1/v3zCIkWkr3UPer0aKveInciwhgjM6TVTOoTQjBavPK9T
xcgXm3y4siNi1pPyYgvTMdmmJJCbevVmdx/nJuAxKE2RoLtBLQCPwRGNvKhODdtqnLtvRTdLpgkp
2XOM8fE6Fr6LbBt4AvnhElS8ovgIgaCB9YDFc2qrOSOlBYyrQPhxULBa5yoWnl16qfsMPEE25dG6
LHTTlYRYoEgxNTnIw+TufxNsaGyt3eaAZMOgt6/KHaNYRfY70u4dIR2btzOm97puwypKuvETdF5F
7h+FBCf4wOlYO2y65ci4QrdBSkNoDszQlc3OSLwYPQ+ZNpQAXDgI0NbUx52t0YUK6UDPlX4ZwTGS
7L4P09YF9ruqXkGK2ZxBavsBGaHGn9W8vEjmJRdJQ6we3Inl1S6o4fRuO2hkZTih3iLXkYhd/G7u
Ylm9iq/Rviyn+vitiZmhXUa91wRUEWPgzjH4C0pzKasmBbWwF+mpx3GFTssjnF/RJqyFSoyMA6GA
NgaTAT7REpkr1DcvIvUDAGWLVpXbgzh3VFW10iu9sSOZZ7VnQwaRvw9GGk2ldoXy1FOYBOVHp0cn
t+lvfpXVJUHYFdClDR5Y9waYUhH3vWINa5XCrt5K3ZBxaGY4KQS5hUHUEnUhTJBLFE9nHev8wfw+
MDBC0qCxdozQNSK5ZVBdCF9kekZZAwADKnjK/GYHxtfF1QliDil4YAMYaEg3/R55sUxasBHxxCWk
1Gpud3p7XKEa+4wHB/0QyxWFNkvWXfQwgRyh8S4hvHzp+snDJTXr04XDo3AnMPnBokgFqTtr3MXx
vlyMba1D6JZwkAF7kFWqBiGEnd0Cd+6/m9pYwlhm74wIPmYr9yYdu4CNrfgfQOtPrLXwHy9B3h7w
GPGLSpxxY/3TmV0b44XPAJZ1do+vlUvkiX2tfekRra4iVS7EeSBSnTw/6yucUKDx98ohvn0OgLzL
V3ToK4GwBmlXv9bX8XmZPyuPI8l6vEIxQTHXX9Rh7IclYj9GWFHCj0eFfOTFngFDCjsz12I7moCZ
OeQmNOhFtHO7qJL9p4e8oWjUAf1NAA5HzGuvaeS+2EBjSFuSIm7VB0d+eEEMxSVxbKBNwqP7XQ00
S/WFCHENwjdfni2w/RpyiLswGnkzqqshUpK0z2GGTNuzDWjSItmerPVsvRBRuHZKGMPZI/5zt2vZ
KOfXmxybi34LEP3npujXMoZ1h1ICLPkYf3egyx9h8gAFmC68jRzBNakbAW3pv8aWyOMrFAT8QhVa
JZQlBXAzhP6mHIaIptYwTcRm0wkKN8cd+RNW/aecDO83gBeJie6RAzais2UQACvfVpVyvj7QA4x2
ABh1s6jaUHDBycGDth0UkaMKspYRDlyHYD4looOklg/EZ+19DqUjeRFBJko8NtLah9PA1hb7uYNc
LO9WzjI35S96M940VJIC1uXJbY+waZSNaMlKXRlrdctLZqJL0Vn5Ruyc01D0cB7X3olv7pjNxNHe
H2Ra4HiyJP60KstY1Sss3G0te+HIaqFmEKfQq3Huuo3JdUvG2GBQVUAhYuQG+Nb2gi4cVVJ1CFWL
OdEU31dZ6zYo3M56GlyNrxfbpHQ38atDxV2yHyi+6gQBVfTS83juAuQZLNdCpDFd7awYQC6fIctd
rpz2svusBSOjKPn6W4g42q4UGN4TLBI3MtI576RSJzTCJFoZJY1OqOeuQ52Z30YbzUqBOoYLln5H
wefk6vFW3pZwLHEc2LDNF1XW0rjJsRDtZAaiz1ZdH3pRoSeNMWjEMeSc8R+ARYc9sQK81Taq1pXL
XS+/wjg3nmBD0FX/zui1qKR1REKsc2h7jdc6LV0i+Q0+BsdDr3Rvq2xjKmiXm5b1fzFobsWKXP9v
jlIhrr/ZExLQNP1CjL2vnQJ8bOS46sCF25L4S4tsge7rNO3Nsy3+MKCc706zNeQN/WMWktn+CB5P
3Uyf4lLD0ncEqgm2mXLEowqdt+D+bskGbfUp8u8ZQuvcSSP9nyHQKla7afAvNCNffxToS1y2iX11
ZmUd59nWp1EgDMb/HWmip9dHvKLhvaU9+TH3xi6RO3TRs4AGFOzvJ0PBBFesDa8jLYUhpY92m3KH
ijO1dHne1LB1BaIVdlEfStyG0e7OVgtSyzNzaoLJ4PPCrEIRlbJT3gVShg8T86prWSqx6EZL469D
S++HvF9NQ7XGdSfAGg1IIVdFY44Y4Fpva1MSs7Wt2He/ZWHFPad/EIO4HqMRfKnVaJMFUyHLqSqw
p+nQjvZqcGCpIZ6ivr4yCkIEdQySATfxUXiCOTxPUn47fy+8SyEdqAp51as0+ANcG/VADyyvhiEA
NP3u4Gl11fglvSHg78DIMP8xNL3CVCTdYakDqlHPtghirUYi4dB+yu7ZZY32bJ0YM0r/Mjc3HEYw
vAgSWwS/e2aOeMOWTu/iLghQZrj9uoQl03lNgFGqeiXab+dTodAfMDMxOwQpMoobqyxE0RW5g95j
Glz1X4j86kFMof6Wrng2aeMnbrTa1WpId7iQgGzT+fXZC+tyG0jwh1pzfAKy2kak7FpgemP/iwg4
Ra0CNTtDPfl6J9cM96FU25p4tA6KXq4Oe/Dclpgck15ejmOb/eYvsfpTkxxEPEGV5LvD3xzaw1cD
E+HcYXMyl5xQ2O9TdpFa9itenHjR1dabMU+E/ANPvghYBF6kiBlwR56IYq9bTus4mZwXbVDqpeKx
AeohEXB/PKKN0KohHuvOgkfYUHwN4Jeiae5/XNp+3raVzYpoZx5qLo0vtj2XQPUqTcPIkeYKLQRd
OTk0VqSLBdelbJ/z+zFZGD/XiDMWzoagZjir9wBr2IG+rK90rMXa4ge+qFK2aBiCclH6na3WMThs
amlhT8Zh0rcTSmOifksHaLvA4Z6SBo+CmUhUUFYkMsMzIY7a+5wOPuwnGm4eTjNscgjIkKNI38jW
AS9G+93PHBO5J01ala6f4jnfo8Oi5HS0Nw64IR7tYtUDoIiVCObDtaBkl92loeUWyYvYEQBfmQSj
KMHDOfmUTlDuvfqavWPQe08s70EkvLgQO49T9nnQYvgP5aXq83c0jFlSzILPHRnIapC3Y7uNLXuK
SJ3t3DGTc7LjIeDgapdJE33ngeJraxwta4jaVI5pbmH32Y+GcHa5rLpzew3mLxBp3nc5+MV2Xr7K
5TLzI6Qebu2tnWlAn2DCCtHwIndr+YQj+0Q3PDdUDaOwSb3KQuYPTRJCYagAFovSKtVqXGWnQC+e
uzZbcJRAWyOLL78MxDgumeApvKVunuwvzEJYZMZHL0CavU16iQUOoWAZivP2E3l/sSjzMJerRh55
uqRbaDldU4zi0+cyYhZh5CV+75ZPe8hMEywTi6PTpdgzDXaZTDHTgxT1hM9nNvIE5BJ8iZ+WdF/1
/n8m8C7qcKbgMlopoDH3mQptqfAZrkiR7HzlfduupBceb3Vx2BD2NpKZRif0pQhppGUBqSLckiiA
gAze39tmZnN0F/w7nrjV2xFaKaJWbMm1uCmuV6/JtKQjt1c3YC8Us9kMs0uD/UeYf2wxV2eozCuS
Fk2LxcJIvrbp+E0iI63ojYg2sj5/YUnyH6I+5xe29ZXbXuD76ugkI1PpMB0DMU8g1X8keB5kpCIy
SmAEdOhlH4CdpI+W/LbJ/CbqLqIt+AdyZvPlG/CiCrwZzh2Afkpu7WtlMuLI88aHhgTuZ97BVMSk
JVI4UDWag6d7yiAnZGJrJGEf9AQntaB/Z3eTVioobYAWPcH9taOY/K6Mmc0gBYfnZdtUs+Rrrjq+
R04h/zrzLXabhLRkDocJX/RqNn+w/Uk4jHZYiK2JjATRGdSeYv/12k0OwwuB0+9HnO87HXYStscI
5RCk+6XYEblK5+Sht6NVv9ZU5278mF69WAoeEWsyc6uxf1/Gyqct9IB3SBZzRkuqpa0J7wr7vlsK
/+ZB+URJJT+oWtDhs2fHhW+hKtrz+jMMTPn4X5B/BhzpH53qnbwH/rQNxnsCMZL+aLJwzWDJkdww
0I9Q5G61weiBkSXYoHU7RwVSqJWnduULJDznTukrW98ssc5BqP9qFiyc8N8RXsslCwey73f4UR9F
A5zHB12LycroGXDnACKO0XklvKDg14qWa5SpLRO1cT5DhEFwFEkLMK+QqUrQ3G7oxZgsPlLyLlbN
HucNai0ZHEmcVRLuvalwek+zYOga0RaoyeL6Kfb+eCr1BYRrMRTaxz5+eaK8+IfA6BwVkdlukTec
S7AoQlONcTI8Y5gFm5AZR+pjTasv2IhLOgQFPL/3uwV8uY+LKFM+JZCkNQBchUBIiLHa0P9e2OJe
C6QMTr5yqgCMorTZ/6MfTGDnqEHlOmPihAgS+03oQ5tkPyDfWGjF3FfUuzPK6Vp7kzFIrRV+2euW
BDhcFpSxPJdHSmjHn7MjT9O2rHssJPknHFUigr/jLSaXQOikPZNOoO40nuzGVk2XCagb4CCJ2rVb
1FBs6zF1+FEgB+qxVz4V5LFQBuky620FhDT5mAtdr60egLohgRhuPMeRdmTThXuxLj6EmgwItDqh
oywNCZ87xLFaQnx4eMFJ4JdO6514cws8tlgL1cxlTKMM3526qNVgm5RzbJhgGMLft8KS+eMcXlW/
k80+vf6h/EzYu9v74CvKNoTMXAXoTS9FTEHVpG8HFK8hFU9RFNbgPbcRAoKF9+r2v1edlbI4DMhs
++hvAi44NqBCJWiCMTlNhzRx/xs9hkT8fTZSSVO2h+U6Z304yx1R17KpVTX+7/RHMQCZIci1+oP4
4rBjtbHq+55TgsmpSigh0zbSrQx9bVh5i28Rn2JFuvXlsDUEvC+3ASGzGCHvrhTosyUG2hn2tjZ7
JNW5FF+xlEvV1rdZAs4J9nQpzYn/7vR+OqfAnzcj/2pzCkk3p9ovVCWbLn+IakwrQPQPC14M60bM
kp/EWuJuDVeG5NgSx2IxFrEFJfiL2EtDihyhdQJGwETiPKwscUFs+OzOCXExfXd+uB/5DwDe+5Sx
aLc6HfendvAbedipYDgVlsTuXAy7NpeVi9balp7ycsCHAo98pG25FFZzPf2I5/7BuKPs51usWJX4
BDoDpC587RtzHx9qzvwX4vQpJC4GVmaBm0jWtksrYZ2Y39BNX1xNTwPHDSbVqyOCg8hKRgH/8vq8
TgUELggCjo/nZR5JKhYqWuB+5eymoRBiVo/ZvxIA2klLnfMieGfsFxY99jqzJQeN3dlUIp/5YnQm
qG8/nvDRg2PfpQSG85k3s4MOmgQjrqN98balczFv12pH8oKx+nbtLkZmZYMs5ZPlIZHveMHLlqYi
/BYB7/BHUXCvDrKuzy/h7fV2NwlqrbfBuZqdIjSFWdkbbHBlcGGZElUV5WUuVPVM6+3nN5129+Z2
VoG2D8Jn/4WqO4wKnI1KceAqu32m/Q/xgqFsc+FOMoj7AL++9UMBioGk4O+N/RFy19Fa0NMn50sV
ek1RDyYwKZ+gkqnkmBNGUKcn3TUkS/8gUnnUGHYxjtx/kJ3C0m/0we0x3zRqMF1L9FSulMYQrZoV
l67uH3Ddnabj9OSuY4wMtgdyLwULgz06evUaWrh2CPzAWXDLTv5NZPitcPx1b6c1MDAmU06j02jn
OyiONYbK2ps5b53fQMmSSEecFQjxkygNg2zsvKb+VJ2idReC3rcvpAgecMEHlHKzxNyQWtW7jWWh
sWwgb2Pnk79EOjpCIfgt+xTq2KUXRq1HpoDPGQNvMyYMzYHtMNOXoHlAktxrhG3Wwaq9LO+Hm1QK
9dmV9CCp0++Uii4mlB4o82pTmnGcGUnDWYAhhs3rh6vH3e4IMUyIH1gPc/y038pX1NWiiU58k/OK
MBWk7xhURqKyRou7Fje1DBpbU6284jNgNO2S4Vcfd6O0AeAG8PpQIwFfOHBS6K1ICwhugkE4lrvr
f6FO9U5dZLZSk7ddKax0BsXmDgbRwWozZ6AxPTJn9b1lrfAjerpIdynjB/94w6lZjHygR4X/aYhY
WkUB/w+s/MBu5vAk3l3JQaA0pG75Jq5diQjC0bMk+2bf9cBJPQs3MVH7aJEsb7WENIBkXz8ytFsx
0Wr5FQV2z/RyccwmsdWuz8j+9+87FfgoOTtisEvHpJHBUH+GgZdTE0KlLsoZJyM/gRWrOgzF222n
dFMObPRPZfhXpJgCXmZQh6QmVbDZBdIsNdVwyzFZLVh4ck1IpLvPA//LUHLJASuvu63BfL13RJng
VoXr4fg3qKUlwslm4ZhYQbRfAMEkK0jbTvVBrNJDvBmnFAmCJl+w6MuN0f91uNNu+gyCioqjo7Ms
HNwiUGXsZC3q1z0yGsBr+ongjy9MaD6TKpBHFLBVwYl1amh9MD/dr5VF7GCmjTFGBKg6Zd6Bi9nM
GmT6uHy7twCrivmPIvdtgnl+IvjANxxp1Xzy6OQdxNNgXKf2XUEjVQ/LBjBgKJnqAG259bjjlkZu
RanFd3KqVGEtkyLDp5+Wij+f7PGYM6FEzk+Ay9utfwVStmDgEYjQlwpIhXzeROVov5m6YI1eIVZq
muu0+VkPlSN2pGpFLh2giL44NkcCjEe5LV+UKbzTMbaNbXL74Px7mL1ikUjWWUQkyB5y8vb1K7u+
h7D82T39VGQ8S6WyRo50+VJnVjiO1hXYnVKm5fEuMS578sfEpqLKBRYOTfg2G2wjnCPl4ABCEtbp
8Wv3hdHL00oiGgeQiO8Du9cgNWAZLS6osRiLoYizjA8rBDiG2QIq7XJOLLAbCbwSNDMa+3UZEl6A
bxmJ9YG9dAMYm7DxlD9ykiW6q4Zo4R0/XUBA6KuaxB7B/+OIeS/nbqlsQ7WZoGDhc0s8AavalJYz
YSGzFGkg5fOtyWGsBIZODweEiFEw4sflr0T7pWYJan2tinWoF0U8be7RWvVvooAVsEWpvVcpA55l
k4tc1AVYT++7SMDBh2U+kuiS/PYMBwtt0Ly2yqxDmCPsqB6lpT2u/TCti+ylUF9kX37ZxtUUtRfV
e30VcT0M6hdsho2aFaYZfg5S6jxtYxVDnOezoUDbTL+EdG1GA0/GLySCGBRd0q0PCaHh0DVC4w5C
8a3Wmlq3DbUqYvZMp9K90DEsHnn9h3VIHDQeiw+1WfAzi/m+GXm1FtVbk5qRkyVyxZUt5upKLeBN
D0/LEoK+l+yGlbGSAbrhncrsyQaHMd+pZJxBIm/qBXkDLenhnvZqwBPPtWTQ2bIpvwV+ECncvoG0
6MSbgEbN7YOz/5em85//LjfSQ5uK9mBYQU0QIUMDMEFkWCuWaBcZDyfdYw3WfVITay5N8uuMdOdw
cwFpfh6sylcf1tIXRcIxywR7RY2JzTvIpJ/LdDf7j/STbWeAV4tutpqOm6U9GKEfAxOfK8v/hwZN
P5o2DgSyPS9YgLXYgdFXw9JciETaxEDj816/wdOOBXXETPNgC1wRrMKkJYsLEz1IgtS5sNzGDV6C
TiJGFBIuu3sr3nkOn8qS8xFGG0ZlKPkhpDts76OaduD7ZPyXaf8mAD0yna5VXpW15WL1Ic/g11iv
xQCLBigmFHrYjWjwJ5KERC2MvB0Z7HC8ftcLTr922huCUFXOy5F0fxtjpvFW20SHawhMjMWRqdoC
Vjt5m8vuEzBxWepcf+CBM2LgJ7Z9rq0x1x9+E6TCnHpiu8TabSUB5G2tLnslgbh0HD7O0wfEr+BL
Ht9/3aCF63uS0vX1NB9emGgCvZmjPPl9sQUE6VYqBWuLiLtDrukrLujiEIvc/jo8/RZ3GY1uWNYP
SWoGi9kSb/MuqGOME5XxVDr+FL87ilD4QTscqL0Iw/+kGA6mS3YYc74DyoLQNH5l5T4KZZjYUd55
fr+d2Vg7tUnS/JXG9tdq4kpwCHdiukJWl/F8ghZIkYZKZpyjEE2idDVqwuQZOJUJu1KyS/VpyQGU
b6EG1L3CS2dPLjy9kzbbBQobsMNkCmbDUFnfPYXlJ8tKUYPSMMx3WBK+YMpm379gZEYwdNOQfaGn
8M4q7FQxV8KdDkb92yAjcGXg8slYjV9OPTfL1xD7TCRa+yA2QaIcpBvLjLJUMqpjgDhWAysTiJbd
9945HRM5wLHmzAKrDES24xEXJwSGkxVXBPaKmMWEb8w/eh4pEPpJRJYCk1wwHdL26C7t2eLbG2Kp
A6z3G/DKG9ecPhVbK/ifenGtNGuUamrpS1Y34gc//bVaah3Vcen3g63rWbxz7MEhrQm/Na4GtIY3
+WrAE7lSumsYjolH2xSJ87xZ2SNEyFSqtmnmEa4TlUFNapEGFSllHJ1W4PDrZNLZcEZzZxWY0kT1
CtQR6gesfPkt24YLKsLRodtSQFlby4b5NZCtJksM6ucUhvvnfkxiPvvKH67s4CfZZwstbX+X7qFi
jWUj/QtIZYX5dG2l+RS3VXV5gc0IZlSa+HDUW4xkMMjaYvEDgzAxC6eGxPzxwk/g1IcuhsX9RWRo
zOUZp5a0GDf4kHXFeoC5/rvDfYZhI5T+EmhLqzT3DPrv8q84jwPiyCrMPuQJsgl4/QVikulHDj6s
3pgJ+L8njiOW1Ts3NZmwE8qB56u2khL5Xhfv/xH8pRjgLSsVIi0YDHKDmHyYdOVi3tDefnBEQ18S
Q+w1dJ5/4y6RBHXFFKOEfPtsj5C5LpjQBZUOOndY9K7OVm49z49DrIHJFJ7wTefLoI65I3YCJI/i
4AupwklqnJozdV8Xo/2JOcmCHvSmLP6bi+bsGT+AdB9hTkAhAMI6GkiO8aEg4L9XIP64hth96oyQ
Xdp46mvtnuh8U4WjFrdSeMt3lh7aqw2nSNKrhpIBswVQPg3yi5j4HhTX+7dwDZkJ4mL9n3o7OBsr
cY8lbjvJQM174pUS1RffIoILoufbaOCZx+sfv91+txoV0eF4Edpv6mOv+ZSzFeWx97cYyNY6Acuo
O02834tCijejaBSroH7jKopoNMgQNS74tfqVMonZICQLpMjvuXwCpp4T/1y3ur6Qa1SY/uiYkzHk
UwtDUiF2U1/Xvhiifa2NOV17J3IVHMErbG5HlglNAqeSIHOQNw/4ri0QZ6+7J5wR6yodfp5InS/J
est3bVw96BonBIVbrkjq2RGQ7oYkQP4Z0ncRetsGtVMtPw9p/xRUD9quMNG7nwz2PLYb9+DgWY6c
DrMGw0IKIOxoLsxyYtHQVYzpDPnVRbDiYgoLba3NIlCCBHic61r+0m4qdSSavwsq/omS1GJtcJ7I
NpChQbGPO+QcG0bc0HrFZSJaZ87uSzRLywEhQqrC+DTzYQ0KjaJ7+bPDrN+/WPOaE2uwP+Vmvzmy
EckMCxyfzhLou/0l5gLdN4Pw70BMSFcAAJNSGh/cGimVsYUpeL/kijgeAvmS5oV/7LIvXY3A7Hgb
6D3WW792ZLehLUKSp2iR1FyKHNY7haSwOINSSgwI07YYQ/quctJ8iJnL9UxMYuNKcjJFsNTCooMV
WEWxTfsTI/R2E36K1GnmE7EFbV+80OgcsMgv/sf0PPphJpvFsgmieIx0jdBrTVX145VXwaMc9QJF
gHgV52OoNoAKuzaD25o9RFMZ6xN9aFHM5+jqUQxJaKNJDNdHV90egHm2PjljfEnb7+y9nIf1G6eh
azqTbbo8wst9c7/ANqsIK0moiiFLjGgM/sgSldISJOcpQoPHEWCzTeBmEQzctBx74pNnh8VzMb6/
yN3h2IAYWRHDs2OMspe8hn2ke2ilSjdlF73+1r6tllk2scQrUq/Gmo2kjOzQacyDHA9N76F9vLBX
jib74MFP1CFMeGe+aIr6+r9iICQKp8kOYKOSimPnF8kmQRdp8gF1HDwi4LN8ni1JscrVAC0JQnGI
qE4muL6vwJCdbKoDBHjf9Zi3dE3umP95QdANNGM0O9TW1AUfkaXF9+hxl6aINMQQcjLa5s2teRmb
J4BcxEObOeTc4RznbO/wwrQASDTy5mLjhQOT+N8OcKY0C0Nbe82wEWYovPFSyNdHTJNqI7IA9vKv
6cV0yOWJ9tZgPkItImn2SVm33JfK2mDfItVoTWa6tL+Ub91NaXWIgpGri1mo1g/oOYjsPa6oo7Hw
ofrhwacDvstSopHVWrqZI8Es1iM2jGVVyHvrTHmXulV4jBcsCDMlKaiEOvh5XDgTKY1rmXh6ezF8
QuVXDftabP5BoXfqQtz1tBy+LUChskcBJMPztV+ptL8g8R3kuEq8tBMFuN/os4C10nEInoEAm1xC
uZax8nBgj+W5ZwUIn5eJCF0ejNVNPRyPpqh2mEYzI/OvOBTbT9FCS+fVnOG0Z1JQ6uWuTh3qK37c
2T7yDcjiqmllWXEhnWEenjnb1J2pFelchpDSaeb9fVxPrNOz7/fTBnPMojzAq27/iIzVtiLzzpV4
F2y0o82ttR+yd6wbBF0YcmQ9vS0V8t27EmQRzyYq+5UYXSNdiixv0bvwgdH5oeHXKg7i598MikAv
vu0oF6EDDQDeTRIXVbMYD1CR8tRsxwwGOzfuQex91CHii7yuMwrLRb9/3eTJIPbk5MseesmZ178n
T9CjQWY/0PY4l0J827oHoXIOVT0rpHoM84IWohoqd9G0YT7Tm7w4H3uhCAsrWc5uB24mV1AZJwe4
QMn5i+G4cpk6fLUIDIOCi/T8EwzD2iPRGfiKZN5mUNPdBS0Q+8tQh9n3o8+Z2/H0JpqMk4aUcMLi
f9y/lrA0SY3qKcsEbW+iD7WVK7/eDR7g4E7uTtcWivnP6xWcReAt19zI6TqGpXgfMCSa+C3yi2iX
+ucIZfY2LkwQicvMSO9bY+DRPIoVbYA1nxY3GaKTrM5zJnLfsr8Qhu3nh+pp0x1RPYHUPYz5zlWO
9shMUeFcid/nhdqvmmBU/G2VdyrF1/CHzbvlAHvumOUd1faqJNOkhv2mPjS+FpeMNzUryPqGFZUx
bhfHBXmRHvRISy61GL8A/KaZdxuKExYdBpvGSg8dpVLgVSZZu4jZmP6oZSYfugr274DldgTyd9rK
AWAy6tulsUOf8pNG1TzYcqcWQUWPQ9KQ/OrfxnxARr0WdGT35XLrrrs58DhlLHMUZ60qpf0non8J
NOXKpLCs5h3PfxlExd53jIz9/dDYWqf+05yh9i83llELf7u841PuTJhJoZySwdJLheTQFkDoB9XR
74b+DW6IoelRQf+n6dJAu2wtDmEd89wPREUXRCqp5XjcbSetTL1NbR8df6W8EobP6avPdKPfG4TW
At7mToihoZftuYcD4BQ5+1GDYl+tvXk/ZwzLLSYo22ztxGwxiYxpDIOm/GUp94Irnu2iQjuCBo24
3iJQFMlX2zvq7vShcoGeSPN8bSwDSZAyMf6Y11IU7rXH6xiN8/+D4aOt5jHWk+lVfZiHm202j8/M
//Oc0YlgWiEoXCvGkRIC9WNgsZUzxl33YcLcyDJaDLAWbyAouI9szsrr6N1ThUXob72eiTY/ctrt
/hiwEJfMcQfQt/yOD1HwGdLoxyI/Kcq2x2oXUTKctZ2SlgyhCBiDRpuELp9GP05vfreRMVlCDBeI
nDHhhYNduURxgUcdAmrqiUCMj6oDyXV8xh+oLwffL4ovS2dN7ACBCJL9OKF3OC5ocBFsQO257M/5
4ik/bOV+gozMc1OmRMk9Ylwg8BHVMyhLX27AHgNeLXYULmV/WPeykaV6ql6mJ6Om3MOCuG9l0std
T+osVrFLWYK5TWu2Q+YgTJkR6pRHROyUhsLcK+cO78LVnoD5sPEGlhsJSR0xneI/CNr1WL58zXDL
q4L/Nw8zgcK1vf8t5nwdJrOJIXl5UamLlTyJt/t4v6TVQQdTZEo1y0WBopyxQlTWOfe+P5tO2ppI
PNKNksXxVS7ooEWUXNwMzNZn1WcxqXedjbHWRrk+x8uQNyNyDjdWMx8ptloaPQSBKzlZzECxplLU
rW6v1U5LJl5ExyakanB3ro5xJ5l9aMup46RKVUcBw2YhU39aQHSky/cx9RY+3CxSq43lvD//kAqd
UCdqsbozZpt2mEmjMnxt5ZoVhBuFUw08LSHaNeMk5ZfYdABtsp1np7klwlG4wFJjFJ/d5IdSDa6X
WeLPddWA9GIECqggR+a6YuBu2mIluyQbGAa/338GSA8iUqZ4WkyAawmqbt7aalgopV5RW5FVOFao
MV4ioETNFc1Idf/B/OZenOTvJsep3+GhkdsuzSRuBYz8LZC8FJ0NoSYN359vLOfSPfdp9gTTl7fm
cHxN+2CJ5l6eenAL8kZRrMygo0L+bU9uSygT4BdSmHk8k9ZKi8FaA1BwbdOZeU3Mr+1K+Y697fVP
SyDDtFKMHMggvCqi/wa0qn9JCxoUAYttHOaQxul55oM31DF1yVb+/palacl8dyeBQVTaUcDaHtkU
+EwW0ECosfy21W58iPwoHphElLzIydryFfY6vA8T6AIYGUPUrtsDGbDD2DiPmoCccO1v1+liWVqZ
38haJ1ZEnrEy8IAtd0xD2OFA1TEkDliuEPiIsr3PF0t+/0U0d0U1DFrQcWQKp/X1I/bQmVMfnFfW
ONwgpmsSRz9HiQQeGSQXha1siFw9R2qHtB6a+0DVIxS4T1CcoP+Yj0wa2k409OBq+6dP3P3idEoa
oXUPQoEjlwxLlI71/F5zhobCFGaABtDMhs2/zhd/pWGbtv6vtDuaMCEOTureHUe5zy2XTBmgtqfV
sEk5EzfpviiAek3Uwe4Tgp3UH8PahINSUCV8n567TiS3sKFkZoccdnIU6eT7zQvCO5dAO2di+SCf
QXhKQ85CG94BcO+z9AIIlBjoF8Iz7Fg/tDlaHWprSF+ODBR37cqH5Oqs84oIDeRkIPQJIG/kNk1x
CKFWw7Faz9S21KMh7z54gK7cWfWiKrCgG4dfRzw0uk7GmUe3dSII7Ev0Tdw94h6eoY0R9w2nzCos
I8bhsAthCJ8wRl+xkmE0NGnSwdREZAuSVk5s5dcOQf61yriNYT8ssZj5m7K5pYhD9X6ilH6yxVX7
lImTl4BjJkPllL+4vmVpbQgiKXCMgz28ttBJFIrEmmjj7hX/uNtmvXusPJHFSF+Zoj/zbyfHceKO
hX7b5mT3DWTyV0ipQXUL+3tUYd4g2CxWEJ4/5vOp1XMpyIxdU9dh5EYi/QzSgY32YBdIvoz+CqlE
tEdARou8kn0tU/KPwRSsTsLOitUT2EhGWIQ6w9V/DI/R+Npi2il2EITZuFBr63MJ2RO2mE4HR2s9
2EgmugglouClcNNBKGZVmZ1TljXmykzdqO8kA6Hk7VItjai1aHUCJoS/1RgqrvqLzx5BvB/UGlkP
LXGNLWfAzvvxAOzalctaOlfg+XCm36mqNPh0lPxkGSBpjjTA1hfkUnrPnq0mCT3QjYvZ7xpgvD7v
QO3+g4GAJkJrmE53EM6q6i0fKYygR/Z8//Q9QB3191BuE6WOLKnDzuhOkrdETcjCSii/dIEDw5Da
w4R/X/erVvuEy9QsJHc4CVnIDgT3bE8SHOGNcb8Wy5Ux/fab80IqIsuD9MzfCx79iwIQfYbNnLtV
RD27WCMDj+JVOutIBdfOSAb/sVAJ+W6VQ53prjhEtAbRINjcUtUBC/Y0zbX1AjZ0i87Jsm+xjtYe
sRNgLnpzGKQNLeTv1FHS4Cm5XxEnpcJyPUGo5dzWG5liAxOlYolD0w9of3yqDsAL5LDljIuagZ4m
qN/IOe6mz38iVuSbwJY5yxL0WFHZYvw9nCFoNDBKssGPc66FtC1wqhTQpFU2aG9eOGGJ52CpCz9i
AKw4hNbwXBNmQATrQESUBn5+QBhQyc1xkmA+26xX16QUP4RyQQEt17cE3zjeYgPjBfbhVG5+Qqng
Q6fK3vfUVTl0yO3LjDDBLtsga+D8KR8eai1pT7Kp1koYZjorAgLts7M8f0V46XkybsEAUH+GjgJg
kRMi6bfVjh1QTg0+UIiatTL9q6uQxIYNPKmg+gcOkP504LRCZHPSvx8agxJjhZpYLP+xtyzTbY6m
299xyL2BUpxEGw9jq2DY1fCXG/9pPLXzTTvSsDoSaEBwN6fU7dBdoZOpBtJg3KcWVUNWi38UOLOB
tNsZFvOXQ/EYmzw23OmDRhkQEsCQ77SE2WnULki99j6FlN8rNuZT6z6HblV/y7lTvPDq+zyRBD+x
IhNMBpWWrojtiq69mT+r+jp0HO73JrJ6gNiDOr0dBC9mA1665xSXDIQVTD2nuNkj21wqadVwNOsO
Dg4jY57YHZU5AAXvKvNsihy2+x1NMIX0ji8M17e7mYXOfZ8a/rQYm+cuaTli1PZDONT3WSR+l/q3
OhQ95oWKyRK7Pb4iF3p82coAMeueYCsyg/NKnRwukRAyaHtQZ2sk00ZnuI2xBd4q28DHrDrf+p0R
OjSElovHluhVB2/pOy7m8NqZTjr+0uSI5B5BkYg5RMiA1JAX3bqIr7KvqTifPCwRwE+uJxMmrtVI
SsnFnqpf0tklmTHPnGzvdBw7oM9FT1U9f3zQlfEcOKQ03/uoDVQQ9SqSEE8gxse9eXatK7l6DtBW
Yzke/pE0az8QwB0NRZNnMZr/I3txm4XKDXwqMJDHRcE0BZK+kEL6NNMSIXCGuJi1W37UfTrB18qd
pguqHeN+NK83qv/vCgfsWBsTgtsAZjFf57kdjlccKpsAPDEIXIvEMmNkQCFqM50qsmIxk+dE0AnV
vZxUYFhqenUPvE40AXSqPZMEjPk0iEn/CifNRvotjy3zawUVC0c/40M4qc7YAXMInRwIo0gS+nVm
pnrB1UYyE3+vZDCtWQJ3PtZzsqkEm+Bm0i8MR14yMkJmgxctuh+mzcgFgbzBNIoph5Dko8udpGDq
e0+LK97a54iR9/27RW4Vcd6D8gM89bKvzmKm5pvWSRQIEHTG/+mnREGw5IbfIMh5JM9FyMezWDAx
B58GkaEW/KfWw3G2X9Pg1pKoVk38eX5wztOCz65vsVdhRcNSiJn/WOKxwKwjznKO/BBhDs+KAl+6
G8AMR2jQ47GfKGVT4px8V79HYBXnkcImr8KfRgiZ4nTsULbKPmmsvjp7NUK/0E/dYpaSPDGYI531
+t3AjEdb3Tn7+WlN2ITlKtHQDaCcYyN4tGWYBI1zYkjFIy3XkrJzJA4S7lvs8oxW+N82IpDxx2fY
hn7YaMgShf8omhA04HWHfeGGWdNPGMMNP6kY9noomdD+0mWGTKsSFjrYL56LdLUngQ6SXXTQt84g
SoBrcLh74NUUu73uigUqvN4uEwgzQyt9QYHTWWhAXC1DRMgkL61hWAftmR48t8cI59khoDesbp6v
5fBzc5z3AAgANauEn7rD5tEeewf9iH+aPFfKBH7zwlGmQWf75w0aSJKMq73ZFH8J0UstyYdXVfIj
MMBnIisYTIzMlEh2GrbeqxUM2EFs9klqaimwl6cJAqd0p2lsuZ0YN2ekzc/Z1R1LAXk5SZQPMxJs
F9l+hQJP1BhoN+UgwuLK5nEDEEhwKoj8eYF58+lDpW0QhLM8BHBFVf1dBiXsQdPnvE4JARCFX6ph
VQSQ7JWWJl38QOcqSQBHSMABrcJLBf6UCfDyL6DeihXzNVTyO0szq4zdBb/e+Z7lZ4+b+UwHPU+b
IrgsYkGYOnG9cneiIrE88Nn8l2gAqK7g+W7/6ogY+F7e0IVaNjuu3c0zS1AW5lbiMR/uIYpGw0La
IRsgNR8BTWauf8lbmGiqKr37imWe6643wyvguxPdwLX5lp94WrSkGAwTBnkrxocxwLslRg7MtsSp
ez77vIl8XQjxo4QkjBQ53lo+HnzoIXS6Q2nUid/lkYzHxTTFeQMs0AeI4JgwHfb6lP3ncYFfVlGl
YWRwdSxci6ZyZUnbe03rngFn24BAVcMxlme0objlBz6RWLnHHC6q8RKlJGNvpHfcHk+jYkk09UeV
FPLneYPiXVVZCwNoIk3jCCNKIhxmhxzpwLNbH+bm+g5mcDVAI873BfYuoBh/eKqezTWlsoLdixul
QvjoMwr7P605snrZj2Ak0kN0QWEPHAyEnzsLh3E2SCrMiRJDHUZijnCT8oo90aEw/LPr273HGTc2
OhIngrAHbImMW5kp9mFL7Tfpe6Go58v3ValVX7J58wIdmyqItuB5MXOa4stijwb137dYphxwqBvq
n/5iH3HquOM1np7LqoOjIh80wpknW8oKILMDGHHEvMf/o9anrpl+g5LV3Rb6e7lwe9pP+yUdhiVf
XFlwzEgt0eB+WK2//zogEvT+H4cec1BT3Ar0PMm4Cn1tWus4Cz+e0lMPaT1mEyqPH31TZrbjKLYI
AR9wOJ73HMP1N2q+NhHV/ETQI3s2RD15z+vgmwp9J5g2+K6mtpQGuoeu/Z3a8g1l8YAY9eVmj+MU
jHociYm53FdhwocAUMBsTRYUI4zG4j7w8Q6CZYEb+Zi0MYQahheCkzmIbjtOB1ayoJyC7dJHWXtj
7/SjuURrf5FBdS4Ztp6j8cwuNTlh5YASZ811Sz8brg/Ct5nRyuhx5H8Kqxk9VXlVpsyes+D6mltC
7VxYmva6vTk5ptOPRuQAlJ1glWY3IR8x2FrQNkhHGWO0W0CaFnvsZmg70GlzZnZfa4IJvqoAbTL2
wQNwZO46VOsa5YDSs4gSir9DWQbz3qW7w5qnF1qKM6y8mksd9SW89B0yEoh6Xy170hIOI4D0fLTa
gE09eoV0+l0RXtYqKmqcyDICglApu+URxtJwIC04UuoG6T+U6c+OtbSqO8mQyCkJJ+VFni+Y20fm
sT/BEWjn1H5yCLj36xUsbAPalsazYpzX2xg+sFkwuH9ypZUXzYAUNfN6KxMGruM1A4sg/NYTW4Ti
RWPOSwvw0q0hkzoMrNVcOILM24fj5uvF8EHB7Ua6wPAAGk+UIRAjQzcmYOeEfngrwjyo3D0XTMZR
APMQZvcxx7gXxKRmmqTIXdthcyYM1LsompotSaKzPH0J1Zh9sJgUARsqNYCaOdpPEK/jTOQhvvTQ
mGTpR0wNe+HJoBIFBbHFs0X9HPXJrxzu6qIog/pblIfO+13IVc+MACIgHRLSdqlJbakhTcJfg0Lq
WZEf/D68jeSbHoinbZwhBCJqdNte9J53DS/1SXqro1h3iMF14iG/l8d/Zc6Uy+dy9ERelnQr+ntN
L01H3uyFbhGetLfHMDgv70erPdJdZMZbx2qU/4YKJoqCFl0JppXZDek6fhQxE6tXIlxfp9qFVxPT
q1WpXLsl42Imotn7q1ihybnmiB7OoeHwVUbv+BjqNHnI1GAlObYSdhBAycBgSQhYCZ08HuKKE6Vm
XjR24H2gI0ptguDAnDVFFOvMmUEbWslf3IA9PrUBhRXLshdbdydlRIhceA6Fr23g8GesjwxpbirN
n4yh9kTVj2ea58uP9lqupq9qd+Tciyc3U+7YT2DBbH87kBYgQnRwz7S+gju00Xai4dcUgY43S1Mu
0owc3JK3DP91sksaT3ab0wS0RtJ05TsJSXdK7NXVO5veQo/gZT+FeomaPcM5aylYBxViaMTagVX2
UWp2Au9w616VlPL3XKNAp2Z/meWCzLgh3ngQmFyu6VUQBFnqH1kRahJTvWb7Y1ciN6/MgN13tzyO
H5DztFdSjfVDTa8vQ8tSUjcpYVGOQSLLyyWLvknDTGgr6Ob4nKs7yWcqHlLkIN+DSnfEc62MxV4S
/hEv+kWliAJy3TTP12YN59zcd7Q0SWHoTDfU+z7i9wkJa7mVkfKTQZNEtm38piLXgT6LyrHv0Ezd
nqM5u0B58OMX9etxJwayQXxUEkwBoAyrMiEqlTGUZn+pGmUYu6cyfn0PR5z5Q2W4F7/Cus7a7hba
hDeuW44/td7D++alkZ5CMM8B5FjxVXfGBsqzjhiF6xGDo57DDOiyw2Gy6L1UrdrDpMuZjHsmI7yi
WuAMMigYOEnT9UJ2R1G0EYmpk0BMeNMudKVJjvNtpfZKGbVJ4h+2UJXGoeB8rMUMjUk6vxUMljvx
ZUs1jVc6NJ82GkQ/FbZ7g99iggOrzR5Og33In5ViGF7k/O13iOGKDRBQDHdEqDfkY296rQdMHfEy
8O0CD8d5Ha3zDbBHnzv7S/CW0HWyCq75iXulpA51Fk8IGWURlP3xRa8smLpIKrF13/B0j1rXZlWl
tkqzrVSp1kkW6ahMEVGVH+2a+MV9Rd344Fuo2MDKn7iZ6D0h9H3JZvzMMEkLpKyBXdxwBi/hkMpQ
2tFuS6exN8ZaaYo2lVND4pIiPeBqSlxvE+tKvePO08GS4F5fbsnue5jdry3qOsOXLeLsg1aCTVZJ
Qhk+XZjoiOdO6OITTJuPKuKxzwU83QXB+CXLxvNvzfR3VVsTZmkbRDejlM+iBAmLw0alNGMBv5SA
61wrx2NKTN3rwWmNsj0XqRJ7pFxgeRDMePf0f3AEpsJ5An62mluDNWJI5xygvm186SzWQwP4MXUv
MmcNED0kq8oQrnYIAfNUqV6P5Ni94Uae8WvYvAC8MhSFv+O3W3+CwnVUmc6CgZgYR8KX0WHzFP/u
WmR/Ar86y2dMVDsVV5V5eVnfD8i+gmzcaIkemNrg4U33YC48iQ3cFdt3KiLv/HWpS5WR1sk7pOGk
pyz6Q5CE4Z2F1mR6B+XrFKAZcW8oOGrVplWkUzH7g3u1pgScW6CQZjHWD9EF8TzapqlZ5/x9IlCF
97FNX350aCsERSfpF4B5a6PvS5OGsIaziu1iAn/q3kib82UgEcCs7J3EjBfpjtL5FmcYjJxKIMY6
oaHxMJKzmng88+ryW6W8wOl7M66eja8qvUcMuXgrhxJUxmcWv9rgJpHyLl2kpFWd1hoTuuozB5I3
nbPIwgW1EaxqPZ+ac6y/SGSHkIaZrnwvm9JULX/VAAWPTPgIz2htnmAiBM3rSfsukKiyB2mcBMBn
1eUZaWTCMdnUBeD1Afy6szHLcXwfEQ18fccpqqVHAoOn83e4svDIkfa0Cc7yYWqVl1C7XFPZjMfP
Yt8JiaMGXr0tqFKCWHxB+YTKcSVjqKZcvmc/jGglDzc+G/KS573DqKSDa3CKseUR3OEGarcv6BZT
wml2o05TETCX3BFF2tX4tD5iMk0mlb7S2D7Wa3V5TZST0Dw84P2OYFDoLqGjteKsfrOTQvfNYC1k
5quu6nxG7l18742eeblOE1SmRJQBLOr/BhYBLu9bXVkgix32+8sxviW2EO602i2X+y4UTQnreQkE
dTE542hRBlXVQ3Sg8jJkqs2DV2dKYhVoeKgtzaEpObpCGSG9xVjZGpRGvSAf6KluunLeyftVe4Ep
6QovCtNXE69bZoQPlL4Bzg+DBW9hVVOvH7RlaxCnoiQJ5fXvyzft9QHfCOcBlWZ8klMko4G4eE++
ZRB2UMjxQfBidZnlRxKYj0KsZXpxzlcsF9PuTQKBZVjsbdbVFo+hzxfTg4EexAghJrmHVckTDIe5
/UuUUlDKd7mdK10eS7TJFwmw5MIRXFWJ5Klvabqk/6PU7OAK4dGVYFE1HEs2yZTKwiuRlPtNrGTM
srqABZ6HodTp4+v2aEX2xKtcekBGwhWGVI5d0PLcgvU5iQOjd62LyzV45eFZRj5Je3nMm42d6GLa
5kdpBnivpKY3so0dIJG7X3e9ClYtNVYEczq/29ebGD74iMITGva3RL3biIVs5F+rdoS6JXchWDXe
kVJYgNue4U8DEOhxV1h4UnNk4wZrB+JnPG0n6N9+kBWzVIwaK5m0sdBKpSbTDnOnmSwZ4MoZXmxJ
UcodalQT6A7rDztg14wzD7oB4d6zlLJ4wQI3gDJYh5E1nV3eCVUEOOAxffi24qOX0nHb8ylV/hd2
cTX1ccI+21sodAmHsleU3QufmqmWOchAWIFs8aK1IfUfRR+rK83phj7kVGDC1JKtsIFQa+24N6Ch
/pluA43Ympev8Zj5vh4eY4wvC6tTubJ4vtL9/rwDI/0dEmvEHpqMP24HdWMPkEL77KeAjOnWJ/3Y
aYueIgZ7ZhCk163IXjMGewuCYE8X/LUoJ/vklEBZq+Wd8tjEzyRHbLlYsuBftJ572he92pxpFVwn
tl5K1blmQkIf7HNY22SKH0MzRTAkkd3P1alsbg4nQ0FPQ9SqwC0xMePhcWa75+i06EfoU+lfxglD
zmHsEUKGU2LmcgvEk+sGKLNBEkihEYrZ5kt6jdB1uSqbqDukioioK1kFiC/+dm7KrLZSqjH+TtwF
d36ckzEyTJOtEo4fvotL9ZLLp9O7YpMC1TnBVDdguvww+0FUROwuQVo3C7jDFGlr+MK7hBhb5jhv
l7vH+HgLuBVKAUNM8NWjtrKLpm+z/B0AY8SK8swbFn6xdRe6BebtX/1EiEuThlaeeVRSWdexK18q
esnPGBTfpmkDR+IadAyk/tHeYLQDr2QXhpnCR6FkWl5ruijLJi8kkJIgc+267kuwyQ4DlAhM5DY1
5rp55V8dVtJMCLfZy2+ZqYDCH/ZX0pi7bwnbqiYz7+zprd24QUdeBEScD29pCdZ/dyqHFeemKLAu
FcQd+oOwtoMK2OYosxLsX+Ens21tnPZr0APbPEfkP2W3dN/xZuGL3LPFneyikvEbNv2c4aEsnGdP
rxMHZDY709b2G7wxHOWtIvymewTOEeUO0hXfjv8uvS8bR9aU20+Anj02I0HmermX6eavS8/0ej4H
oL9D0KhT9KpzSo/1O16CqfA0HuG9R74uNDsMxaPJw+ZGvIGQMxdD0YNEEIALdZSo7tyoVBALlXqS
wnQuEF/3HQw3FKKqFvYzS0OS/q/K7/CaCoAmXUkAPWFdUxJGpxppZqtQWSYfy3Mpe1h3Wwj7VWim
65AwRrxYhyY68/6Fq5Nxn8Sl/3Y2m6apC6JuGNT27nfzioX3Kmyf0jRseiM1XMxzLD8e1NLv8USd
dac56AIqJAx6nshfaDp3/WpjbRAQ7gDcaAcYFvmxw9S8bOgR1HU8pwr5uM5oREPVbEHV/p8vvqcx
kXZcVo37FfdbMGXO//nexdFBFGrESxzGwHp5b6Si95oQpQ50h8eNTfYMk7hznZ5gacwmFpLYc5cO
xYfYxof+mFyXiYGKe2Dn6e6iPeVKzJDTvW6agRU5LGEnj3lHZ8uVm37GBfucCx9idGYDzuXWVRFY
iaq8tpwVF8JTG+E3Fr0KR97XN5nCdW58yD996jzny14NeUI7ZNRhD8b9gJdzLY6ps/kKcgBaFJp2
13n7Tqnump12sBEZkN0Y9lqlVqdqxZ/TITkxT1wDv/d+B5vSWkxAPxsHKoWQMaGHlw5h42Z2jmYN
DzIk3UKpY081IO4Wdsz7Nexuh1Qzb2Rhwn5q97uiHDDV1/r4QBXgoaCL49OHgbLhpLm7b+rDWRnd
yaznvPSnZxlZEriBOOu7Woo4QevwVf8vV1gD6mDGzvxRRu4t10TPkK+godyq2R4AUGwCo2HUCoHX
Aw3VJjTpdgykHpsrBt9fNrR5irR+irZiI5OqV4oNuyBenujLv6q1A9nnkwn1/ItiBh0ndDxHk1Ny
2m9miwh2jvCblsbplFU5N4gG6v3rYqEmgX0KSrfMnEdqmBCK3RpYgcvbEWSEUz87t5XsSqDgbIkh
v6H4BYCWmumHk1x9U9IZkxpa2HmAqZUrHg37OKRGWuDVKhH+sBN9/16qtAL+fl4955SvOSAWtsJC
LkGIiWcFTitGnCVA8eH4SzG43yVT4OXimGgVZ5xLhnajlDEe8dhzeYAl1nuo2fuokZ92679Wg9vk
PCKTcS0QafEh2q0DtYHQmVqEWhGMbN1tfcCgBW/punA4xHNxA+JqwOtnOd7t6ylsTv6jY6W4S+4l
salPHt2yBVoC9fE4DBejjSNzPtDmItbhva+1qujMPdEa4qWH9wkJkj4O14kv12ngqccXM30EOrdb
aGQNgNlv/WSKs3S55hnk3ts3V/s71dBogESabDE732wKomsI3P1ovFcidHhbuRPQkD9BnqWFMn+n
HzjOb455OKLWHqIevs6mHfMarqrjokjIOjKVKS6W9cQjF99MOQYmelh6HfCa+uklO83Abcaknkf8
BfHCfLhKO6ZSqjLFtWDf7LMHWX9++Vg2cqiADmPc4keqvr1oLf9uTPTNI9gq9hWE1CFsZurdDdk2
+qC54iqUMNWAN7/WDdOlWDMW/dJXoM8HFGlPpL3wL+eIr1SMew4brzoD5NikZkppUevJwV2stkWT
wxlWyXY0oWqXSEaCTM59EAozsCHx6uCFqdsz6z3psPXOIqcg8J7GaDMhcVfybEaCejiHIraU7ULK
zWT8YKbHtil1+nNfNbiscleR2ElC+EPKSNhEokJGHhQfpNBYBKgIG38N7H1xNAb0n3EiC9Li/O48
HNXWeMo/98g/U2mOVuLLToj533T4u94PFq3RaAzbaWCp8YH0Fu5Dt8cH2R6KMHCSAS1vFEiBMg2e
JXSRSMOurkUT2WJ0PAyXxTENpxooa7axuJRq6Pu8pLbWS2Y2/vEeSX+RnIwc55EebbbSd6OWFik5
SA8Z5r/hbeDE6lpw068Fz+S5he8hR3u4F/aMoa9JibSV2CCNkvLQ8itg/Fp16CMbv1CFeYnfdu5h
PzhW57idWOR4DNFzb5Gc75oxa5v84m6aTMtf4m7hBdR2ptnyLxQVhrtg4PfHNvSOkoVi9S4X4ebW
/8HLDk04/jOA5CqoXmjCr9Nw8qPxpO/jdClA0QBnhCJgsvSPdOQZ6vLv9nn4DIZXTSQwsm+jhbcO
EIN1dD/Y7XvT/yrYQF9luDPO3LTmcXw/eVPZ5CQ8Ow3y+suYMERyc3h7++ErtOM3uICNf8BsOBtn
Nr0ldlH/ij3QtNIHg5T2jK4P9/tXorYQhnuC6YsLZjCsorcRhpQMEVTxfRdk8JMKf6lzs0EEL+gP
H4d4crb+wfxo5hywBF0BmVPzooNN1ogV4CxECTohUkVHsGAlBM8PV0QJwZzB+4jOps94SkDPVWI3
HM3P/E56n8xLXkZAV84OMUevECuHVxZ4yigX6Qp4ZmJ3ltpBxdgMf/k9JPjDZjaxB/tFsHAfc9BN
gPA403ab/t2tFfAE8MMRqqkR3dsc+2p6gDZm22NLX6l7MDr52tEHMJysY8DTUv2QwoWaEwAE8zVw
b79sUWO8i3Z74IeY2YkAtAIA0gdjD21XnHDtt1AvbZiqfehfsZ9TLY1IohPaJuJhYhkZetOlk7JW
40GmlZ91OOlWW1VRbtv/JBg5lQc7ZSNpeR41/DagshcnQ5D+mgs2XoKESrnz1cDMAh9VP7EsSbv4
7GM6B+4HgoTp6D//ZC5rIt+FA1+Eap3vDEdg5Ul3Ajltrxvc8KLI/ZRWT7R3/1V/egzCpKYK8C7T
CXo5CwHDF64EG+AYSh5e8FHF6e4hojruUXMpbXqLxhTyeV9oCh1Lg4ZJBuYvX6zV1pwo3s/IGIFh
1szmsSIfCx/yJm4tLmfwTLE1ukyJoCQsYRSCeeCtIKVQp9tdGqIEivYpRcRu1I/v2tuKezx1CwpD
PjWuzdcX5YCsuqnKlntF/77pgJ9gDIzqTWIeg7rTQD9ZI+0Bl82g+4h2GxxKkVPjZ2wq78KlUAO4
wPcHM7nvfrrRNeBMXctZd47VDsDRNzkLvuGTIQyu1KF981KgCi0xEDuW2KpM18+e6a6y8J5jCxtw
E/f8w5jLw3VMWEq69kudq5zOqlXAT1a7MSG4NrkuWhYA41gsCRQUzyG9Bp/xrvPkJ0CQ3FEgOB2k
lKAXjFIX0dkcTB0eNSRSst6R9maqMx56/SUpuRPqTupiRIG0Nbyhqi5WFWbKDDWIINA8WSKrkIfB
Y1E34wdn2MAkkXWDFZDWxJ9qqc4wtXPdNFPmWe5ItDWRShWRvjX1bNDnqKui1MGgNQlifbnE+Bmn
0YoduDwqQ65+PL+OoDBqfWHEOrxPa/+8tdtDNCI4sqeN1MLqtVJNaezhiWA/r7wjBQ3ce+eECGTF
w8dqtVK3rcGpmwzOFTQ1DFMxiBNGQvgXzj2ONlLu46YolLfOD61UuaK+rSB1ynH5hPtCvO/bBBZR
cjpMnhqca0uSJeAPabGdFM+3DUdeQa8AwGhlIg8Ayb0N9IBfwI88Zix3Vi3b+4Jnc8FYIwjgl1NZ
tXJx+Im8MKOrwv/PAE5ix1Z3Wd5ePCXdtosXKvAzAjdbdgckCgzSa4BikrSeEwnWOcYFm+aCAsZN
1XjXZmPmUBhbJoB8YvvOlXErr22xmQ8oPvp/2jJAmaDCNgHIbQMLY5rBSxipQ/kRTA0PitQLM1S/
HWqozwOGOtnsfnvgnypY0d+5MAknkMQOEQnNEdbzQOin/7xA5WvIybGjICzJa9xgnLe8YCsQr5Fm
J0R91xwHLUjhI4sp72ZGURYUGTdUHCSmAVipDRcM7aONH4BYfmKDt1lHaNLha12sEMsy6TAqDWf7
mTah8oP0JuXNiXdgh3dQumuLQZc+n/sNqNDCJEZiDT8R40DISOjaOW6t2S6C1zLw46aUp2JZNOxt
ppOk9uPCBymoF4JPWvTBBwaYN7j4MjGMSXzzyM6YC2ZSTy17bGs/Dj1QvNltHZ4qSE+tMPLwSvob
mjV2yQsDGoKSOB+PyViSBETUe69kzIkmgIWPStRcnsG7JAgjJh63WoepoTczVeWrd3I6+abWSafL
7B/k9OtH5JhhuLsBVwvbTG7oyOriviDJahIO/w9YXQuTEsSwBXeokoXmcCguSDOHdJoRXgz51gKJ
R3pISJe2C+ih/r0li4dWM30H+BpMKYsUw0LUORaAfoA0NcsmiTcMFLP4wjvmM31LmA5uM7zYhqDp
zM5P72OMVj3O9yfcaepYcjBG2N9DMoOyZlvf5pSoqXmXUtgIYrQO8qrKydwZP/cwhpY5EiE8qQDs
mnfcGiOOKt8SeWdsTPGcTmDlKbXzLggOEOC1Ej4QQLzFDMqv6Cigo8ed8YJB9Mxkhb3vf8JDZHod
zwK4cCXkNzbeqXbl1rpLPmBhT5LBJYm5jhx2t060MjJdvIa8dvCCeVdE7USCWeXX5DdPSwwNuOkz
oVJnHRnvv9Dof6TKKx6lfY0BjeB0DBQl736ah9g77MeECLxM1B2MLxWoPo7ePVmoF27Dnc6RpKjK
SzWyvEBnWVeX4ZGb9DetWNbu28zlfMeHEBZgIxxqywjNplgmx1jWdTrlW5GkBuLiqq0CH+aTdVeM
c6aUM4w5OEghVnCuqnEA+iJdk4vDc/rIt6v1SZFNR4IaoKM944mUzbrOkhNVz7vTybic9pS/6oMn
elYtKCZCQEPFcs0kn2zS9F1qysBBP96BefbfaCtcIpKbCLoJqcWoLoaTmAX9O/oo+Q94itMNeEDI
k4h+vc/ORwbww94YKaD2z7Yap7Jvxx6TKLllP5D/UPigoL52IWvqLt1izLCCsy5XA2Bz552LfpX9
YEnjMlM+6BPg1D3SQ1V2t5y+lhoJPAIQqMwc/0G4kwXoZTc9TmGbobCf0/learkI0Nv6tIh3y6KY
Xp9UNx029TNKMgrYTyF3GTatjpemUpIRP1ICPcGQfX1AvwsOAJ5Wk6aDnf4REDp11CEiLbb1W63L
jhdTy0M1v5i+a7dwAVXddp560MMW6YuV22WZY/ItV1jSRGRLdgxgR6LykZqxJuwFcLRDXXazjOfm
E5YZrCrrBv2Ihywmsycw+3mOKo0L8Eq/Gmv7GjgDSlORLyhEFruJh8m0GVX9mCNgrPzfHn2kfzT4
3D/QpkIUrn/4KkMkluaNnOYkKcNwBVRdRXv6M1AdJshbqGX64mnM2l+2GUJ0Z74gQLBABLSWJPvZ
yGtBjKBRtLfQ7l/BXTRw/jLZ5svnRbeqPiuv+Ix+W0bvphiLfeekuQ3I59zyCRL6HYcrt+BV/awR
0QmJNLPHSq5qj+rZ3sMyrq/gzTH2GRRLjs3bpasz86FAJkB6Hb5oIlcowf2Y/r1CGGCOt/3w7jgT
LZ/IO7B8n1gD1cgYMd1FmIlJ9vrZekfcCBHP0y5JoLbpjPVGlJbDMP9y+mxMGUfsXvZyGcMVmbDt
nVI59dbMWiO6qPVUY/cCRIauJJ3cwt+gR1plepXzjxMxMqBqKsA7B3TwGtG3S1uMhUm2Szk2tDsz
kzWZApePQoWMS32owP5lo9HlFfdXz3tlSknSRUvTdE3bGoZ3c12f5V5uiwiL0TCqNVIbsJcJxiT5
/JM4qnmY7u/ygyKCKzu0XG0hmsJGhZDqx448Xa+YMysYYUk2peleOxWfKhPaAffJ66OQrFhiIwDa
KJdR7mIWnRIIuXisvVZhoV74K3yJ5u7QHExwzeBnCMf8P56Ih+ty2q03NEmW0z/8cUVUtyI7NOAz
IhTNO3oMLxg9wJYvxk+Wpocan6elJccaORBU3ZB3tLq/1L5fIsXDjLuJPbCECBTlgfCKy+kaCy41
hvuHy5KFyTQ5SinkgUwwtKH4fgv8HqevedTQniTLdZGeAD7pKRtLx++vJhjMFBmBmW62G0LxvPxu
ERPxF1U4Rdw2QoeT5n6Q0dwWDL4GVYE9+C/skCSHCGG2y+/1cvbkSQ+1Mu3R8A4RHIXIt8mWhWfm
csBnz8V5EMHoxguwpXw/ZaJsHIFxMzinF1dIxGdTn+0IqT4BoxGdrcv6MWeYsB+lkRmdyPgdBkmm
QXywLC+iRbdjE3z2w4sygdkLiQu26WUZyPF5Hets2hStkiCRJ06wZ8w/YcMWGV7l5RN6/ZvPi443
yz1gUn8lrlAYyDjYWHjVBBIMspxXVyBIc54YRyGqsbM6tWUqJ/pV1fl+9gV3Z9SgSfbPlGFG/7jI
MZ7TjW3TEzbvw17WMhzr3VFWmLfdOd+BH7glb3XhNrDLKWbeMhV3XtopYN0mQFr01GHRWJ0+pOMU
EHyKOUwAUHdoa6QVsw7sIQufqoqej3ewIUwRBaidyXMYXnYEswTtNxtBfJ3PVH4ob+hoLrZQmMA3
GOIiAVTqOP+6B6Wst07M2/Yz5SqrCs//WOgVHuyfye/yYBZq00Af7E2ERvZoXDcV3FkujmRXIVgS
1cmC/QOJK9qD9lzNOQZ0BW8+viTGnqi7CB3LCEy/GQp90JvPkGsQ+p5cD9hxKkOU8O3/l+bnE8K0
C1ReE5xIaRAakDZM8fgY/osaOs62pojLxlQ8lEN9xUZiZ8gspEldfezI1UOo5tP9E6U5crsRhP6A
eMHsiWdbxLMWPWniOHJ8Ld3E/Ya+y/ce4cZpATs3pz+iipFbK5Unh9oSCNDUJzUG4om7eC1vEJ2o
glLuYCrs94wGmhMu4FzWzk7SxntrYA1nMzK+y5yVrdiLvUEjcCi/CEWFlb+znyI3fGVyXo4Cu90l
fvtHAJeVWzxxDMSjxIMD6lzJT+E59Ume/JmeTmPe7rml/8592aKrQ8ToocLamSkwz/YeShAOSxgm
ryr7elVQrA7mouyG9ncmKcMN+gkq0VVwBwfpAJ3daljs0xFVMqN2WAI35gU11HD/CZ/q8V+kh6fy
nNGFL9jCbWeZ9EyUPacX/3g92bJTBxdGGpLiTA8/VIAWanmftdHnwcFchXOOvdJLx0ancQSPS5a/
RoURCr5ZHVqUru5eZCUGizE34xT4UwX2osMNdCWG+00H2OcHROKwUYwNIdxlwuK4IJsASmUlzIfJ
OhswK+u9Ph5ewRzYSQeD8CVwEBAa2HM8tuhm2txwj8ZczORlowCxXrkXZYbZLH9Slxm0l+eHLOZ7
OymP43MjSqJ4PdhEITejytPlR7riu0mLyQf8pgVACX4X4F8DIk8OqpCxsvcpyPNvQSCCbk1nuwyl
jP5iuBUfZ5E3FqYrOjHdAJKn/Gwj0ED26DwTOVPGEyqoNqPIBZ++hhxXAhzCosmXjsMhP9MP0f8I
Sm0/TM37P50Wk9tlVaHuPncP32z0kFcNGT4w/ltonqAci2HaIKeBsIuduYeBJY+pj41C7KUOEkJK
A9Gqf3g5v1XsSd9FRlNCuPtB65Mi9ixu0OvK3807s5xXa+CIruORv0n/DCEMGhWArF2DN57YG3Nm
6CBqOVX5zWZ3O3nuDhqY7mJQdDwzSVXM24THu03zlff5P7Cgo7BbxFORV1Erzbj+FuVgJGH7s1BF
IihZi5MDZojd5dXedr5FZDmoQr5Zc3oPlSQ/dPoHHL8aAb9M3CpQpeoQVNy8+jJKWTZdQ60pZ6Kx
5MG9UylxovxIqKYR0Rlxl/dL7Pl9ad59Gc+8uArA8/KtRfHxsXE/opyDSXfMg2Ioh+EEb/JbZa0f
R2XtNT7QN3jFv1vEUEdK8l+F7sGwJuhVCUBoCwvBlVjyb3Mz2u05+RNLlFciBxuupNMtAy/+zu5b
U5/IB5ZfVNQSXhBQG3k88AhWjaAHFI6iWFzcpjTQb031l8f8C9cfpBCrdu2n+vd3SNosNs+ZvIoX
IRiaQNRDYujxgmkBs4A/YSstkvuAkVTJlq6rO6+p2lDiddVGDCCsIoRJWwoOcpqRmZUyqbNA/83N
/8bFv6BuNOmVnhb8//zanEUDGtWUiiovbnqkvw9K58DySFKXjuJBEKD7rDAerRgMb7KAHYciqvp1
N1AYxoMrpChwk/N2rjTorMVkI3two17T9KZ09MDYCDq2Y+qkO2DoBT+QlRFfQtGqGNr75y1DkxQi
AL4V50qD6qLZNemvtqX7p511w+4HOnLLOG3L0txYR9SGKSzVR5zQy92TWwbKPLAgEXZ0RW3yJ5CK
kMz5TR8WR3SVXZRtWweHIr/Gzb6LpCIWcJ/VtyHWlMQBMg6aNKndiBbAUrQ7aUcPrURzgLWk4s//
J7PdMIqERjTgXwlA69piN3IPwIe1A5U37LMt70mH1O1gdydQlvnm59xK3YeGlDDFkUO0sXOFirW1
gm9g2g9OR30Vx3HpVcZd3HrXg9GTzochiqLvmgvHv/J8XMwssK4E3AEyzb7ursTrZB6yU6hOj0WQ
n65oGpD9eTzRDitj3cIXfu7Hms/b/+qcUlChoTHc5D2h64vp1SXoVgEdwzAKukWbEDEiR75l3z7/
XxScLO7ABoW5BFwy1UDuENffxYIHCI8Gsa6rz9WJa49jPQcy/HkmbD5cx46SWKt70elPRmLDJ6qU
KAq3dhu9h+6XSGhApmLhe4NPuyopBiNl5tqbjges3i/rzfe7ApRUztmE2M7NJD7hvjpk4zvdUl1W
XPB/2/NqyKNj45SlTIR7Gkqh7G2y4hOjE7LtHtxUg+Wtcg2hVYmn5nAWurBxQLsdm1xVliF7NBWq
0v5OCo7hcR4D0zbz/iUfvHIDqwiBjc5MFLBoyuUgR7bzDDa59BHXr/MpYOz/1AdL+UBK9/e+H5zt
rnsQbdG0Vdp8v6MpqqKI7PPRqFlMXj2+obSI9nH6WI5LXzuSs0x5ZCFGoySC9T/EZ3MbSfXeDQmn
mpm3Lx9q41bNlDudYlkikYKouvl4koVj11ylEZo4UO13w+byFUMXeC3JTly0YX49GmWq+W8RD36g
Y8C1oaZjupR1QPvWinMP6MXE8OMQZgX8W4giv1m+X0Ej5I3gNQdbzOjhD+XMzhM6fbOb64h2k8Xd
VLnkZf89mzUELdQ895eRih5+SPbGDUfwBk2alp0w/NaWridiecHb6znKGxH4krZp7sYEQ9RpWgst
7rZaVn+pzKnO/+6/+cfK4PUw82XL3YRe20xQHcIlD2GzsT+uthc+6droidqIelmmqEQVKppkIN70
awgCHxJf56TNuiA6293ZZ8tmd+K9RXbFGclLzO+5xpc0FIboUsU29TXWd6pXBCWcpfztgmaM36jT
1qy11MywVOul1d8QgMa39IOXiwam1GIdSFVurM7mzPlBudAt13IISKcdTzCWzBgT+SvU1LpTEHh2
UQQXuCWqbX1aJXp0wHc+ldeRFfLbtr8e4z6+nJQY32iyPdj802H3Kq5QVYUrlw+0MmNl93FU4fWB
wToMVB/gCRIX8R+OG5P5XJJb/jqUZwiQ3M6J8jUtl4+IzPRxyNaHFWZsI2ZftpnjB3wnNkkr1T42
mZk4OEwvRVgMQ2LsSSObc3fA1+gNbTd+31g94uYede7kj/rUwLmzNkz2hwoMcbWidW712eAah7qS
BOOCEzy6BmQLzi2b6VK22Ihc6cpwJRJNNXjjwnHrfm1q/dtRGZ1XApcy28R/PYh2ohv5n15m+P2j
zxIhgQDwV9Srz4nH/tpPph0kOaoD2F+1A4NbcTJE/XQHMLh8TCnyytNL04ZM1fWDGpt5t91PBtr/
CHS6gsxvyl3glrqPRPBC8NUwzIESodW5wEsJN+EuZsxBzBD9aL/CcSWg6hapMbF1g5ERrX+//LXQ
7oMw9BU77glF70853DK7OvCmKpmRiKTSizjs5ngwQnulU6bHThCvzjpts3xBT3q4HAhPcvRCjBtE
dGlK0bRsvP6Sw0iM3tawvt8Ue50hVPM6eCKWs2KdSmBhrplfRgY93oawtVuAms7Gudgn8Np2E1Rj
CFIWToa9swztWWfrPDy7hX0wjPsLZh1pHpg1aWXBHpi21LreZBTbIvqiOyOtxagDXPKuBxiOIihs
jcn/qw+JqKnuLXWlwgzAKYHEXwEYb0Tequ2W8Ejb6gX0aCgUh9bC9hUrNdfMpb24HIjjucB3jxvD
s6HkOsLvH0RCn1lZcx5FHLBOAuO0ZE1bw+9W9N0lO9wKQ40kTY6byls4JPp32HNkvBMAVfN7oTyR
84PN+OkpfRRiUWGaCuhCrSizEUCOQJwyvFfg/rtwB5mFgN9+jSp/kI1Bomlf5UHlS87QWTvu3/9A
FZqy0CuWHyKIC2C9dTO7auaCjggZNi3nuAqtcTv9mUChyOOc2WPfOcV73zEcACFfGrFx+xveuILC
1tiCqAZPUqLOyUHvXSr24wJEu5KnQMnq2QxWUcBNkJzJzx+IqwPAqtxpx5DXtVNOhA1SNcxPowFl
kpyFtuMIX66rXxsVcNwHi9TSTOohnxVbq05Lx68dKYQ+Ex0ds+hGqFGh2PMC/WmQds2HAjZqw1CO
8P9PohAfjzGEJk117NCm237jQz76u4xFGCgTmuYaROEr6Di/QQWRnl9R5aJzcH1makWFcJMW/W3H
IkgA/zs0JNvTnVE0go5aUeHfzJg3cVtvm7NEvf4p711SnExu1FvpCA8+GL3ttjNct92t/EUamE1l
K/kpry6czNkjPMgY1gN5t8ZqhaQPnxUiR/8gdt1792Uqu9gh6VtcQqZkWLKcc3z5xc4D6Vy7toJ1
zp8Qf6e9+2PDTio+Qq426Q5wQK6VvI9a0sKjaiEW21ntPl3M0To/da3Z2OuIYlcsDaC8SAmbw/jh
SYQwQx4IoHSqWWi80exmHlRBuRv/UhiQ6L4pfn1s/dSnaA/NFgFZK1dCuVJCKsqPh9bw4GpC0bsi
pKGG7okOtpReUCyfCAC7Tbp8pxuAljZncM7zbhBjhYGQnn2m//icd3VZYeVdn4GuT8d6tvN+FQ/h
9e2bdhGm0JkyEhxTK7dLmiFkiV9CCphJYZGDn394JobJwySVQZTbtcXRvL6EZZVDW7+THsfXB93y
Rrsmh2MyIQXYKPg6pfrZhOfrNMnN3Qw5qi0mtMHOlXzBxTFSToqn4LvoQnoKaGmEPA7N8Rg23lDs
aBaCjtajZgmqowst6LQC82kPXqp3LZP9aaBfRGMZ27zY9aLxm4rZ/cfAi/uowXjdj5DAmV58g24J
omsmk1UXM8JZ3wXupYMj1VWk3WAJhENKKgjEh4JQeI6WAw3dndxxDAcuW/msXaSQ/J/vQwAB4DeB
bp34+PBinjVWcCmbOp5smfLPIt2GpAPA7u5J47r0XtL4jcVG/gk+7feeeCy6vQqFfjXS+36YjzaO
4iN94PXpsplDM37IBe6mGLPr1Yag4PVjzuuqM5Oq0KV6S7byBHvauunvOpd/DPTlTLtN7YC8OR7b
MvG9JAB8xY+OGttfnSTWHmDFbaTlPl3RV8W1ffYE+DDqMIVd9F/r0BtJg9IkiA3VcEXzPWb5AQA9
m2qXi9w0h8GAGUBoERKzZitiCWyg2+rsNwPgOXjqixhFtqpOSxVQrb3hts5LxvBoEhYYv2xNTU/R
r9DzWg9SUGMnlV8sTT3anyrFT+9hY5gNSNvk6+3YU0+BM+enACdXehQX74SpqH7H1rh/vSB+UWhR
SGm79+IueKZc9WpkN9wyWCobNSDA2w9VIq+y3kPCqOr9+5kXjozB1jEKBkdhHoARzRNbl0p587Kd
w/DDD0u14ddA1ANkIjJL9rlW5fwKsb/IJPYoxXwTFB0Y0Nz1F91peA4xFRFJRnYcNpoQ1xpy1QUQ
0ICkxgvzgx/Cck+sbqJfKUF1sw5pNXOszIYv0cLDdWkyoKuyIKaO2SByiKUanjWk5K76iqod3e4g
NYEy1KautNwJIpGY0sUOPcRkGPYDDNMjlTxWFlR/ydA8/wuKWVTLjUftT5shZ/glqVzSPw8My+7Z
YQHTy5JL83LqdAu2gRQrvO0vAIGteKCQcJAjp1y3UNv2rQvgBETJKiYrZlgGySpZYppqcB4PGpc8
FXwc5QJlY+uC5cSLpibF4qKwaodsFizHyE/MDR2xiJujqJq+zjbIlMDKa2xivcBD5I5Rxn+ubcqh
NYkff+SeINHlAV1fykV4PeL5GODjQP11BUzuMEqPsxPZSFDuGUcMwNvIQBXBwPqUG8qp6A6VmsGr
SwE5fxyKKv5b/43Vit/Nn2bQOuk0xXcspBHwI7wY5nYnjpr9dCvEGzx19KHI3rvSLPDqnntdkhfN
NW5vCI4hMhV+kIHXh6773P+k8lmqQe8szZK99rvC6JSVJqlzBs4N52UYidAHhbBVkCqGWgvHbpmW
cEnMMs4pT0PADB76UjivMMrs+XEH2a9+pQS1RHJSe9LdILDPXDTZvz4lnZFXTe78qw6jHP2QpD4G
ipY50jMXg62/tsLhDVrnhr7RLqUZSlnilE25mZnoEEn7KM5zXiJFKVf2bIB/Vei3Eij7LIFhrhIx
D/YFqPcSCQprQIuKEH4+5z4eMDwmJ6Hjx5+JCaXlZw4gF3AKLZ8W/3aKIjS8ksEUr9KWWPdqjY2j
4LqA7CqYU3vqnBtEe2FU8ptw0v2MSrW50XCO9FaDN+6tdi5jMJdSL1c9kMXwSi6R4ifRYMPqH6cj
GL9CxTXfMvpIAyouSmI3anipMPxRvhuxHTW/POh6BgRGrun9abEcTaX8OCKjoSBwpTVKaihDJGjw
x0r/tER5MRmKm+IpBwDlc4v/ZU6IKT7E9uPHQt8eMO/kLHfieuRk6/j92Mm+XAJrETuXZ3qe5+wH
iIC64wFd0ALlMIIGy1BjnfQT6bGwAxgnkGTAWW4pZfQb+faRje1KsYnbPkAOHmAQKPxFUk+FUUbU
le+d3F2+Hlhi18bqruPlidloh605xJ0fxyZ4QrpGM9p1kxRAdvWeGJWLcRXDJEerHd7I+Twk6EdS
2r12xX1Ss9A7MkFekFW6LPPxTJy2TAKPzYm83XS0yKm949hMi4Ebmyqs9gYtUZpSqvxa6og8HqUF
RPNt5hN6pj0tXrwJ44nl1R3qJNaC7g/SUCKFwPEJHuCgLfqMy+F6uilT/89OF0lP5YMYMeI1QnZ+
7B/OiCTISfbocrUyFIyOSbNwlSUxzlwFeDAEdPcbU50n5JcUSOFJZrE0bNOzPFc/vzhKDlZXsNSc
C3BjtL5B/W2+Mg++D1+OA0Xkk+B/C7NLzIYQoTiA6sV3SPJumVJ5W8QzHMtgEMw9qurDK04navaS
RU+zoCt57yo5HJvTzhZWUMnirx0Z5TojCS5f+rcy4vcZrlHXHKM+KKoWKdVGnRCcAXbMoA2h5ExI
Gee6pja2cfC66FCUHOVzLzhBDEegKmb9n9jZdiUycYsv0x5aqiMlBodXM2K4aW678gwJ4kNCBL5z
nMHIweB6FRSVYb2hDqDYJMQhOZHhIdXYWBl90PmE/YQY7NBpSp/wSK57i0WzQkTZJXTgCqCQZwIj
QBwaSTiLw/WzJASjIwkEIs6P5AJ8rOwiClkD3nGy1tsvu2IbbkrhKvwO3d8HYXNuVFC+ce1sbks/
GvVTp0NhnRkCFjhM5Oby459+KSfdwgXquow0AgKRIfIlIcaTTQmfRafitXLXeCoY91Vz7HYZTz5k
xxWseU346agfsingHLcOgd019t3/BeQOTAh+XS14P2s8cLXjeL5wH8E3RsQWcUDUPjD37Gh+9RVY
DNP8NBdiZ2Hth7P4G7xnFy++FAvlD//iqsSDyjg8vzgsSAwAfLkzioRhnuG9mCBvm/xkyrP9aqVm
1sV81vulo2oG2+OD5RRMn88d77iEyLbYiOGBSjwmn9AuBFu+5obL7Gc9/PHWBr5EDOlGaenf0oi1
JJWSPgDqUOSQ1hkYlujYNYlFqRg2WswYsGE5eNcnnUpzlRDHurQDS8t8gVpd1g4EFURhO59TJiVE
FTBrYSM6SZGprE6Cr9ai+Ay1hPhyibUrCk7jblncCY3/3Nz9Fgn6cl5A8Pf+q1znwjtnM8cIfo9t
8VFjYHz3/oNnGum/Q4Wlao9Nzj+POTc/Udet+2+BnwoqK7dA4g06Cn07mAXzuoUFgq9cVUo1gOuS
WzNdw50rzo3DsGWDgAqejrIhyim4XpRhZN6rAiGA5XDU8F/3q3XB64AYx0hLy9DMh+cx3MBGqW3N
3GD/RM0KEsSYQpkIAulOBINVUKo5pSDpSyleTrbbt/127uqMEPv9taGC867XLX8ZjKG7sacRzbbG
ooOe9f3XtK4PXaMSm3hDs20omu+pozodAEDEP+MhQC/jQlMcsrUm8yaRbihoWraXZe275Pyh5fzk
XJjDN352wmkVmZa5RVZosPbxa58gQXPdjdEA+t0SqpwimYxVsXOP9oWC/bGLpcvVq/WgP/O+8Dbm
mWtonwFzRbX4aTS/59IAYRfvdgbeKPaLb1TaFFF8AXm+waY/20PdW7PtS7mD1SaYrLe7gxW20FL4
I2rqhq33XAhgZCjtu3MXyXQjU9bDdi4/9MZIZKcxFPsTydYSVbkA2lOKSLxplBr6Dikma/3f9yW+
GYElWbr6qkqjfju/21dYsDw8SoDWQ64ezJ0ZXaZ5u9WpPYeX7TJCp0WxLznWrMsT6POXLZNlvC1h
TxVRzNBlkK2TvivMX44lfSUAYNdgWlskftfCKvFJPHLYBFBMbhDQZunSgX/uaUIQ9vAU8xDcNgH9
W7PmL55CHsonBquZDFr1s6EVwFqlUF3Hz4oloesCmjG1hb+ngkxhiBc5cliqhy9IOuDs9R6Ykyb4
PCQ4jr1s660b6l/EbqI50yLr4tiy+jAKf3LL3OOJwl3zXAzysuZ0nMPD5v/gpcw2afqK4Zl59Obr
Du1l7d3OiTqtPJsy0J5J0ej/mA8whu21EHmIdzlK5EKx6UncERsV7zYdvCUDMeimwliJiU7czHTO
kYr0+AiHB92V+qXKgSGi9CIakWvHCZzVPzLZcoRstLbVeR65Rga8KIypUz+IUaUrZhJjADWwJOk3
TVNLOox9M20YjecxTailYGWyczDqtleBbU4c98GyeTJXueMPG/PgkzucTwai6PQILspF/F3Me86R
OkNyxP8J6XWpTpPaeO2xR+2PR06tYO2UJ2zmckpR5KkR9xHw9E0Bk1HfSpzQrbKv+vpobz6LDy0Z
B+UhX5V222VYT9xaD4XbRTp9Q51ZhtwcNhh7kCwOEKUjUe4T7nJ8kNmW81h8010wEkEh44wXPr0d
+BhZJ+hF8qIwGWRqBp9XOAjoJCzRzZQkJr5gqIanVCYRwZjv1PKyea6IcSDB8YdLsOMXaFqMH6Hg
2OTA4xMaH6S30Uu34Hi7ItBiA7R/cZMOWfOY6jrPe6j8jggmsaFp83kzLeOp8owaMIHefBHIURUo
As6+U9+xgRF4SzWINiAr0b+d3OJD+6GPuY1KQjpLdBHhLWsUQQCSsWPENOkTAWiym73UT1mZRWgI
uvL8ejaDJB/N6Jtat/+GpjGNWPy/LZDfcxjOuQOHRKF9WEsZLwZ1bLj36tkQjOPN/2HB2u7LKdlA
X0o2IYJWC8WCt1MiVdsRbThOvdSmfXSKu4jZXrwtxJozNCqRlqgqBKmSAEMFr1HxdARjtFJRTyNw
VLZa+NX93PV4uii0keS5sShc7+PXfohJi0BeN2Z6WBbVxKjF3RSLo0/L0xshoDpfJb/Fc+q/f0y8
mFllo3qnD1jp4P/XeNUkFCShuK6mvD8AYY3YjAKvUBxnm9AceRf2krdEFE0/WVwMRpZQ3iKI0q3a
9BsxKDn99M+lXQihXzjYAY6bykeRkm27XGLVyN05g9TiEC5VHprWkuEn3zj9/WYoO+KbgHBZgVZ2
A6kMKzPOpufDb1bEDX7xQOS90/VH8KmNvEDMWBqWBY5Wtnt+SHt/xooWhM7HCI4IxI7GYLr4Wcym
4E7yS2/z9/5ZUsCW27+RAn8Vo9PDG+psX82E9282MGEMxzKuRo+N5LGemJMDPCUXNqjHghISfBXd
0zj5o6yJNyaO8/7Qs5Zp5WF1QDC2E6iNTGkUyAIrjLWPZLLZbp8hGy8u/QINVNsD79NKJUjAta0k
5nvPk2IIWQkIe27vL523i6Za+nxrEJgzXJK12Hrgrh7KhQhwKVHa+gtsPou4aLfqnO03bcSHaEzi
XpqmIQj1Pr3RMnjUh+rsuT6bhFOYAcKrk6GiadXaMLLmUK5TWnpHeAqakLIGmC3A1/S5XAfEO4L1
Y/ULOpsmM20/sx14iRG8xsiZPXnAnDP5qkHEeOCQstQO0QEnOsF+jPmQgdDUKpsh3UGEQPTmOJGE
JOBYLyaJXG02aA4LKKOnk12IKesy/odZ+mz7YSS0w0MZiedt6Ch42OC0rpuX96+W2gPeJdMT6c/3
sCZHb3FKYIwGO5zCSIq3UM1Vz8hlIaPAiTV2D5odA6Foxlwq3g6Y9ZOzx0tBhOq586O9f6mL5hqO
CLYkWUS509xjIoWwwD7zV7XyNrhVF4uwZdfoROQmwaYeMLP/R2f7i1CIkvxaJQnU5Fn8nghJrb/l
ouTdfEZPayFat2YcZTSmIyb+HxdKYfa9kVgjasy+qG1Jy5twW1fdF3vR6j+oKyIOVW0fi5Y9kGU3
HREhEZ3H21E0Gyr+jWr6i+oV3xfqcwrZauaV1S9IIlR7UmlKLzc9SvQ3dB1qQY4hNT7ui0Hnl7Nd
aL21QAh3rxtmFXYWfIeMkqT2xjWhxFz/aU3bZUUhf7Li1pkV/bMM1eQ/k1g81npgsKZraxK5nc5e
/SN/dLjPLXfjbOUoKqsjkp1W8ea0Gh7sV5+HxhBreZXRllyNwcwgIFeKUxrvss6YinPM1Sh7gMCc
6sjqKlUjajvlHcjJqWemEtBf3jq5AMu8YO9Bo9BppH4c3GJBL9/SpawfIlRP2Yvd/VAagJ0eVcgq
SA8CXRrVlmHEtBn41QYCOnPMxu8e5wkA83CzMY8J3rLMTapWlrougxMlT+9goe8YkrhB8Iq/xjpH
whn8sK4S+FpWq+ST0zMXeY6RSJmsxJsJry2y/ERNzRIw4vlELuER/NUklohp6ZQyup0tIIcyj7fr
sqlKd2sXAer7+DyHRYcw0fUDD87TqPvg/M9PeGG+GOqC3G8K+mfARfVgVRp27KFqOOWKLjQZCixp
qMrnS+3kZbo5PPYXsJh6pypkk+v4jQsdQsacU0iaCub9vQsZtCOSAjkQl98gxdPcaJkPvvLwPkzd
SqtxSnjD+PbXJujkNxpjVlCIq9lRshVqSPV8LANRnWoV6FlTtze8/ABic9LqucSZgvxdPb3rI9c9
7+99Fplktz0leQH5sU3kAgMyO4EhrmS3HWynCuPumjCGgRinQ0NlCOnqHpqdlfq8Ogazi/NtXXTR
j1amVNsImf12AlyMK3z+n5KIPFDUzK3+WzjVDtNuU1pQegXfu6N6PHxnuCR7jLKn6KlAitH6hcGp
IXgLDRl98pexVUAVXwLe6Ob77E2ijZPdVNMR62cQ93FlJQUsa+Nwu4SFpz4aAwt87QXEitmJ4uvE
8kGSkKGDZQTXRRCXAPNqqjeL87IcuEEXv7Mg7olIrgwbhl+VvKy16yNzeT9wL2DkbwCQxTfKq/7J
l9maBxbgM0J5Cl/9Odl4HjASLvwXwB3B6S1BXdlpAgO9hhpHnYm1qjaB9Jo2p7lkPwTvDX7twPRS
+0bbT5zwsYKFvKF0bQDbMrEvWoffYrVD5IoVECuP6QeQUPm1NUWQ/2YKwTwhG6PehGqmt3L10TgZ
J1nR5RxQ6V3pB4kDziXq0YBWLR8BxLIAArh5uKrRSh2cokU1K/cfvSHwZ3xAMGaA4mlmXP74XHJU
n7IXo4CjbAFy7Z39xWW2S/ehwg3Olm44tkgT8D8ho5UJD+ZkQW+LUifgCS2INKMlOhjbqm4SCHkE
iSVoRUHe4UWfQU0VVBd9azB4cFAd9gGxrksW/I3ED8qvChmvvxb6uvj8mWCVv73ISyvUFRF4283W
4tNgTYSiGFzKiEd/17BZlwn+lNlWHZvEIQz1vmqg7NdFIh0F4AKle5vNUa7yPUgfGT6afGk5oFyd
Gy4G/Nm0oCzb/x6HhBN9dQND7UgBwZWDCrzdZrP38uWaCg//aG6WPTUTVEsNOqd05GWr/rQpM7bx
GBr+3CTZ2pcEWydHvFDcDjT+Iod7G43FlB9LzC41PFMZ/DqXJEpGZmHMI+NNryYf0qkAfwN07l1l
Po/uwIuAkkhhi/f6QlbEXQdR4HfIoSM2AO/JuuSg0sXovnJ57njGI7AcejrvVhNAqRighnCItVW8
kScTI5HrC7xs2joMG2hruubnc7HyodM6SMQwbng5aYvr31FJZgV4cqCnCfOW0JBY0OHr3ah6cTF1
ha6FrJydPH9lXGe9OzGGWn1Tvqcum5ECN4HsuYHHjTlVfbHvNc1tMEaFwiM8o+gjiqLS/30N4Vc2
arAfrE1nXaWLAfVFaJZfCUQrslOAmNjYQduoQKhfdm+tL9O1vFL+JdSj1ZMi3lKF4djgu05omwKE
drLv+ybDFbp7mdkrSt83Lp7y0gBb98TNx+nB4GgHGkWQCQn4BcQwXKPzIRZV0pN3mVWGqQKni4Ud
09rPiq/tLySbXHu85inveZud0XpIAGsbSWUY9aMkzIseVAIezgGUSTni03MrAXPuPYdl9QAEtYcd
2BHw4KVqeVJTDcGOZAtDLFQIWZQhOhwwpwntbLSXm8Ba7ymlIMlvJ+Fuww1L/hUYJ8n6otDfT5p1
cyuANJ7wUwKtYA0UpVIbmRa+olHPIw22uaopamUAHc25/QK18s9GHXWp6FHuGCPLbfl0ze4Um2O4
u5WOBUtga+WJZYoSLdA9ScyAEYsBYk/H9OyNh6qpD3buRWZ64AGYyHDwwX6yrdp17XJ3vU2DSdX6
28p89Fbtlw/ytuqXbNLUPqzhBDI/uMpS5mx+cCAI5a+YFep2joQCBZuFUnHW4/g0uN/0IpL5hZ1f
E+rU8+k7fvMRSWX122IbbUHbhuQJwChLhctqvWAx2+zumqY9dbxpMR0s4vatAfnWwDj/+bo7008O
Yn7Dee6gDAX0uz3eBpbigykq1/yRAsQTf3B6NDh/W4fnlHiPOm2VkpHzZzADMQldh4yk0n6m5Cow
oJTHHJ6dHqjB20Rz43mpAREzn3eVHvhPGS+YV7JjUa0+p48qmDrX5CSVoWtjCywZl5jGosv0jxEm
APC92HBxs6I9JhjCUpdlalwzFUce96bMc1ayT5OIOZePQCRwJYtwNB1NWlhxDGryfbnYIeleH5/w
Ca8GJcW8ARg4ES0Iu5gmNZazwaZGO36dd6ImOYHJU2G/8LcALgFuwyuXwyT+uqKkGkv0Qi50JeYL
54lgK926K6ahKucVepewjMmDwoFxCn7FuSoNWATvnwUNpix6pUFp4A2/ZK05y+Elbu09RNCHE90N
LsBAcjvRK5DYgSFngnW9xTufZ2THRMwOeDEhvP3H1VAjcvqEdAMZcDv1F47S/NP+qAUsscEb4yA5
fRBqJmJdmDW+6k1wuYOKiBPV4IW2don7MnJdJXXl4rU0gsMj4mx4cgHIrq3DwvNjNqtjcAZDB3o3
eL8R3mWnpU7qz50goN77Aq0eMkD/C6NVSOYpLoTNL6F+KZGlW+WY+buDqhoBZN2SLC+zh/1FeON7
R8F7afaeN5sLjyb0MmhltPbalzvr1EY5dEPulaMhudO9ZX/hJiMDUbQFWRvpMhw6+FA7xmL5maak
n5uKEL5BPd3GMyrdP60DLwkZQTysLTKja36IDqfCKKxG1Xo2c6AX/2uPOfgbEotSbl7BmUPLWJf1
JGhpdnEdzSbY8vtij7T6rMbkuhyF4TQ0+PHXu771TimfjqYlG5riHY5D32fl4bCUDlsgf1G7QhIv
UwDpBqA6Q0v83bjXhMzxUyUnY94FuYCWHDhRDY4GVT7ldm9Pr0di5ehyx+0fM3vArFCeBBHE2N4X
yMxTgpPDvXrk1gALQOub4bLceJRC+gGW7CQQxGaRmb6hQjT/VrhC2+V/qCJgKtRyv8bsG4BahdLo
GfmfYODP/k8jByknOxv6NDf+02HMIAqSkH6/QdSAS/IvfgXdL/6ZqUivXSK88oTmM+r62uHaqyxq
i+2VM87GsJbiFsDn5YojQhDVZJHek7umlJk37rfBURQwpcN3zolIXPcYg3cd0HEx8hOON0kAzszV
epuiFwJBqnWt/M8J5Rr7BVJgZEf3R+psMp/Yydfps2oQZsbgkoKTobLCz+GTtBJm/MgJm4nKKw27
ZAK9OkMvg6rIepvvgRXyGKU7ck10TNxBlmbLz70J/1tKHLHewzIVfGTG9TpSZOx4ljIadjz91iFu
4ijLiSoB0CN5/EroG8epUelIZUOUe/BEOljyrfgxLPVJEO8Q1mT5G51K5drRWAO59s8h4KQR3m8E
CBlQ1Aodp0G74PHItsjOgpipJVrmGiWEBDjkJFA4IHgTUz5s3QwPvDbwaJgG4LS2xNXu347BFCCv
AsassZvUzb6LP/9WQN4SoQlxN0Nu8b0gF327SbXR3jpsp3Mdqyp7EFrqeWlfg4uMoyeI+jx5T63b
B3Fd/ENVkesDKxgAIwBFM8nXIQPiJPddb0MoJbPzdmmE4ETrXHWC3aNrzhSFtkZi70asx/KzGpsm
UNIjUAL2CzuutXgP/q/iguh7/XN9JTEyBsMfezCz+s4NRvmlPWOuyDWG7j2mblIQSxIXyXZFv/Lk
Z844lwzABrHpzUP4buuEeveANTNMKwnXKPxf5WSL/8hZyFMAMGOLfTdg33Yq2vU2m4qCvxXIBnOH
zdz+UGnbHzcNDOIgdA908wPZTJBuac8qv7AxrKOFgTJxO9w9yrqGNXVlFfPBHOJYATBw2RR9lGnk
kDDGrumrSqr2y3m7Zf4wiUwYO2Ofqw+zxMq+N7mOfLvajqo7TNRE+B8ax6+TgwPOv5nm2u6gORj+
DW99o5fgp0SXtrthiGpUAPUle0en+Sf+ncF7JEMt1fJw3Vwd2Q1vHonulCTJoEeS0IvAL1/6JjQX
Mz4lKcE5QKUfQK36uZc/ebcrQU7cyl8GNI4rbKkT2+ZDWml4crK05TvoDUUzZem4PJ4n8jCD8wbI
QFY959dWguOm/a2fixJqd8vpFfO+l+X4wvzUiB1QXWozMAPBA/MLBLjGsFwXnZoINGUhFRNR+kBZ
s7Ws+nQwhVETUG6zdNiQeVl/umm2Te+pc6yTmYxsXZcI/zbvcbuUry1dgABWOMHM2nlFBIB043NE
GkBZZoqPI2KtJGWCoOhdo8Y+cnGFfpEymH3nD7tYgN5a0uk+lSedOZMIRysZ7JWoGyqX5w5kpNeG
79rWxBTqv/C/tFQFPxXyp8ij6ZB2Kc/CZOAj2UDWI+D9xJXqNnFNnU1JVNDlsPS7T58L+Ulb4cuc
EcPViIWpUCprJPXsG5r8dmdGVCAzhwmIT+PKG/QILZOBhiEjBfRldottROdyocZnwrtKfZvb71vj
8T2P76YddLYOE4SImnV3ZQm8IB8MGZigQPkHfTbzP6V7pTq7e/v8Lp4LP+JBfbPSBV/4af82GIMd
V6CAGQVrKSfs03QTEfv6UL8hFSHrl1i1ul117hor05Notp28FddQU3WqImKay2DAFz1F7NBI/ehZ
XnfzZcVHXxwoVdQ+65jGi17p91BFgVPkjlptmtvaDcnX1yHxKzj1YbaQOes/liQl4VzO8y2m5AQH
4fHpvaGnKSGZKiUJqsdwpWxYF2+sBXgcHLvYO3vqDF3vqZ2NzrS9nRu7RmgH26lUwvsMt7fjMhFL
qYT+rgeVQAQ9aYA9fZ89DHZbE+2G7FPzelYFBr0/9kSUSVSQb1dkeZHj+7T1u/l89UgfHuYcHf+j
37ZGDEMOgugZmzmtI1lSas2rxsDGs+b0cMAIBxhXoeVAmJRAuMQw1hA7SqY3vmKmwvi/uVVarrlr
Da5Gj0A8tBodZQX+Wyh3yoDJVzWjTmzgKH4vA/7zaefp5ZDdE+DkbtDdARtNdQftE+cuMZqwPRp8
AySL8jDEZf6B31uvB73kaArYwJ///2kJO0Zr/AyHkUU76WoCbZEL7+thXd2v0q9rsDKrdserqrYi
HG+V7GJ4pg4Eq8wlubxNM1GQPrOXB4IbiI8Rab3kDt68GIsLYg4M6sAodQUPmYEAMTuCVhXngM8t
r3y95PuoXCSV3Zt9DXqFa2JOn3S4MLBmFuvwZd7byxntD4VO6oPzSzk+0hynW4MYzwhKJHtgwoVN
U1zWi9wIltiVyYlEZYUyHsZJ1RiPkecjpcQqxohC2hMirNLBfPYS9BJsz9WdhHo12H4N6ntNZWSx
yodNPdpVTJJjGpnz9y1zjAzZX2+HwyKjhsqOuoZYKDT7geQ2bAZx91kI+/O156FV258Ol6Tcqqgg
p9c7GY2d6LCfxlzhwkN8lkWVoZ1IDrm97iZdiy4i2wy8YT48O5mRPur5P66Lac5IJwMkvERGzWrr
6AkfWjKOlrInH/Jo7mw1/NZIdApCIHN4r4iples/5egK8uWSN5ad33Oc0fXJYHBs6ezIFJKbqHbN
WWpW7+rTT0YsMKRY/YrTKL5Ienqy1d4/jzaJVupZhgROYVP3QB447iCWuTq41AxdxVT6i8uvDGyp
D2W9bS+K9lKae0ZlQFRvRel6/jVKx1P0Ry6TgCUx+HiGfq3khRITrzNXkNBzzZdyVVNxylmNdDYi
wEfFOxEt9Pl9RUAb6x5ogQRq3qCZ8e6Mz83WAj+GMYKWuq5lloBhbITNdEXrVoBNcFgl0zDODeHC
mhG2lHaQrKUobppCPPE13Jg4Wy6BtjwxDiDxopQYKBas+qLnJVbHSZlPEkJZeQKdMCXvaikukiP9
wDJlP+LqRolOO+U2S427q1JxL8VSStPtQVXv3t1mSmdebCZCo0A73KIM+v8j41ev8UUcjelD6Xgl
VcxfjxKVsWpd5DN808HsMke4iqHCBli7/rJtpSU7WGkOKPBjOO15uphnGiTB0Ta9x1aJ9iIzsNR/
Egg9zXq0xVH4Gt6AgSRU8wq8f/5n88YKaFGIu7n7FE9qQ48ddY9twdhQfiJPbHhEZ7VaOoQKJqmP
dWyT4SVPahwFUUEHAdEvFyJlVH7CwUeTRweuoeBbOWiYzwYQu2qYFMCnrQyULO3nXxugipWhN6Oo
e3fd/AmxQvd6Eq/qJTNIgRnadCdw6Ko7ZpIFeOiV1cLAJ2xJgyroLuS4aBLPAdYN8awryDe5Hmiv
OwmcQQUtYKL2sa2ldB+hFnZWtoN3NM+jyffDs83A7CMAHCeDoyOluCiSRqtnEdMPR31e6iFrGpWA
dH6DvtIQYxct3mZDfC0KDXFsyb+4PPKqR+mdTFlY7TT2UjiEz3fUotUa+mXz+3ZzNTzxri2PbmbY
zPdx9pK2HYlBSyVn9tOxNS/sROhIl6MvOdsPc+bjN6ugl4b4Srhqb/Wpbwc4UZNh+GSzIXNjZgMi
xaMYcRdq4WzZ0bmqgwWNBEhlepDh5nAvJhRKbHZmgKb5qWXfPDh1lOldz7DcgEJac2Eto4ciuP8z
7a0rWMyEd4bxGdGh3tq6Pn1VfZHWoyo1jj+Hv9m2lX5M7bxPYnvR4pPD7oaHcvKY5/j1YPQJobDh
v5u7EhS7WHa6B5z2W7AX5EVTqYgvYTZw0/vWmNUPAuPaEjavCGCZ1lzaOwc8/fAFpAR7Djz+hLJI
L1YyW5tOrr+oEagUDfgBfe11SR686JD1Z+TyaYLcTmYp/Jqx+42/wgErlzSHd+IjESbLvIaR/LU4
OmLV5TesF9Dhb9OEh5uSt+LNUlWWIUTTPimwsreEVmoDrNxUwrx7OesEkJg6Bp3pTQknqtTvg/5w
x9ZMrufuTST7ggvQGSanrfjkObwN1UDf0nNwl7jEq9Wr/jLKk66OSxr+Vqy6EjqZ7C4h3y3eim07
qBZX+cd/dS3D9UzLjPi1Jlk3thxdzolq0QQ7oSUzaBVgZhdOiQoXCFtIEnvFan4L6QmPyT3fcgCb
IHlrG6heL8tLYWZx0y4elmNm6ldZc5Y5BzklwH9O9HaFRuB1/HHnglKXZIZQz+ztVR+hCoin3lun
JXt0b+XPBXhrIl+lzdl2wEXXauxIAuqpSqjQRQEj14P9RG0JnHx7LB3g23raD4TaiW0I7w0QCtyY
W7Z6KfPpYFhL+61A2HsnuCBW8j4xQsELvXm43bpVh/g3Oich6N7A7hqPe2t0KT5QZnY8o1I6pqkV
ibNX1eHisiMR19QR0HCIB03a9/uSm5qgOWP9bFgsfQgZQYse4wZRA/TychcNRJWRXAfz+Bzh6Nty
gieRTnOEE+ZK4CRnbUMts79vsGcIIWw6EOF73/uaydKG3aNN05nrFQONjADyTp9VfkrLiFjKAHtf
cKkRYAC0u5UPhHVwg9ctUQp3lhGc0NakUKpIbxNy+62s03pzdVckzP6TSYvvh5lV5mgwU7V3kyz7
54TIoXdqRvfDWO/l6NeE9CP/jYlyhzKTnI4c07w3Xsn/rJd0ZGemPQ/rAwtuDDC9IjcXGw8OtLQG
Rli0Y1boi0TYk7f93vkG6zUA0RLT/hnWDhjJ5flZFY2hCEfd99J0GLE9CpXbMKKOxQ+cz7yuLqJN
99IleUdhpCWweg2qeQES51MiuMHAgbBMDQAZv4750F6zj2+Eoy8X3RespDse52clXaMLRKUjpLXt
B3k+ga6Ha1ikuYAy+ZniZiaJohB52P9XNZSjYWkANmPlUBMyhXMo5LggyCD0f5YNsXtOjZm1ivjg
2DmLozRZAXT3JCFYEvd2c9GwMv/VSVVHR54mjUJ5ER2X6DmukwrVUE4iLEBD+FvBG7BhJXYBh+dk
5a3BYT+cPhmzq2ZhrVdHFbkc+4qWzl9ynKNLj7uZOEOwLDqQDODkmn6y6RGDRSANMtqSSYolRlAf
5dchwXbiz66VdRBeKa13keWLGWQYGLgkxYxenr0YOPQ9y6ZHRUsmeoCsbECTiQN6HIziuWbZVRzF
ic04yJjklDZLfIGkN0Y19pDSgNak2qhVMoSAa2SvOBfLtSaJO0DOw0asuhf27SamlZxI0eNizZd0
dBV9IKC2P0m4kYsqztlXyVhQQreOk/br3n/AvYTmf66avys+HlnGumhNK096lPhd0qz7iP13TfhY
Hbhj13FlYPs+8GyGVpz9d+GnjcaxNlgKYrA+CD+LwxyoP+fsqB0YLDWA15A9XF4AIRqmp+axnLVl
K64FyAabPlu/8mWwRhfWAsvsySU+DIOfWujQXROW3hxrAttMddhDqypHvoGVjpZqJkPgIWJCGQsZ
jaRPmK2BuN+mGWcrFrMoaifQh2obhSASSC+H1T6fidD/oXae30hA7xlq8gd7dRp3YDmMlERFQQcP
dqPhIJ14OxJ6C5L4t7WIzd+YrLH8Gcq5xYVKY7xkQHLk92DAVFzmOoVcBu4AGl49/FGIfTWTIN+x
jftqiIP6M7bJYKoIrJkFYTrs7/bQ3pYaGTGOFU08MnpHWN3v77/IOOCf02KW+0YPu7nU6mpNRXAG
5NNqbc5hAJfdTVUXjONKE8vQbQcoQGnVgbyP4NC3fNasGiedhMUS/v1FLS5XkNzUVSaBcDh6i8Yd
qfKchVpymMEaarFS4SLdqFDVgbuli6RA31oxDYvY5FgaASyRPQa3XAzRHwwWHN9Wbj3sm9jIAkZh
FbAXWCDHkFgjnhHK7DVqxaPLBNSBG44bunqBiHoO91s57z+HIzBrb4eCtOTygvAtSZMOW2EAVbYM
q5dxCU1/fgn1xluoj/pxQtm9ZErXmlc5++OaFoEAfqz/P+I3eORqu7y7CWz52JsHWqwiBu9+NVbx
t4kWGl/CpurwDbLC2M2fd5ZfVBMs9UtojkXIo0YTDfBa/H/SpNIdccE1nf1rZu2pmqZYVltRvXHJ
vMLgEXlDvmh6PZt8WjvaNp5Eb1mK4sz/hMiq/2+0M9lo0zvaEMZemAIB28E+p69CbxPH1LepUWMI
FfGBXkmGfMHWo9CZmTPca46UJNoWYoELtapiiOfZAtzQV8iiAYxYjo0MtDR+2dVqHcRz943WBNdG
kKnn8Tv8OgJ8TUtGOfRAu4YjQgFGozn9P5Nh3dFVcXGkQKEiza++hesVWZQzVE4eDb1/qmi50M4/
ze4KOUXOXM9zHXvliNQEPvWd/LhUhhsH/zwI6tFwswLNdZ01gScr47DfmxR9vXR2Pi6EntWdLgAq
57NVFSAW/ghxPNWRX8Rny5tQyYBgGG+XrG4S7veCgF3IblllJ67Wm6dnUS4BvVFx47uyrRBbafFw
DMOCM1fc2qlczN/Hnw0cd0v6mkyMr6fjhR3DV67cQHvGoRdKhg8VLD0EfsP1S6rMKwmL57B7IFTW
VGmv0Ua+RznBQtjlDs3KaYF/C3KpGBrS8ilyEAxmQGKhylK3htqV/IzHZEYLSze3/J8SiAUIOAbk
Wf7yhx2MnZul+ggzETNOh1RKYXgkDgDnmNjur5qIdedTZgeFcphe2BzML5HoeH90xfFsIXFd3NsO
RrkmrAyvFF8OA8Fx2UP4umZZ02+IDjfw04utortmydqHA3Zf1ykkyP9RV8/Qiy7nKxtcQW6GyFMY
zSYR4HWoV+aXi+hw5ZgRH2RdG3MUy/qM+nwa1XiLw1+c5YU0fkBZv/oAWRYU8yAVJgkylfRndfFh
AEvnMj8s5cg8GmCFjht22LxN3VRPEGjCq+0/b6p4awkHY4hgbJLlDdbQJ2YcVr0UZlFk6AcTYx8a
YDl+rrw791Kv/QsXxxRvZCe5UNnp1GkjzOzaWX9dnwtdwbeCytW8mHcXhARNS8HrdbD2W+blNSOx
YXVYKRB5gSLWVepSKiRIsezLNR8OdMiDillqWvGc7J0LAS0KQOhFp7UySD2Lm7S2la4EeRaZPhO/
3quJgHNcFf7phaHTB8oksR2N65uFc+ZC2YmX4l1jruFIKZTGTn+UFY2LDisEkk29SAzDeIAgMDXO
uJ1FojQuqtdzcIaIAbW6cXWqPw3kqsv5lkdkptmzKhmZa0e9Ct27PdJ+OmohBGQm5N3h8xhlhVLt
Rog9MwBdEW3OjflFm3F2pvqgEEXzwOxEKYVTJ1nFE1E1F+679vAoOOo7XFpmX2IHoQIuoVLnBmx4
FPjlHVcRJVbfzCpTVZru83Yp6RIDCt+g230rR7j7XEWCHq8K4/wvS436R9twY86aiFAu/Ep9YVqf
v0GJn3O4YMRBYeqjmKkNifS98N4ysHCEmO109HFbsi+MWeWKCNvgli7ZlVcs3FbJ5tDr5WNK0FRV
oc4I8w+jDCcZyVHNjDO8fdfZxOEJvatrXiej/uVM4p8K/BPE5scAhWDxllTbPbq75SFjQsKuZyeg
y4kF+w2U/4a9/yLP45oX6aENvNcePB29IYyWYsDyjKBqUKWrO+4pdxjrURBjnFXiHCdeQmLk3A1H
2nlPxF3ltmsKI+re/zkWzB5KUUp/vXaepZWIF9Pn3MEUdlRs5HD2A/I0l7UnCsKKK4HSZVmVb6h+
c/CxXal7hYKY4eCtyXyCTqPBP49ahY7Dy9GOCXzRQv07fNIomneBTM7iwoA7LfkUOgXV3ueoBE91
rqCrAXkFf+Wd7+5UMh2BraY3Orpa3+kAxZr8i09Kyd2eHOClpCNhlDv52dYQCtAQHA25No5JROEL
D9/pjYcF0qGn2QhOSwFgUUfXQdImHJs34KayYDSD06FHRy61mn+eL4+FF1FsDra/+x+zppXMyobF
vHBtvXt/QtXUxFpS8i/XHfLRusXZ4ypzUiyVB48YmxfUAHwneYM5QwjeAztv9uxEVX5xCRuuToXN
a0M6vR20F4zEV7oN9CBzyjB1slUrQcJSToledhiiI/8OFhPwe4VPfs0t9qHsGMwbufo94IMFtx4L
Ff6SExttZ8fHysXqm7yx+4E7Q1BJWufxeKqFazM3D792b18BZd1oFycf0D0zsscpBqUEUwDa9jrt
A2cgvHsMYs4H6TWAW2zU0oLOuJYCw6LtlBcghwZP5F1I6IRvnt+NdO8jGoei1aaPkZzEAdQQtfN4
lEOf2TfYRTajhr9HmgGd2WrMYZDq8bpWjEP8vDHh7qzvhi2u1RFxbzXtI9mvweAgATYiowidNsy2
8ATpS+l/42LhkbgokPZFfmuM42dFKXwa7RC3lsowTfnn+ZPjCy5+FB3DX32phXba+krizOIVx8M+
LEQd4ylfiiNKv6Qwha2qa0tSvM+2a7g8C2Ne8cfQhCSMiGvWnNg0z5pgdIBNIPO4WHki/EsmEv8S
YtjiC/0ynWjw6ReR/35vy6xXTuSJdFX5XQ3njdcXkGff1V0V3+ivgfj8RAZ4mix61d0C5IEKBmvo
b4ZqW7m+GsoW0mA3dQQbf/shyUxaW+d5QmQIzxJhQHP/GgjxtzD/CsZY007W4CmKaXpy/HZHHxWZ
pGldSr24pYiNkcTLeXkA3i2yboZ6cTIhhtJ3U/PklLom5Cg/4D6onukzmXCtRsb0h+phPNf74z/A
OiL0gCePlZkeiKa1bI39rAwrne4E476Vr7Se7mZz2q90qf1q5JlTI32BRKW8EtvnUlxUehNwblh4
uedAXN1K9oSnIlLtIVy2cQKjG5QiBSsoqf4eDRA2u+Z4TfIkaIHlW3125Cjm86ysm5vpbQ2DdT52
lmak7MLz1uUaIbCHuIIqsoi6pqPUOkrO5m+ShPnmQNkAyDlRfNqpzWiiPbqrCqNY/4UmF4jkS8IW
xWDsfUY25gFXGCeqsZzJxg7XMC46E6OZ9KulP25CNOzkw+pff1mWZtFQUXFONOLpdXHwCMf4DSs6
dNSWlhn1U/XtbCpjdq80CoH70rQH5xU+F4Y3BD/dGP/hWHgLyeNSTlJ/0X0oGtGbelj0vKB4Tr7O
jjl5IIQ8tTvoj+spwD35KrhTeYwXDCxU68FlifbTwoSw4SDSU0mFzejXhdBFGWhM/3xMVaj4AQlk
I550nI6zHyM/FBRKUSRlWlAub3fmpuYuS1EfunIVcZvTbm1HWHJDz3EqFqdtPz6FVzjo1Awzw04v
sYIXWz0FdDf0HOEZNUegIe2eKV1QnWTtffM1nuIgplYh1tCNUfPh9yoB4uCRFokaoY3ZGC1fHRuT
qPl9H8LjBO+E1C7aW/84mRQrrP5vgeqn7cJ5uj3YjoOhuYW8LtW8sqRum4mPFuG4t+grLRP6/Lva
vpS+4pTSYzNS9QyxluNHPU3Yz2rux7y/0D3M6JFooq4eT1UgwCtf5Xde7Z7EA4DAHs6gMhy9TCnG
UGtldnhc0AlNzaZpUnHVqZ1pBWlXJM9T8S8WVvjWX2HAOHpp/jIR3tZzrlupW5gxiTGEEj2dmTXT
8+nU2k//Ymg9UyEBgVL9WaDq76oqFGN7OfxjnHRtBkhjESU+FrpKaowVtXId6sDvhBXu6HSQtQA1
Fj0wwUpy4H/lkenPBbu+c9lfvZRvAscuI20Kia6BMEuDlnhtuJaj40ecj2vGf0xq7P67eeAv+IM8
JOyVFYp2yW1wzixmWU/AEZE1cdHMpUMS7ZSlaw+qoGBTtilNUjcYGg4C3NvrFxT1Gq9cSioC2Fvx
tfWOsvlsAcx0AparHrBor/Kkws7VKY2xwM9sxI+osy6zWCBLNkJAdWZfr28xP5vmwelJIoFoUFzE
9NHQ11Q/PTPiVzBUDosC/6nzSzxaO59M/Ul0KTXURLnv2uqbfOsA7B/jUGRsDEux3n8MafaX/32W
dOaP8+5Ox8l7XGIeZ814D9Cf5pE71GZRYaZqfxjvpA6VU8GLNbzGdWJOOMnHyuz2pf0Tg2l84F7z
Yan5EuJLay7q1wJIMf3z7VNDaKytjYWySowYHy6bBHgfMfnPOFK7jQwuRSIQ/6j/FVT9NVfhTST6
1uBAoj4kzoQZoYe/fuTHxLQtoXP7D0yM4PwbCpvg283IwWTl9STxVNp/7bnr5MJobsYHcwCCzmxf
uAjzIlsfb0P0bkmJivtAWT3U6jAqXuKS3LYe7Imspz5uC3rMU1PWzR1Xh09XocccpxNGgRtL4PiI
pcnn7euAr9QCjohiN6hK6cSfQr1J0wFbre4y9lFuZHzgNgQt35LiVepF4/AzlFhlfMIEApATRGi8
7GNrqM5jnR2MTODVkuAQuWt5CwcucyYMEO5jvEp6cj8KN6+KpC6etSo/NcmAfBfJzDClwlAVQpBS
9voIe2WXyU4Ei7oOsQ6iAktgwaR60++vZRyfccl5Jd/pQFmAucG7G5aoIOdaRZAc08DDvrODTwiW
uU9zuuwrc08/2UkZVyCAxu3LVAxWihb0Yyd3bDBhjLOCpKPGWp2Oit16au1BQ97N70OXTcJm4Gy4
BF+nksgTgTCA1mKB4ZmOO6FWJSRXppDLB+z1VDu8a9eiiFlyRxlPH3Imw7lBCMTZVPEBVQeVybaG
aeGqKgMDb8Q8zlKtbr/xhYwz03B8w/0IrZxofpB0DLKu6ouTghpAhxVImsS2+9SvP0+Ab/hb/i2e
IJhqugGpTlvvPaC9PplcqHBrRFl80vQBgzF0dfqjQC5XMbdNFnRPvboZyMoSzU2X5Yi5yI3xSEzQ
k3vJChm7Bwtf7dnGEdzDZw5JpQQfOV+PVd6OTDBwBffhkTIAK/kMWIiYZnaJORJVQDbtbxzeBItk
D+R49aZyNRx5PLWV4HQXkIP14m/xOktr0+aVFpxKdFx7P0mV8VQo0HWSIemMOQ1X02Ev/Cg8vw2t
6GgPH6DqXL1XoYwoR0zUQzuWyMlEViKrSgmOV86cW6Rs2PC2qcVkUEN4hIbM0TdzuvMCpUa6QMTD
0niazXIOZRkDzFkX+7Hh6WLnqszAQ7kbfuQfHBDdUWiGYVMRDU64d0heFae2DOKsqpwwwDHpPVOZ
bvdaOVEGlinsHvnXJtwG8ImCaaRFDMfEpQrDN+6B0TiCAsT615VX/tomkaT6mNz1Y3HpZk+YqF/t
/ZGCeouTb6rNHOV2hhwRZS3iSBChRvMFdccS271MLm3+ETikHdrBvGYane5o/AEEucCE94tdEwKA
GAO34aj/hJz46VWcbyAE2wqL5t+YQ0TKpD7w4IMvMWD09gUorXaQ/+7XUP7Aar7T7scgGOUbfQS5
5AF+8oj6LDCzu6sZstYVCfui+RhaI+B2jUi/PSSBGZSnZAeYzvNX/q96LEFFy1Z9dvIkY4Jk+BJ6
0MwxxUy2ediVUJTsKAdpilOAbMhOktRmXt7P3iN8l6zH6q+zOluh8uwnR0hFVtcfOiKhzaRNltZg
tLMCeknPGcncSJ8d6HMdtQcKFFef0XkcspS+42m6x+4JRP2MNZlFoTiSaONx2AsKGV0/IMcIKXXF
Y+S5x4ogaZ08xXh9XmjCBriwgPY08+kS1ahNCRGp0fIF5yCCqqxqGe8IFcGHlNjL2Rh93vI8Oygy
9isZptHmXVx2pO3NBCc5PkPUfy8IDJxu3cZcl8PD7D9YmThm6ISdEQ9atIYpH75IJVQo24VerKVS
aI459y7XbJ/04+8wl4ojhNaDZWnFJphSq3/QwJfmVS9n4LGrJVMQjbricIRopS5pvqiOh5naX8Y7
NSb0Jy0eFh92bw+1b7nkZHd8J/pQONc1+14jx/J0fBRdoBILQ0BtPCsTqUGi5v+x0mljk70Ihp/b
VvsgK2t2kudDpweVxoU92lkcMwHVKPQPfRxop3g0jMnnRnCeCyxrp2A1/IloZtxG0tjA9N7Myy2s
pJmIHPi6We1iaHmaaKxReWrjPsG6iquFJzfqQsbuR3MhP1/wtkYJIOCcQDOPONeik9dUm6QlymHx
gWxYvlT9iyZPP7jtjCEZfp/hEG/hu31QxwfW19FFKOQa9VAlV0MVuxX2Z3Uvs0XB9paaspOPdYKD
eg4D1jAXhaAXKfvfSoOuU5HW/CBgLyht57X5Rx7eiBn5Dc8AXUywZiZ4dwxnuKTig3ZqZjqXPmsW
0jQx3ObHQmX7xLEcN7e70Bc+MefUkqjgfE/ZyGnmDaXwgm+mIawv5+hPW6qQoJxqM6TIVdjtzgxv
dmJWUocjA+kDWJfFBrym9+yIPtWQkepgolk/JOtzD9KTjc/mTX3SFPu1P4Hj3RI6FPpZKbkgTHzu
V9fe13fhvShHIw5s3klKAQY8nu09n3HC+0Cl6auVtQb//v0l0iWOqV/E4q0jlfApjXwpYUDiDrAc
K6DP8jFQR5eYmtm6TYeo9vzQMfKKT9l6jmjmZg9EWk4viC7fU7S+jaBQK2uwHzoqTG1SA7nS3omv
qzr9iZ7QvEGnt1thGwoXeTzkHwGKVoXuHOfgF7H6l/MUKPcNXzrU3042tlBRItS6i1Wi2suyecHL
MZavFOHw4v3CltgXxgB4n7ZoMPC41QvacG4eWocvFdP1knGz5q1wDthimalxiKXsnUJ8dY2EM26x
0tr704+H9vd96ZEv6+2fKRaadNEVoGX3Zmx1kvGKZOFTQZOvdof6Afo5WnIUmtNrU3MI2A8zGARs
eubzopJ8EeI5MyeLjPn++Pwossh08Z9+rHsCyRcgP3vyNXKqPnR/jgABBezWK3gTWbaFq4YXzj9V
IOnHq7k7/QimQCsyQJLhi7kILW2xXffWQQ0Lt7WnCUSFBmOTfQnC/iCJlupptpy04Wu099oGOptM
B5qM4Au8+gxJp2NbToi1O1LxuRNSvF3wiRSX6zewIyVYXhmkfJOBJocCA8a/StUNE95wo7DcMIn/
fYgbsNBVeAiyLWi8GNZ+MCBcvPG5JINyFEeFGiTPJEbYsan6I7WkLZwXgw/qWZN5eBLnfUAWmA4o
hNAH5uJgdPSw58nEEHXNPLb8elBz5PhI6E74Nc4811ORIJwFgFAM+gAZZZbC2qMOhtVSI1krKcol
T2LXE/HKNqRzm1JaRwghl5MzzsnjyDg7LBho4VEwMUWFuiAyX9dXOaiPAFK5Gxjbxe1etVCZv9XN
SfinQu+B7g2cLAswjPV10BdQckYlzSKUZFvNBQV+JJjBBoYyES9jMDbwUyOPqZIvVqJaziPgjgV8
Wda/Ds9Y2M2TEISDyRXdK+MN/J8MUAC1nPYLR3Zhk5pLJBuxobrvshoGBOm8yEnRzNR2OO9XNidR
r+iMY69eG9uUW9T7anKUpA8m1KnhLGkYjfp0F9r1fp+SsfpzGErvtnIUv71IcQMb/YHJJQnRsZXv
NyOiVVvkbwUGSQPd4MR0aHWiEQG9Jkj48z3SxNwi5tmy6cqkDNLkOFAl24jeVQERi2qt5qua/Imh
WWjrCH3S/qK3vQMVcFsUHDJ8QUnZkwNJIkiTbmPlLBi9wACZgRagG8BRGBAjTqBqH0jNmeDnYjCH
qxdiroEiTsqSf+KnHbfd50XKXOO3a9GJ7A0kGNrb9gPOh5n4/IEUv9Y79OAPqj2kyg9RmUGb2RDk
rF+CJxTVipDwT76AnHgSZ8VlXmv0+VE59enlyA2/h1QzBZp4G7tmuDnFkHI03V5ragthbNSWCkhX
A389VMdtI2yEclS0MwZ8r3koUxTMgv3p4xzPdBznA7ovvXyFwbIGzKvDzK1uK6uq/vahXIlhjGPL
3sAWqwKzSAReIYeYw5q4QqVR9JAduqLEO5bH4RCqL2diQ1SIl7VRjl5kd2NJE+Ibg3B/kdKiGE0B
HQGQHA7O3Unw0hASwK0VfFWT0f36L5CwGOFj/7iGuhwFxw3IchwBBpPgy68Sm2SCBiXqoevnjdoh
DQTFhsF3Xp5dzZJ7ShR0eCukKudWvkUTNdGj8pTMeWQjC1kF3q8CdGGMXwHTn1dcAE7kE5MaH/G4
qe3C4t/X1Ofy/Toj5+DDir4johLM6xWHAffP/EElBbvsRd/tI4yde1Y8iSDRYnTWW3V0JnSRuxuo
wi+KbtaAm3iuT2B+wsQbwEwaiGDJU/tIf2q9z11tWqqDaNVmEEn40/ZA+cSJ85oZ8GeGaY7meO7L
Q7xFCdI+70EEq17K2JYMmRp/HcjwZZDALbmaGoezRHpLgrwlpeAO3tAuoo+oQRZ/gg2wz72eurKn
hj4VhtWkoOD+xao664GVynTUkY1qAQcKQ37T2dLz8ujYoBugvsN4WTdP2xdNkw+cGGtOekvp/eN+
dINS4r0sh3qhI1Ro1H8+80+55sbxBNCAoQBiOKKgV2W9lH0PbiGiDx7/Xqyi9soDk/MKCT+6uqZT
7VkAtU3gDC0vVxWzQVtkx+lCSjPP2/4nAlhtWjx7HUA2lXgqilD4UlwTU7S7Yv9B4lor9X2nZLR5
KXapMkKC5I80spW6PmmyoaGpJueDgEuM1ApUV7OxF7prEJEbNiVBU4EigjeYdL2j8goOQW2iOJVv
Fe3Jweg6xCVLQY9B0vuVcWmvrKYgQ5O9Ql9KGX3muOf+OOW25HZxTCmbgliJ7JZioKCTofLQRofV
94tLWR3l8/ppco4i7Q89jrU9th6Kd/JvBddbO9KfIYVmmaLQXv+zHaweYs4uiIyo4hOCAm6DlsKf
ksL2Xm1dnH51UtvzlmKe8WOyi3kGpb7dKhRENu9nc5kbUJXj4nMvH1rB2XZ3Zp+UKso1FnJWDWRH
6/ioEQePJvYhFRuYFd+ferhTACkuQX56FLk038Y+j1wANPah5w65r/3E5NBxzfsUeSfHrKGTOAPO
7v+2VXlZZVdyNCAQ2WNzBdkBvHz3kg8MDUrd/DXnDH9JcO6kZf6BxAW3Bx+BsD1RRA4LdB18gvK6
0O3B20TE6QnWfCm43X87znFEJJrenvVYjVw55z0Gp87qjgssjBTSKh6LIPkfER1s5mL/EBfyeZ0M
sFMVSWAYoTZxnnXy4fFS/l+gTBKz1+urrHSfgh/2REtjZfWQJtLgxMrZJk3HwnrHWU6hr7QAG4j1
b/7UowdwtzB6KecHkqvVWOuYCyXZNQ7Qjr/oAZZ/q1Bk0cB1QANn7G+p5PVb2qpA4NCcBTr5HjAq
ZGlfQ4G1F04JPeFTr6MSHF9kizEwS1Xpn25wLPB8gpfkMQWInfOcZsP5ViTeGgPjLcQ8R1XmfE0H
lENsbaR/5Fk5ggLtfOfI0ttpEtzLgBc8jaMxDhb/bQHBWRfLBw6A6+Zgkvxl2yyNYH3eHvmVj35b
v95zbab6t34EWoh55GJU58eETOZ1xkLoZ0Bmvao4suDRE0WVku5K7TeEvPqXciVU7WYLrvzhOn0l
WkM5UXn/XeThKKNOpUCPRgFzdDW26ZVYik6kaZD3qyvE/cSHQgj1mN/dlK/WtK8irK6uwmyOavrt
NNnBLe25iJ7uvQyvHJS8dA/m612+L2SPcYPR0JX7yzxIhWisBmctLN10lGqF3tLmFyGywEgd1udJ
1iOgBnHwDkuAypo2PBsx3o+67SO9XdaPYxO/SBVYfTYjxvRTMjC0xmQT819jrNHehgzML4p6jftL
ZSdvvwXKRek3AvczBo6xJZty8r8ZT7S7PuZdO/EFBM46IQ3dRdn9CWRvB4KxJyXsI+e1WENi+l7/
XrsRjGtwkPIYrwGQC9eNfUG3nlChCoVV3vUKbicWi+9wSThztP/A2gm/MpZCHXbyeuNbxyp0qcdX
RO7d0qEl8AHUmUP+Ei4QKpwPcHMHsvIO4DSCfkH9ap8NhLjJUdNchcmNgwnqk4a0fsBbGub7FTsg
/lbxFJsFl3F3Tnugx9DCmoV8rb7VazeyU1gVybAwO0RHeBl7KMZQO8dASNQZZkj13QSIsWyk/n1C
9zxewWo+bbd2rHMLn5Gw+CExn7QJk3ylKcSE7X2CESSVkB7/b+NjDtOFUHLOSR3GQ0TOXLWeBDgo
oaI699vSRnyC+zbda+dadeoS6aoeFfVy7ty1/iZAmByUBpF7UhWgBkvM7khjDswQUcApbNcgzAvW
42/WBxjaoz+5Y180D25FfHsjt9wGBRD6dVvG78ghgKxBQpWekyJSTpAgfDkKeqXMrEsSdiSzbeaO
tHtSPkLkJPZJwQ41EktDEEABNPtNOPMVg6B0RVGrfwcMzOGXMasFaGQr4M/JZjW2z2QVU0/o0/aX
mdHM8PL+O04f8NTArZ316ruTy7gsvoihhSHNVO96C27C2NR+rw4CzBU46F+CQyyhwaCB7btAIqPF
rItsMqiP8KXkNVv2OPGysycOe8N63soglv0OIDMpzvzja9KLzJXERHhrqkeYC3l9o4n7T1HjLkaU
sSYwTYBTf/yxzEAsGwYjebCn7SNKNuINtupoAJbptU8y6Pkz2bc5jQOCFHK/7pok3rqgh4pY8QGP
PD/uodjnSyGUgefW5G4b70g9KlUIlxgFDX3ENmj6ew7dnP99A3cMhc61ir1jE7eTmU1elVAoe2P9
ODDBtqEGNJMySHBBCOKbHYQi8ry6lDnWDn3MwlEKj5QmHNN69OUrHT3RkK/8DYZtFwHR1H49BqWB
hE8T+Lu+3UW4E5OMcP0l0PjixrhkzRsUwLiBju89qwAli8lAgnMqEwwx0OcfydwCAJZfw7DswShi
tHGkeY8nKRDhqLIjb9CcuywlLfY+RckYxarO3pwaBbfwYJO2EKyhn+X5u9q8uf4LOfIeBvNWszyB
HP8voLCaBiToZcX0tiNU5NYnT+xaAvyElj02SMpPLbWab3Cf1f3uQjkhMhNBadkA0sLRAT5b/YGF
wxstXZenqPWsDPzaBaXTzG9Dhg2BF/bXw+NpEtL1vqcczKuRxZdnL+6mVLiFF+Si4mLVjtp6+8PV
rnMLAVVMu3J5A/LqDushG+q6Lj/gu8QpT/+rmkXJEimMf3FGV49+szQHAQ5pT1ncxQgmwcZS7hhv
qk9FXY9nYjoLdeK0dUrfI99pFJ7fLDdskp0A2TKB/YZuyfAZkzrqhDWbeMiOd2Kjew4RbMv+iJCh
WmCg1zUBnGjqsBOqpkuzKX5B8QqHR0Wug9WebySmt+MzSAUiiQGGSQnoo73bCeeZrI7/mJY3zSXp
aCsM4fYuTLy2L9GyCZHMXa0/Sq5/ZdxeeO9HF3zqtF/bwjcFvT7gP9CchVHut+eTKnZ8ZfXSOjgb
HPjUahKKOed02dXG+BRF8fVR0kx/sPM9S7Ku7DDBb3Y8xGMKR/zC3BL2t1s5gWIuIYEIBKhwp0DH
RQLyKk9GLzEZqV8ZhXpDrLGj0hL4tSUV6zxLHq+KsGbpXxtyfz1gO+anVKmPsv7VHa0SeldMkYdz
0NsJvcqZ1lOgC2R3dsdvUT+SB32xRUPTgisfh9kty8fxRMVF8hm92Uf7oD9u+H5Yak08PMIrksaj
MDXOWAjr6NtLS5MtJ5GA3/2PzRRQhC8QDo24AI1ntT0kgYp1hB3NrJlAEJfAOyO3Sqr923CapI4q
czxjSNDY2kPFGgwCGA9IKPzc9NpwqVv76YBKEVCS2ilUW/qgExxHgY40i1s1OhIZT7jVgm7JqbC7
zJ8RpJEpxszsBxm12i+QvgeBm5lPXjBD4Dtm3uitQcK6JBTKfeVrEhmhdyEYpMBca8JLFtkmgLPQ
vOHD1CpgN9/jCyH82DgqeH9mPPccsXc7FYxxqINHc5LifDFedI5E42eyLWb3EHlwf3XvmpxcHLMk
mnIQC9mBj2oPtC396DNEpKD53xBQ5MhjGA1jS36QgpsRihsRbYCRyhVN0XiGsMMRD+g9PE8wyHd1
I2EOlwDLDT/GGvYE7pnTCvGt5syGM5gEa+hLfGn6lhbip79p7RRAXPKGirktiT/C4y5OujfX0EmS
GLMBfEoAj35Blj6F2tQo7LDwlBMdqQeV0Atx2AVNTKaPWUiuzGu6WF8I/Lj/lr7NbcEJUP6c8fy+
cD+EHVc57aqq7neSEmKBI4Sbs1cYji/jres1Hp9jslFyG9DbVJq6px2p2gt1jVAx18eEzT5y2DJ+
SMt4OzlZ0b2ffBXX2UGbC98mIOukQwdMIr599OsInd3gWzC6Jejql7h/gc25Yp7SLPSztWMVL6m9
iLPCydZ2KR8ss3XKsj9UxrjEZy93BFo72hur1vr6L0le5AJSOdD3SS287oNkHBe0couvgjmq8gxd
WpFg4AFd3SdiA+20Q88YKZSak95ZKWQNozg8AcTsxb573p6C8OamdBHSWmtLquypby1Wxj01e1xG
VeweU0k7z1GmHVp+Du8I1CQzrqsJXLa8oDx9b7wquJ1JH2ipFV4T6/fJsiJZY1O9RXjQAyKKtiop
a46xEmqK1daXGLGabcw2ifeAYlgbyn48KMns5pBnXnoY0CTcLmaalwYKAF3/7rqcj0Vd8PWry6Uc
o3vDBBeiHBLz4R63x+8UbOAQalZM6qr9aj7+fBkvc6GJlyqZYQxbIWDs9O7mPKbk0z5TxiY+ehNn
SM5L336FD6vIh66+8HROux87wAyVyeHYOGM42pjMn5dzrY/dvsqIFlHweAMPKKmVhmPHAUI3bx1C
+l5n4PAIahi/xNFN/90Y9Y7gQjn7x/+a+HZNZz2SKSTO7JMQK9fKZF+2lCQYz7xHHmtZiUKem3xo
3V1JcxxNILnP2HqD1PrLFemin8BMJIwxT54P+qBPn6+lLeSsAR78mkwb6AG4SwbgSWQzXKenKkxd
A1L6HINmKHYxZxlP0dzIZwQ418gerHjDrcBQLJt3citOFuVkowWuj5t8Ik6gVxO6mB+hDIqjNeNO
XWv/wMYNIN2EGORAJk5gtyGtDwC01wHyaG2RgSETakv3ZujzRAEV031zxjphJvASAq2Z7jNX9fy8
ohS1zK+YHQBTVj/o67m4Az13Kv2AwVxAPQEIgFcVDLNZXk+3JpG8TocRcJPoD/SDVgsYxK9IYIam
6mg0myXekTA3ubyBqcU8NA6v4wXU4aG0r7JjbCKYRbVerM/233W9cV5IXb05cIOjqh4Jr2vmghbg
8aMmcF9NNds6luF9oiwTPW36fF1vAnolOrN/fipib9UBwdxQs2Z4egP2uqc1L3HgYZ/Z0C2Gusjk
x0PXZzto+eQO3V3cC+FBwE0qV4CehT1VayimleldIvN/YvUue3ME8TOXYC37nHakYSEXUAIr6NY/
c1DudzvDoAoXYHIplvCnE85BflUUiXxQRzKS3PdUKPy8bQeBJnIIAtixb8C5GPeMmBCKxAJ9ngIh
ezLFeRPNd4K6OKSBLK5cATCctQIS+xFfhuqOFf3ij6VGvtaHDnT7fWDKOj+aG+dZq0jlf+ywCk9j
hbxr7isGqyVgt/jXGzaD4pNHIvSeDRyAJni+8YlW1tuy+N7EX8WbPe6bY4otZmTotQ/TxfA6vwiO
wHfDC1j8CcEc0eAUo4QYuAXQY9IVBHZhjz4xRuYf7+pk6tpsKApLIBr+tAia8tA/z3nlDjcpeRoA
Ky7hvvjhrPH03OI3IUPljYmoB1neXcobBjF/8/Udf5bwddRQP7Kpmz4fT4VNBIscyXs3J8IXp14h
P3W3kkZBVlyn8/tLcyiRlc+DgQ1w9c2apAsS8b8qyBb4AMrVhJdlNyKLYul0hwW0i9tcfU+v3Ij1
0iCrSGcfNRbhS+7bNUmAMOsSHRmBe7PGefkY44ahgC4GT648k/GNGCRZTPVyQyeGP8UTCkoyv/gc
AyRquCKdbSnpAxeHGzwKWHOUM2COYKap+8Tqq4t7YH/Y385yOAJ5ihhzSTlRDkotyDwOcK3bQ1VJ
O7DsIHIYBl91JVNaA0rS5tRjSungssDh/hxfrAPwhhyRUAmmQ959prPv97jDXdGEealHrtovLSMM
oeUvYyYf5iNhpBW6jOWZxNSqDtx2YP1CHqP5rA4mJOmN5hth2jvSROOUu3dHT+3Ij+9Opjyivtwo
8BVtI2Mtvaql+3JXd1sWuA3jHA2kAM0eNajgmTv5KSharpqGhpMf9S294HP4Jga/EO0Cv/aaO+tu
Fpf2KPx6hOU9qPohCeePhIA3IIkfiWpS96jPtWGDmUfifbK0hWZYCqWChD+CroKa+jJ/5CoYgAdt
fK4fXTSHBhj4gr/d5ChhIg3vKbf3g6nZHt2igiowvN7sJIGObwbcgn48jWyOMklsW71l4v/vvrRX
xJgK6ussM+9GRL3X6d+p3J2DlAEc9HZ4qRuXeLtBPMecspcrb59gVIfLdhJz15T1JQR09/7ZvsaJ
212z/dCc1a6CP4k8dsZmkP+AQQaJfY4hoi7oJTTwwY6R9EgxhFSLE5kUntZij17tqX/pCBuTmwCd
5KAeAN+y6wIVz5G91KwQpwFj9YyUDvnmopzC5VXMNO8VnDZodf7sDGfYx9DEcLf2v719ToEB3/xD
81yOhDnfsSXhrkY15e0HEbJECuZJHbn3PWwNOvnoUQH394cLRnaoGFz8oGjpm4XpBn3uBS+bzJOn
p9s/SIiK9elVjx2mjssbAGgsIuHihJ8dWE53C/esCw8RTUWs/G/dySVNvZM0DCCQuxOTvpTE2bqx
EfM/ZGRGEVZ4+lJ+ypLnFRf0qq6Ny0QyTxtGhhHujTuMLszQsElmg3DwzIjRbuijr9cv8VKoaVqS
Q9+s08fUsFpXG7GAe5524Q4u4a3ep2QcO0t+Aovc2vNk7RSNhOm4WuA1TInxzng76Prd4MRdLjV8
9eUFZBTczQuGB7rVkRaHMQY23tYbx5MQ27trw2C74zVqQmRK+Re7KggW493iPJPcbAQpwYbzJr1m
mezB+IhV31zAwx8q2skH+Buhqt32ptghEQGQS9AgzbaFRQojGvCat1AAT6Ix4qR+NVzTzgPjdFb5
PpHzuDmB5xq61L9N4IaOO8Wdt09Im0KUWed+ORBD+UHNwm3LySRL/34m8vGzYqcJM2zOnaRki+8F
gnpkVE1+BjTv3YXUbaqaRhKqtX9HuTkOCjztB+R54JgCEgAPGs6UDRiq4SkfAzgWwGrM4KSXguBp
gJfr22Pklss0Blzh+iAAgNdfXzdXlENdop1zmMAQGJ8RbE2LSVcKQH0qPNn1ZJBY+foZPoVM+Jer
rWCImYl1dcHKRDsTPSUGXZ9VRIPpsj6Blkmf+LO6UMLBbdH6bK3xoAsK9WNtCo/aDkhhdFqWZrgI
0Ho89aLwRjuWMSioVVniQeGyiaIIuNex2U+bqn8jPOo9mR5hZuwMpoi5KaiQTtPCL+KnB6C318To
jtaUMzK82VqDOkNDR/YPVNyE1Ub6dClXrQIO9L8YPNZYBZt8rvHbD8yO7D1ZLzQnWE3J0OPjMcvM
XZ7al9YC4hHxaHV3xA9yAUjKBSgjZFizE9Wd99fJ0bx6KjIM5xsjiJvCXF7cL+Kzn8YE3j3Y3Tnz
3nAm+mVrbCMBYJeD45jQWmlshzmJ2UvyyiP/74juY/dHcwvMhv/UUyP8yveTfIqlX2wXDjolYh7V
pm8EpzCM7RCZjK9DYDR/CobG6UiJQAepAYqQ0Ns9UPDwf7iYfeRBb59HYsp2qXG05EtXMBRa8yT/
UfwHqfLQgC0ZVcnTWsj4DhDPXcm7mLLS9v/ZN5WVWaWx1AFvDjenyp3Sdws5b6yfPE+BTN4vO39M
VMd5hYbqV/5f7+xkI+cTP1jf4Fu51oYfyGERbJWOHmNx3IcsFWubGuBP+TOHwV89y+Ij3qM9RlKL
Wkgpof8Z1BVIFRkzOCpEtxHFsVW6ZJurwILNvmD/YE/AYWlch0u5kmq8ZP3f+0yTIab4u9egcTvx
PL69KEhEsAe67MZtt+dueZ1a3LZFsNv/idXh6J0ogIHiur/9RiV+hAYWuWx5QFO97GW6X3j/dNMo
sjUZx8hC0yw/WsILmE9Hqw+5t8BwTJMZ63gWdBVafrm3orBXJlTGyJQM4dkPUbqNPUxvv2vdX7Bw
jATZgyO/XE2akWG3d6LADbTrng0b9HP6OZUZFLTDlcM/nuteZjoQkVNVGb17JbanKd5pfRpeLnnc
q7tS05CbRrq8Q+IuhLdKVkxDYurMJkFvoa+ujg8iEcZsWj760BPzoEdfh283wclVPOwFdsh4NRfs
lly1gal9Z5l5GtfWFt9I+zTt9SjxoUHHAdM/vXEIoyeCnDQ81PZojDjtOskXXZn5oGh1Xkqqg/Ym
eiGE6bDtF1LYrj4hh8RMD4tyLCoTrN3YrR0kM44uJzmsN8XhGiflYdz8YLwIc9VW93+y78xuXbqN
UUXcJxIM1GHPZSSrnehr6YoJ5QlDjR7T16t9pr4B4IgbjveWKYp222+Hfd22wiB4WoAgTlDxTYFg
sGpQBgiO3QPj4vUyKphoQA7eutodx9qBpZbfSB3NrpF8xruGLlL3Vi5As+I6B001OpDy7eI5PcOT
saUxYOgDAj1k1DANlPCl+qYYSMrtXWd6oMEgaYgfi04srKn8j1YcSC60cpIPUz6zVB8d33TCQh7L
DRoDToq0kBwumeh2bSwqxm1hkWb9NdG5UQ8lXsc96IfZpQ5l0DpRo8kK8E3aX9ub3oAWFiJOmSs5
dqfw4YmS6OpZ9lgay6L1p/f7TyiFVVEPzp/VaQuSPDrAI5yghoc/254qj6a+YDEpPbW9SwS8uT0F
ARj2mJutkpqAvGSBIM5ysWgd1e9HWSJSXLULyU7TKwJbVtd5I+0pmCbdFqyoaE+8XNhEPBGA0GDl
BWHwW8mY8AAivL51W3lx2lxdvI1NBAusSEKLDm4iVbJdC31IA+3lrwA4qD6io6zY0wwnAlLWKxb6
FlVQE78ydN4gdgffDN9DM9K9/+axeCOAszM3izFwZduEH1JF6WccVAYzNqNy54rAdW1PFkfX0cv4
ipJZD/nQBS/aWJwyfx2TGPwpmbeD7UR6nafh/Mrj7a9TEt2/+mNJ/AqftVKyYYjdUQCBDD0hEP74
QNBo0YMy9rmzeoRwrIhqwpaXy8gLr33JhIxV5o5Uxa7IDh9biTniRqemscwpwLBG7i2YmQoofjc9
PDyvxYPNF2l/7lL/AYuVz/a0zbYDjdXCHse0EFvavaPqTEzT0DmJt/yvy1ldBu/74lJn+oTmoY3o
9+kSjWXNA5CH5/i1mQ/1OrMbx6jk7Wvz5DrXw8dBTrM89lYlLsOTgMq4kxIepggZpr7J8pL1QIPJ
ist6n29UNEy4raaSDmRGRlxbuiLmNIrklyAKmNFSL+m3F74tqTy3kOfOF6c7B+k2CM6mCfoBuJXH
1TAHi5/QeSWleR8t9d8F77L6PvV8y6KJi5miz02Y5KoG6fsbg3eKxlQOIqQyA7L2sOHJfNQypgNa
dBNz1PQNP2Vc2xonEu/yE30mxVrwuxHwjqCmPSLwHAGnyFcwAO1G/r4+OL6jwveP03i2SqxLKyn1
mbAPZ/1uY/65aEH/68gj4phDZ4f/OWF2wnSAgszmsNxHfEYHTj+ab8wlTYzwQoqlCIRsPILdepZw
Q+rO4wPSqvCiQXD62qr74ZJviKTnRjazEjo9zWwzX4pG6zyWNY0ahn5gFC0Y6Q3HsAjuYsaGVNz+
CZ7vY6K3gkDScassKawod69mn9pPB+evdgvKbGfBGHAdNmmew3CisMwcUm0EK/KKYAadOJg2vTBg
rXhm6bAncAVdJ060bbv57N3pbXWX5sBfc0bLMyO9smFYz4KpKlAf1jc+kk4/S2C2r5UHFXV+eoPR
0nPYcfAXKjjUSfZNe9PPWEXxxM8C79cFSlQom4fRKI2hg7R6c2196wBHNi6iwuBBiUH4z7jMgTtv
zN1iDzpqswMweNLjqbRw4rh0eLolQr7+g1IKHx5UyuvxOcnIyeJaA7ic/t1CYmXguZybm5KuyZV2
J3bpEdAS0YdavzcjGl3KAbzBY5m/7MYQhz3CANCt8qQUxKr303YHVfbEsLHqHL0RCHIWnK0eOLla
Bt/gbvlA9p8zndJotrrXhAwa+tHMDFPm/VkWmzVAdUhhQ6sT9a+4Plvk8NmuATWeocoBW5QCVXVa
2esAM8YZiCJ9HdOngtN/mhXsclOzFYveWiYSYeWT4pj7uCErlCrOUURf/EWb0QvsnDT5jhLuwG7q
vIcnvfmSBIA7wcuIXNFymb4L4ZgFuM500HaGNpjohD2I5Gjemc0xDnfUz7esN/a2ORfHB8L2/K90
NMW1ONzScvaGlPQzv3cOISUbqf//SY2HqholkJAJvcm7Ri4EcXG6leMEvk7/vBxxbK3469B/i9o7
3DSNPcUv4WGLpim0IuNvjVsPmc0azg0gDtrPGKpU1WzPB/CWzfcpuO2kKCVZZJQlgerfzdk6kXLV
wcJ8hLB1MGAKFbJDUbZa8EQmGX2dz0FjcSX9kdHDRr4h4xduMUBYtl1gIMpT6ucyaZD4YWmLUe/2
ugiyiAAegZPL1ofx+Ycsw+NmceD72jjNaoblNWTrYLlyQwgA7XpdJR9VhAuduf2aJ20g+ujCW3BG
L9149ABA4l856rZMPsKkKgp4TqZkg/ru9NiN+wIMYGleRdKm8j6o3l9Ns6oKp7mMzi2ntZ2+R3en
A5sIF04R1BoAcd7bM3S4ZBceuNd0W16oYmeT6gA+QR+8bq6vPJC46HK8bVo6UG+19Lb4XZOwZamh
mlR78UpbflxdbbNogA//2PHF7tzhDLwl669/zoPbxe0VwSsL7PVddHWRGNffrwSEsrzKu6BB7FNZ
bjJ+LOzYg6jjHLQPAVS+a8MtEpnS6ItLt3pI01CPMbex/YeKcwJE0i958AbWVJAPL5WGe/WqZcQE
Bi/AnGvEVHKJYB5vBChRG3hiAboJSPhgPNcfwFQ3STO7g902zus9yB/dtNVpD+TDfnIaZoisBd4w
TepwSmdUpP8+7a3XFFZyoSgrp9M3q7lTWBv7Ra3+1OnYjLgRz662tDR0p3MKfB/UvdAnTHylBqLn
o7rgfepiHkPNT1U9QkpFl1Th7TS5jyWkOQCKr/YlrVWvIOORUrPVt3GzyKGbupFM4TqqTP0yBAyW
gytCZTZ9b3UaUlNFjCTqTHfsvfYjwSDbD/Esw06VvfNNjQ+6oeMF7mAVwoNCkV8FeMhyrDyKYyjO
N64EOOfZfro3i9U3xsT5yqU8DRs+zgySzpCLB49YtImG5L63I7hQfJjroejq7E4x38Izbq4IhtCn
jsOKv4m81vRksoLrABVJ8k08daV3s8CKPmacmYY+zqy2ts5/W4AibzceEIS/TrJE4aNE/RoY8DqX
7znublxCuEFBoB3FxrP/7CYnvAxvsUUdPPa2+p5vhnzZvKlCWW9G8apyEhNDim323njTOrRKamMr
sGWDg77fVpGSfrIZwxKsAb0yqy8+slqAL6n01r2YJS+yOSB6oEygaY2//uH021wYlBMcyeEVmNZ6
ZuJbQsK72xCNWId9/q68qLZnF1/MsQQFnngxF0R3w7YyVgPXtmHD78abUq/20sQIE05KY0xov7V8
mpIq+lTVJNRcY0jmcEscZQy8VLGSe2P4koF2xnyvF4Yb6W7kAKD98CUgkC5V3TtuMURAHxqydHkV
LwHTdOZepR3j7VGQnSHa+lrfMFjPxyYh5YHYXMf/a5kIQ2mswSLarRy6P4McIBw9qRCxjoVTPhx0
jNhO6i1zAjwfEDdxFGQ3G4JETglwjdOjkA7v82YikQ8PGE6Mg2V4Gh/agB2bj2i7YX8y4bdVMeTq
GSdqR7e/fD7oDMaiczBL5YupqaRDZRaZahVDSn5/5URyLuBLlWdOLY3JUMSZiG4kirYkfpq/EzAP
HczubUdSUB7X/WLjsngdSOY6ybPSUIhG3ErYMzQdWF2XQiezlfktWjAqdXBV78eP1YJ04aix02W+
WbjAjvoOtVHKz88O6YG+665L1Gopzn0acwuLTP8MCsldTqwcaJIaLu9X9V5bwCqE5EsRAXVRnSXQ
gEoTUUl1cdJVbfnAQ6HJpdgU1CxiHo+3xeo3bq4xJFZxFpgY+MeGHaI+BOfJQNhcxPC++1eb1mtm
iIA+y37M3nsyXQirIZixpZr89FiJbkAPZ8zkFt7f1jC40fLvli/EY9UxJ1rUwmoXeJzEzH2Egopo
RZxXsLx+lqgrmfLkdL/0ZXIKBVkz41BueGnroKbWvsKU36WNYtpYXAoGfO5uofvKOYttGk6JVnse
BD7juEy0oHKZbygERLpD96v0kQBPWWLIsOSnjUuII35+ct03ZmeSuQuAMNL6hIXnxGakuTytB3dO
c127Q0krBJzHtyGDw2UXJ9dGOALH0d89gPMNFvCJRaHjoi8rVT+G18f3TUZkE2YxBuTyHcB+nm7L
Z4T4rj0jVzFjZAEKvBvIDdV5eRew4ItFPWf7TV8eZ4qemQmgHWX6NkNQisfe5CNzR83vmG4mUM7U
YeyBIjEBFbHusIHT5Ord6SGLOoQt+WJpvDppVl8Xv/qeiEPCIGGIxQt5bOojqR7ReT3Ua7KGCdo2
ZY1S1EhRtYKYtfFpY7AidjrB3Gj3Mkow2FxAe6U8b7w5qssI67XPnY6Q3y+apT/B9ldXvDUjr+gZ
29qmhuJ9kEF9wGD2+ebto5jVy3Y6AisLmilhHNsxsyngAOfGlTaffd+V7VEo4Oann42arDSES/v2
yZaARMIa/GO1kQG5v8nhORlqa8BEJtsNQ6SWSX49FQfRxjo5+cbSmPKp4rHRAelJrdflvkTfvKdH
1qzXGM+BtIYwLo5KCEzgoPrl3J4SxLyqV0CdahETqOboFY/Tetj7lzn3p5Nj9tX3nCB5dZA6n1vx
P+dvpGexbtH48sRFdjERPmBulvPWExP7w+js4chyIFPtNQex5CvPOgimzdidM5JFP13oV15BCfh+
uO50xy5OeGHokn+38ZhxAO6+vg/9to+201FKJ8ZqAe4t596Ld6F2ZW3GxVUdmlX1bcykWPld3hFt
nXpctJsR7MPEZAkrwhNGOcQ6+4txwR+wHQ5nvmiQL+BuLJz3DH5SZ2NxQakvrs7BUSMZeCMHJoAZ
eDMrw4rsTYBE4HeUdTu9btrAiippzfTXJv3uYJKfI37rTkOpz8L0HfgviNai1re8UtuwXsLrGZr5
DxeH+FQIYCElc8h58FRnz2i1kv+obJ3B/qWmLxgMeQGJmPlvnvDFvZzhDDshBDggE6hwTbDSlUzR
La6daZrlJG46zYt0XvWVENnvvxy8Uo43pyPpGheXuMZN59JFb6Pkl4LALAgUdJdI/Ah9KjXwBSje
Kz+zhRIjGZLIgOh26yywsaK5SFheqBxiLKYjeVc94zqU5LFnOgr22Pg9K+iGA77ACHv37unFDwmW
KQ/XvlOdMJTvE150sYid58HaaTq1UPeNC/LWX76syj8tqqi6LiUZ4RGsq9JbeBWHSnJ8fGWmwCLA
ciQD8bHtsxDWaJXnAdDw2+d2ZT+vKLRhC8LpoxIgnLlbPaLq3tFh2SxtWMxc25CQsHTd0sJia0wm
Hlf720ucc/mMvT+Zy5OG0x9hu1rN5lGLuT3IrX4WttBvelbaIAmtHlWm9e6dAA5BdXrqnYrJgReG
bO8y3pkZkI4yx86ia7j0RWi6GUMuRCt5/DTR+7CNNHcUqTCsLhrJzS38HzLsV/OpCmoGw/JScMpg
qWllRW7Sa2hsHI2jSIKW24j93O/ujQZRwxWLASaHuCz0x/pP/ianf67lP9OubINIBKX7bLFiTeZy
Wmy+3Dy052Oan/2XjT2KtngiUO2r39EtlOF0OXDM6/ZZHcCQNijfedS9sZoRAivtnMWKI+IkuN1C
CwcbdQaT1LRm7UiPXby9jBkVGSWc7wiQSYVEwPCrqIYdiUADF+2K2qyI8LRWL+mJDVnVmgptYz/H
gSPETP1IF56B67YYZYCXTReXdweK/gt8hvxu5Pk7QNSAAjMH8C86Mr7mBB/rAMsDZSxmHLZCXRrI
CfBVN19qTdNR5gs/1syjaRIuXaaHbJuH2w1JWYEF4jJJ2PleoLSqlbtnW+bPIq0Utp96EFcI6Gt5
UExxwd51lvunT169GEfZdHdxFF9Aanmd16bD7QlhVuVAvr0GoX5KoyiGMOw4qIcm28PpywfDdf1+
GTAUqjCpbACACGVKswZEJJk+Hi77BM2kjezkza9osOTC//zXMeGreAN80ho3qjXrT36PxbUh048D
B2fTLPMNqvbSVRNxscKGNjaEsBXYGvczh3Go9z0pHYiLqQkESr0M1zKrDEsyQSMh3GPnUKL+HSo0
cCg7FPKwiA9K9lPaEm1CSgV31lS7RHNCQfOM4NljKzVaMdnVJTvQTdZ7WpxydMnMZJmWcMnJo64a
+o9wzqgcVuKj6PDHmVX548nWkl6Rans5n7g9ccjtaU/a3dxjrmcrxfLuzG4G9KvSLuUlJ4+rcwJM
kL5MMtHVtIo1Jeva6yl2kAgaOisTJbJPxcmVeoJtONytSxbbuPuYZ3F7Z5fMkZ9o9wJnUdgJHd/h
QprgDwwF0e8UQ9ijZ5sePNJF3H1txMKnp8Z291WHtH5D56/1i80ZSqLMT6AUbGqmxSDlvKxmmELg
Cy9PTbC6gVDDrB7p46panSpsivRTAzVVErjgyASXAFf1oAj6C/K8xH7j/JrX9o5xprYL3VuosEj6
sTZUba24uO4lc5GEP3BpZoVwAeusxBCj+eHVzXtm6Le2ssFOlEx5+oQ89hU3vqV8rDhDXuOUnkjY
P09dNlWR0hA/MOrqJy1ZFgTR5YWS2lv1x0TCB22zhY03FoegKER5LiN0nliabiLiRN6uIb0/wmNl
hyRDpUMZM8/sjMl7hsEBGLO4ZhZvxdpl7DV0BW76Ogfp3vWwakQ1kXazmtbQ/Fmx6bWPdEnj/32Z
yciVdW+OUUjgXhrvppmWnNCDI83SmksbVGuBH1j6Ar/qs1Oo7QE2ty6INqgWNtC9dcHBpcSoDjJ4
KLFfTj59lJsWOlRJsKQZBBO1qIjeDPe3/03zROV+x1w9OHfHGVksggZJV3gKep7I4gPQedFzR7Uo
aVUkLEYn1El3LHTY7oETLmNNmgmzqu92frvEjlus541ksQBOZSFgs1Z1GW0k872jhVSG7jDORH4+
E3Ms+KRTaWrc8iAj8/m4vYmFAQLNJmHnRLe6nmM9GhjLTjrahVb83GUUEcPUepzX5CyZ07bgckmI
pSZ52uh45AnlTPeG2dMdJDz/13UYhcVXGNGi8jQFcsNZDW60MsjxTrY1wdKwH3xlaB+eln075/MZ
dkf6JaUe3XP9aFJN+Y/KqUal0QuAU32NMFydVGhmho3uBxrPq3WYyNDP/7JVEpSLvchWQO42CvNJ
+kZO3Za6Fk6MhyRONHtvJmBvv38Lns/z6muHKEnnLLqfsT3NOFemLwz33cfSYlOovKfmq9XN3mKp
IAG3/pbtxfLBgSpgOc1RKNcCYsI1DjWc4EdgiBtFDHkQ3+odFFtYlQVMDRIMGaX7Jh1/JtA6ENhc
GJp5KdVnyuD2dTwTGiBtuQazdxDFYFM2DBU10b+yMp+2FNfxY+p/408DlwG5umOiu9xVRHdR0vWD
JZM8/ctNve6DzOJ8Qx2tjawKKp/U6ASAvV390iiAb/ADML3l5Ubqljn5vihRau+SGrUkf/5YOiC9
GBjjNzgsrUNvONwYGXn4ssx1t/oYrflYwKNYHHJDGFZle3Q8NJT2wyMWbOWamYlpAvArqxeSO/rN
h2gITqDFmI+4+z8hf6DSaIl8KswL58j/H1hNs5iB0XKONo5gv8FFDD8WzVOuiPExHApwsFXGUB6b
GkXMIIQMUUqCUTgYxymSzs0Pj0Jem4WccKLUBOu2SmiTVBRZFEmXFA8DwqamzbBzsFCwKVh1IURI
J3iWM/TM4TGY+1eibTzBDt6ebX9812/0kmpvcCZTYFTimHNSGlmy8IGxes8GtLfJ1A5SjfUuc3SX
B8Ta3ngJfOn2oncFJ80oYy4DljKpPcsoYzF+sdaNbWBZgr5qEqh+k+TFhdxAPXNmIVLqwS33lC+X
H1XpSJtArQnhjHRU+BaJ3CpR4fA3cDpjP/1n8JkLM1iYqRzlWWNgOXDRkjo42jNFZt8Rn7YA1Tfb
j3824Wfndz9lLWzPjrgHpNF1vRhivGaizYv0z9kR66R3XZBt2azaCq5nwHEC3kZQzQK688OPwTAs
HGStLscBrFIiKwAtn799lyryIUjFe7zOulKgqM3Lvj+RR05vBBbX9q7xXKOsd0oXe5KW5Wl6ndUB
UMWuxeSbRJxBcieiZO8/KLsXyANBwRcXtUHvvPf75RW9kabhl84gyq+i054XwbAKFvuoYGoq+Li/
V4y0iMFiOKTdsmI0mWPeTR9W8rEnYy0QSJeVfN0O7M/BSCDwcSeOTKoq0ox94LiMeYpic/XlrEzB
J5FawHQ4izh3E9/R6tht+UHUGv7b2JhYR0dtYRAgfW3V/Eizn5NmXRn0SLXBLA1PLfAtci2YA/qk
MPz1SV8qb3Z3zGQUG629U7E2aJbXH+mZTBHS9vdTdkiOySm+uZp78q4Ap7HSCDBj+qMHXPT1Eevt
Pb3fmMoWQjN7DhtGaDZkF2jaEHMe7zJSWYqP8Jx0MIPQFW3OHW8ytL6EOW51G/rTAzFk1Rn5IakZ
2KhY0uWAT0F33wJq3aqkij1mdOMNAp6eaCYhrdAW9EQgMM++RnRmVUNelcfkiAzHs6g4V+14Ano2
fJODJX5gd6yS/sVjV3wJUx+5bjFPhkD+U92ywZeXvqxmCpUD7nB7EHXlSJY6BHI7lHGOqxwC4er9
Sn2fEavgtQF4VSBoKzrQRaiQeTUYhAbSTVBv3Yqqih5/8FP1YTNdlP1pdFh47ItQyrTC8wfuNstZ
IhuYJb1Md6WQ9GxHOpAqh3hzS6mFbaTg8/G7XAhUiAiPds1Fxe6mgaarTggVxhHbhSH1Jc2EgoQR
ZQ3jGiZ12LVBvZWWktUKdp2Hq5qg9phjqkL9w6jnN+UFh0cgEsn2fLmeYNfQRd6KLSFn1JkFJjg5
6B4rK91AhSrSGl4CQh/YIO0SNPDr3qqcpfxGD80uvQb6okDZTm9S9cepA1U2wp2Zb2SKiBxK63oJ
k0wEWkIVcJgdIlY2jHHWitcy5JSbhE1a1Sdaykk0hF1c9RLXWbq0N7BtkLPdb592miAhry32xTX1
0Bb/NtIEmqPpSPBdkvJWQsK5gsaMlo5p9hOwc7ZWL9lghOKj7KOreSsDuF2NfR2fA4hkb9eef5RF
AAb7NCQ5I1Ci/jVos7t4pmRnrBbLDfmrr77ikd7ZhipnuDDPceG5Uu73yBjeHoCoL3kYgHHqBi1O
cSG/h8BI+tSfS7pMno3M1g80dykyC1Oz4QGtwbHt9KAAGz/mf1mgw3pcv1vdSwY7aRLdwpi908CP
/aKmjOImVfikWaHg8aVYuOPb+zVPNi2ZITc7OWcEFyFGBeAI4W/3il5LIrXnY4O1wc7o3hqKMLyS
Q5ROUSt06T8SyDJIjs0aS//H/RJT7MyEl82iXackldFq1067osgp7X9lgaKog9w58ZpsoxKZ8dae
za/syyuSWmVefWngteMX371kn4rBtV/F1/vQ1vy/MnQ/qFEH5jEXadYPG9OeIfKXX5goYeodAHwQ
jMU9ImXdvuJjgPFLoCCPYkwiNzUDL36HHIa+rF3N433/OFa1X8X3xMV2BcsaiOGm1YTvofHyFAxn
wNPSPJPQNwkADLqTGklr/2wHhZNcIr8B0nrcsZXRLXWeKL8TWsQLrfSc2G3AIV96ERjcGMRnMx9s
MJuiA6IS3TnJxR8qULDRcZ1iN8j3hPyxDJN5vA20ERmbsbmJhn0S/S9StvZja0DxA2RAg8pwbG38
r4KkxY3fuSbi9Ile+WhBQw86YKEC9PuwuJ53NFL0LZA/L5CUkYoh2zulfbpEJewC7/nMvgWAQryZ
mXTHHMwvwZMc/NGEEHqp7UfPeZSPSx2hR287ZDOl2Drxb0UPDtWxc3gthOseLfcyd/U4va2WYcAh
/suYgH+dyAOpqyoTNdyWm5oVNbH1F0E8vtNtWP34plQ1qf0nG4d9po/Oz4SYaU0myTWQ+bUmaPI9
xEyt48BXZFpzdJJphrSPYstgEcSq9x4JkfcD+GfxZToug1KqDUkrBPWIEPyvZElwULWtek4ZUios
p7yGUUShRaK2e8h5XIlHuZ2QJRuV9o7FPvZDlZwMowPrtRXGFxP3zH0pwsMVInPkA51N8qeOf3+n
t+J1MYf5YrMOJ8UZEZHpVMlKIeHYgCHF5CSxWyZMytU1MgPaLahn8RCrRCiMhUHAC0ykMICk0TXh
/TeLfv6QrZhPWtubSIHSs5lMaJqIO1NUeg+aBB+inSjh0bxK3cp1ziAO+7RP0CMtrMD5nJEcZyEp
24Y+15ohMn7Z32z5cBJOp0d3q+qhJMXPd+ipqkvXKW7BfBT8Qwg4bQUeKse/DQSq+4kYOSnInq9h
B5L2kdRCOxED8/AsSgmi6+yuNYSce2LMjbFoT4X7H+h70+9B+lYJoj4IMKLtOnd5NKCPLZtD1eZL
KDQk8x9lBoaGMpy0aOQ5eVxf4ELps4SBdeOPN7P4OdqsfsxvD/dlgdjpGCd8Eik9XWuSwNdWmwU4
EAml4RXfetpbRI7MEvlUPEixFFKZbLlmFBB5HcXATqpg4+zLajd0Fc0abF/ZQLqPXHfJL0D80AK+
2VEqjCqC3uqdq3D5tn11r0I8PyVgCz/GCP0Lia3TRfTT43/qng9kV4oTPA/xTB5y4TJ/kVEgTR+w
sq8CEinZpAUP6KySfPCAf86I+dnetWqkjusgBKR3T4VEV4nTQdHfRL8hZdrBbj1Ljn7rVTr4jYRh
j+Wh6aYmk5bLh089ofJOkbsl8blRTsHVVVo8rQ4peN6PzW3fjAw3WtiSU4poyP9UYDNK+N8s/WAX
Zaq6DKXauh9KoKvw5ZVlq924g4TlGfF0LiUCxG1tfEtj4VrCgQookiDqBbDAYNNf0f8dgHjQayEq
LahTuWpzqM0sMV+H2tPnfuqJlvWjLUr3eurIn1c/k4zJuiKTzY6yh2dTrnOKAQGjYsTq0nS9T9HF
WMueKMQ66qW15j8KcdqcWLOFUQf2hgm7orhXa6xjhIZKZUbsrQN+VdOiELsxWjdem+rJwNlbAHuj
TZa/+qpgCgDmLLXSmVAJRN8MGpk5i5c2VjE/JEhYzE+Zan8+bbFBT9+H/k3A39LiK0cHtozBKUgs
NlDfLXXmw7usV1H++J782FTo55+kCsAEXU9FDNGVPTX87LwpWOsujPvqa6DotpCxjLqRPb03P6mn
RZdPRtL3XGtvW9N0l2vIbNeMYy6IoxW393jMWhnFX+EwOxb1IHHDZeq5hEgInXdQLCrmX/MFP6Z2
5vJEbNvBbSPE3H2N03QvowMiiqLj1pwOGxAcN5lZyHUMyDdjBEJkruGjhzG2fK3aGgLV3DwRqPbW
BQBp2U9AxEP0Obx25atXUJ8w8ZS8LYxU9cn0iy9RWJtTcKi1eZKfZzpP7yWzicfp8xrxqMejuH2L
RCeLyo5WkGS6AIZnc6b21KJsTs8BKyHedwk54rPR4Eg1pwc2lmRvw89fd5atYDXqTALQU/M5AWAX
8gylM9cOfkfUg/VOp/09RDHVt9taW+c8L62LUBTpYBED1PuemmugarRfylx55pcQCGSENNvBerA5
5FLn6ZojoltN4Tqmx7V7YYG/pbdKjDB3JZ0oJYrQOqbTPfwX9RPxS8tf6Gx8Qei1p73L1Du/c1YD
ytFynOv65FfzBR5xuW9Q0+tgGc0dkdhAa/IyPScWRvH4W81QMPoK6Uas8wxbdfRADoVdTnfalXNE
x0K7gCXuOgmUZigYGGT1Q9cx6ta9/r7x80weTkXdpIBBU1bF2CtE+lXE5NiAJh/S5Ufu2S1W/bzA
nirCwNw4+LKYXmTdo034wrXLmBtiIKv8VBAErefNTOG/0tbreA4RUdF4iKKMeBLZ4V6sSQGUKB7Z
GZlrYnbxhtAAEKXPvt1BB51DZyDs5oCbcnLR2e4RKnXmicrqP3bUWRXw+5qtdlMNVy+2cMY8tqi2
xSKXOxaXW5gK8zN6+DOt1+az3EPxj9LeK3AdmCoQPkLqc2UPilYQXi3oSJ0VO2xiOQvjllliLi4P
h2a4eMw7ij4jcXui4MnhN8vb/stBeg+dhlcsz1/Qsar1JbMSC0lHIgDKeKbA2PxXmWapMJ7lRRF5
u+qYHyFiQILRimGr0jN7zK7Up5Qhvn4Knekj2unWB4i/DZkagsRpIRMoM3ymxPtmHiSr+wOy1Q1v
NxfnnoAvZXyflJ+X3MOGPsGAby7V22u/tZvAtBl/QK1Tr7k50xPmryHCYoSbF5PNNUNfr+4TuQ3+
X8e8Y6kqOkMEYPTxEptVVWUnZ5HYQKNeLNlyXSbyx+l4IZXwEP+XYmVLWdcMEyJmvX/6V/PjFuAK
Uchea2UYiGL7GmiR3KTpwZJx5tnmvxcI1xpAQ/4I3S8Uz0mUbY0Df5XZnssdB6yLyl5T3My+nVuX
R2OZl01kxFfShJaDBGmuuo3BGXOqavA9f6gYznQXduWEIfPZay8Bo7X+sVgFxNtuOvBgkUPMha2+
nbzWmtwbFtUtgznboEYZSSmasBM7ay6cqswT6nYJxLo/W8mKBuMHl+m0tpQF/r0mRn/ZU3dpfxiu
yBEjHkRriOMa3zheSjuKbmhR4D2af9PCyG4Amx+ldkMZLSeEcRogZAvT9TWVS798rlXJYiT9fQD6
QrpWD4KgzAISY9g54KJrHO23otZTo/LCG8l4tqx8RzypbjPyJE0rMOq6kfkdmf9F7ZHYGiB2/6l5
hJrSjjaq7xJJA39wllz3X2wjji1I1p8uiVKDJklsYtfKH7EBftLPzc7qqAatLYcqANkavQXBV03e
YQChk7hgvr/ZixL7voAr3KDg2w3nynJ4mFeVLTxWQmGeS991w1kG3RmuXcnnqSAY/VRUeyFZfCvN
KHDLrfKH1sadIDVsWwbxTtTsoJgf3kNqhhK7EXZPniH8UCx12eJgnMy/AM3lrLe8xs3J3L/Q8xWu
NnFf6LBtUdzOOiRUH8h+rwRNQnct9MKO8htljSkiAUun6bG/kO0ue17b70NC/fFP3zzAlYSn1q8b
nV0hYx6Tw82MpzhV3fc6yoT96e9uLJc3L/T8q9YlR0PQT03rTHq+gTR/GPXkYB0cpaQFcssDk8Df
1dReeffdHkgMBfTEDoUcXmPH9tlrSBmX0FzuXaYcrOXehcZlvEXUdb2DfIPRiHjqbQXLx9TBBOWi
+Y09zZwNH4UU14qUIpmyJkLbRCMk9UItD9W7Y8+QnIqGEpdlpHlclG3lbvCWDCqhG40VBoorhxJT
DKBMxhh/Km+NodrvHx1+LBLJHLnBTKyr0mMZ15Z6dx+0u3BCzowvQPVUJm62RxGqMq/fBw1zowa8
S85MH4z002aeyOmt/UaViW4Rdc+RVvzaohh9JSx+iit1CR+biJlE26nPztl2W4X/d073ohD6gXB8
/YXiq9utabL4onfDpnjHs0DOYXNHzLfahcDrA1iyrLb42/R9fTTB5BGYLrG1XF1TluN462lhoM5D
+J7nT84vVNb9M+3XcBYwAm1Ky1WCTYhJwyB2jcv/sVS/DsyeeQ/8XIGzf+649yiJk2geVAaiEM39
gBZyvP0biK9npR7xY+mh/ag4LJ0G8zjqqCZ7jg4V7cSA8rw0ObflZUHpUDQayVvfTnDpsvbdP9ne
RHRNMLqA6mf7s2VACUbrpO7p1hOGeUe7kLBHeNsCIIhF75+7KWdL73UNrQ0hOzOIMUr1C89nKYxV
n85QrOCFPgn0/NqjFlgdeqXfv7As2lTs5kldeNegjtSkAq2+jNMqavoPGm5CgAQZf3Sj31ChlJt9
bwPexjAfzmMz1dL925kl1moC5FXhomGqoH2Z4lC0+KCtrZbDC3izAjAfWAaTXuW9xd9V2wCMA9i3
j8btNZOxBgLLhcxzOWJKIWYPiEHgK4wqyV2/cpuqGXA4Len2yu1LCrFBcWB3gr6N8EY4ySZxv0Xx
G8aYAAojKxcU/Y+lmkH1w2pGmtXz8MnHYkCfG30Jov52Y1ob3mmOrUKMDlRNib6+YBJ6pkmlJxcN
fbyWVsvbtfqpzdzc7/rJesZkQEWEehWWhhDre62avhx0OuTLFy03s5wYcltVnRj7wzSoeAWj+2cC
Eb+6M7KnO/byKWwRmhPN5F2c4sjkCQIKl7POoEvNFBCEAXfdqEwy/inzZts4To/QA/aqeaxV93ri
Ubc3K01kKFbLFCxUE7eSGrJctIYwIyKPJwXemg6UVeTlHLp6o4/TtxXS29ySPp8CBZNFaDwcoZhJ
TfU84/rtTP5gdMU00JPxCGCTLha7Gf1XUVsXPsPiud3o0aPJds28ncqQimFKtoubCOqlWrlK3PGE
PgyIMa/MkPKELgbR7b2PNh0tBQ8viLphjTZqyr+XBM64H/A7DoUsLMx+N5etos0Jl/2/i/wFGzy7
rNP7qWJx5ZLFlrGbJGuTXJmWWbEoT4FTJ2IYsuiz5O+PixXSXfQ51Y2LpJEob0cqATdMZPFazs+J
o+xSF4tjbLWvk2DqrU8plZWVfq/9FdBYSOeSUQvf7ENFmvnHj9vAQjcuMkCbl5TZ1mj938dimqA+
GS/qiQ3At6uZORyUqzSmHzzA+SPQLbD2/PP3NlOALWiVU8dKvwXBUIxqWErdgt9+APdoN8E8cf8z
FnFeHZ6nNAPJysLl5+X9Dgk9DHV7nJ86HJGXP9K+mDmSAXQIOMGvlV28uXfo2Ws6FljcwS1PvTDF
AgAss+c6VIY69ckTQgivSuW42u2A/aYYCfOJHkfhsH3rb4AdPtSAtI2OYZJ4j/SOUWwKHYfmir/l
8M8FX9HgndsDGkexlkPF2dZy118qA/4eZ/v8Q9+9znnwU6Eg82/+2VULAnU19/VcggDKQ3J9n2Rm
Jo3byPCnx8+up0EhMSLT+DZAbbwWoOaRPKY+JySbqEtGJs1hom8FqyQIBKQUoUaEpiLat754ZvfG
E7OI10+7R2FfFTyOKfMDFqO20mTWzYa32nwQ4GiK2muuqO0wJPOlNZ6aohgwufiz460OCYKPLuhG
dTl3JJgGqHO+9GfEKHW0rzgIQcL7T/p1SYWpK2J7VdZOvHoZ+sLO+kO7AQpgZVbKgqgvzyBMJPoS
hvrDpy4ZO4hkm1tlVXtzIlXkmIlCxGzx6abjJ8RBE/XQ3PBc1nZZTFL7s6knZWmhw8y0f/o8xMY9
afk5NbT05ZstUXSopbZ45EBPIMEM04jEq6zalE8roK0vVypchXijESyXznGP7FUjligqM05plqbd
GWjrta+41Mn6fEuJKEGkvqvWASdK7vrWO2c6kEi5alrk5/8hSifK6u2YGcqr6hlSZ9cYKpWh/YuP
nj60NId08eLKxzZsAyxKeizhrizuiuXl/T1Irn4s6zAAGoGLoTLNvnbgTjjNXBFc0u28VRO6Fb4I
vxdlT5XCTupBN9tKqEjgw47rHjATAxCN71MoAO/7rOUb90XRoKbXcQwgXWp3hXtPc/MM34V8jzxW
8HoXm2h1+S1yAAeAX8RjR0sNATR4wYB7nLIcuInYK0lNlVO+GZvhu2TSYyL0RKn5u76hj07bqB5S
qVQdx5USfVRpb2p2Vdgju7MVYoTHKhfUVjhSZ2C/gpFu0+IJeNhVBTSxNSptnXE3Y6FxZFioWOy5
dEdlTg7mHZuM+5BffWAcoS1jiGIRYM2xgyY1TKUSV1HPI2apjqKtVBQovWEx8v+8+Qj9k62RjCp0
N60qmLtjYDjvstNBnKMxo2qA4rLBqdq5KNpNjFUAQKa0irbbjG4fmZrxAO3UNzqeUAvMUFe3hin3
OzGinCxsAIaIaDDFMEqw7v93Hu7mlrY3LrzB+D1EBAU9jA9NzmNcoRzv9Gfc8uyzvLmc3Q05jDwA
FbkkK6FAXyrI62/W96+8bqbrCR+BZz6rfwabxXIM0MANvP7osGgqr5PMnNrNwn8MWeJkf2NVrw0n
vEcF6r/KcwnYHwvFFLimkw/aY/OFnDXd84BiLNC+J0M6laSqtOc60MMvGiumlUoy1LInDdGMgoL0
wq9T09+Uy+61hvRtH1sHlo5wptjEdxQDycOUlw1xszcYtQvfiOfSW4JDeWb4DZKoa5mXrpt147yR
tbqDsmbo7k4+6lDF7rwn2Bf3YujxkuSuQiT3TJscw46u5c6v8kInzhmzsnAOm+Z5/0mFF4+Xv5pI
XwCrH7RRaSUaVlqTmXRLAAvtVicolnwXQeCaBvaSQJEZkl9TWFLKS/MrTj+UNaL+m3wH13jwQv/V
ABmn/D0jnkZNmrguD3BzHGQ0MPI3cKm0qujG7IdUlGhgrGY5dudlBsLUo9IlvKELnFHEu7vC9V/Q
LrHyF5REURr0ORECi7sxIXa6SATGQLH7jIzI8G8+ifcM16VV82LEGvi0kPm7Ej0IDIrQHF5QLGzV
GvGto8sXEJxuN/2qxdCOsJ7EofLtDKXbLJEGxwcGJPbJRg3oMRbky/x76Flov8vXr7AQBqRRkSV8
nl7yml8a+KKgar1oNZ2pWCi2iFa4R3QdGki8AK8SQI/5H+UVPL9RUAIZ81boPck8pSW9MvdknHip
45GDpVgq0aAsf27KOFvYZtwTqnisI+u9bjzfHj+Xus483S+Lude6a6sJCfIqVaeOmfgyXktZ9VbY
lRBizSEjNnGKPLCiHmCHuravGuntJ7luhg2Wb2UZGedipwDEmJwEeW5fovh3mNmvmSanq4cRjWKE
9mAcXeZxlvuCrYpfflO7YKTndc4wv2PVkrCY69ydJ2LGACdlUunNOFjGHIol5ZVX7Rsq93i2OU2e
ahki7F2a35v21lNQ5bfxJvtM9c+f42w6M9rKd1/s2aJyKXcn4N3hM27r5qeA2dkQYNCMrdpmaxWS
zhMsK3Oo9XqKqzH0eFqCveEbUajIMR9iLeJvekMin0gyuyiPO999lME9jlzcefxfkPP5AKB/ujj4
5Gjmeo2oW9gn6eMAdvWEosEBD9HqLtmSR2XqK1sxicybWifJIk0S4Gjt1bfgMiRt/dWYK3oILJ3y
3+9OkdQjkEFsyiy4eRqCkbDdhwpNs5Xjxdvnsya7IdqeJjd8e8IRliJTyCGvEXk042zM4VCAygN+
dLy9vuoNw/hYKoQjxuK981YwmP3j//0R7cUQodq0agFb3p9AbXu/5/KAL4vSojl5UDusNgP4WR3e
eueJ/0tQ1IcDLf6CCWPLWKQM+tPeh+9LYI4vaBa3N1xUaEobPkmGgOeMMCfvruhPnJPePADL1I9A
IFoUprRzwOG563RGpMDhgyNciD0WmXWzTsX+Z05EKgZud2farghzE6d0q497bhUzxB8PHe0sL2IZ
GL8gTQ2QfkaDnFF9xkPfL4yK5O/miKpERtwpgzBL5f2vay/X3V++SIyiAoWEceCe00U3eCDLvS8Y
jcnwuM9sWzQFjgpGCyllp/TTRfyn7zib2BZQ/Tk3/zCtH4Kpd5BZbMoekjVS2BJcbQWWSS/XeNMT
6KuLUSktGA+CoQfR8S1cNpotiuc6GbVrPI+Agv6D+X+rHgmUIXpwwOJgHGMMB0shbpVeIr6ID7LQ
nctFKWRamVVkeBHq2maI0ZXvW2EnCmoDjmUTMJZi9t7/EuorXm8Gg+rtK9VTnE1/7eWxPadLw4Ax
CHqvr32WIGTmpi1KUEbLy4r7DSqlx7EZd5JREI2zdHSILx3SQAxap/ONPyssFOknzQiQcwyB7ZF8
5BbFqV4UNmHarNWOpdTPixTqu8ybO4ATGb5OSnfpzBZ4IvNu9uMiXpjOdZzVkDIiTBAEK3DtZYWF
r4j8VXNmzu4ZM1JHN0fwKLlt5vjeCzcQEyyXfziyMIzGnktwprjde8H7q2TE5BHjOS4Mc5VM1WEV
jeJmYQJeQfrNEMePPULqPZTPwDhIC++QQQtD6wfz8PMaEiiTuvb92WVC+NwoIvRSNUG8JDx7ME0v
gik0YWqcelRjYNgEja7XzBvhEjhZ5wch7Naua6V9WnB4lsy4dE0DuTGLw5DENSWQAtYHoiKSSS+G
SrY6hN07BcKOY6oCrtmFg6uZ77fibVaNX4Ase9zV3fpKhX37LVEa7jWkeGBN4iofq5EQv9lEHuBU
ttbsDRWxgP4A8qKfNtGnZ1cvw5X1AQY3hjYabRXfJ+WxcnBdwQNI1+73ffbMqPwLag7SFEDDKFf7
T9O+nrY2sjntDny/1EQ3Xl6jJbel2L13ZbPsJQrwixxdc8ZVXARi0TFx7zgw1A246vyKy7erMjzU
TmQwCNcn5su3VNNoXidvMl/v2vIU3/tv+dDu4aBXodFRZVByqh1r0GXiAjYofh0PbF6/lp/aAx44
6t7ZPMfXzOerjD3j/8C67SOIdLkcwDhSl9nxhkA9uW6zcq9FmCaWqrx5HEXZpBVhnSRYsler3xRQ
aTPqXuUsFqMPO8FMZR5Q3bMLZNcZ+v/C6rqxIWTQ4rJOm6R+gTT37mh7o4TLAk1ejB5TexNpK+KO
uLDtJYEjC1U/CY2wVuCk0CrvPsEmmamH+ZrYAMkdbUxWYM5nkTpaenRY/hFvlkF0xfiC3l7dxb9A
TsRS46cO74MmeeEnUpdoF/nvKPq9msQKK1TSV4YXOeaqq8yQvHd78aU37Ab4kz8hosA0W9ioYCca
89kGVj92mlICWLTW1WcgOMgvYeo8FwG2ZHJ20IsCG18vjhnKPG8LWK5eMdS/udPt0Rhw0n75CB4H
cRv+IfpMeFdK2WKScj1uR0jFNYyPQLW5no9QorxtCxU/ftSWLTVoBkKnb1IQt/7sLhdT94F13NN1
qnuR7OlFwn+cDZ3ERwWuHx2Jhi0v282WZpHeAdN5y6FyhONYn9c++6Kg02NofUMcOvkAyneWBgjo
eP/NpPEfoZKxzmSsGFlS+Hu21JzISdfbVsnTSln4ZhOi2Q/26MSFvq5w+k3bnUEB7bLr90S/WWqT
cPnM5ijXC7O6nGIL1YlZhKzo9nudvDvF6zfBD+UBbAKF4itdOM2Uz51nZiouY7eX97EDACW1g03A
23d9H1OgxfZ7xjZbBKdU6S+5ttBu67mF15p49epBzJg+KZbY4Ly4CCTJjQS6BOtr3FeRSCa4qaUe
LPA/0KMSJGiWM0b4ha08zEnD7TXRI1jF0x8mZyl5pvZKWyxeiSfNyewD00SuA/2/DFh6+JoGRTbP
5DNtF2Xr7l1e7J2WWZOOWTnDLPoAJFFVkGIFYR/89+Wjr5Ouh0JlYg/pHgWRCadcO0mrea/Az0Fd
4vradhU6iQmdUJvuXxl68aiz9UHUNAAYFJIPkprwhT4cEMAMoattR8ayZU1Boz/K0Jh4o7azFldN
eWTjF1Kll0nYV4rF9YAf7sIrFHaF7vl2NoH4uq0CRqrME89nxMew/Yx1fYSkMLrdxmfmEQqhx21Y
36XqjuVyTtAXot9HwVmwrGngrep7wiVXnBKYyq2OfXBRNopvIVNsb/f9iNnO5XE36gh9dxJXroR/
1hk2cOX6KulDFLIDGWqOtiezisexcxn6bYgGCEqglV+VPUTlYNsFG4uQKvt3xqvmy9fgNGCYHcJd
eAVmVOT45d8kBvmkMWogotyVP/z3hdBGNRLUI7SIfHR1x8czNlGxT+Ny0a0pEdhJKqPiDxq5/caP
5FWxrrJyo7ZDsbH7/G0qc1DedGRfo1h2KhiwxCMTZiDBfunWorjf7WyZ5zeAP2gk/2DaRayp3Ehj
bgBKm/MsREu+CThqj3B1c+2FKEnFNa8IH2HnwhOueJ3fMrSbanyluXPd9/QM6Yd5lrbMqZcOzR8w
mqSYcVAnOw9r5vJKPEtyDw04RIUFfpxA46N0GMtDrDSNJruG8EEp1gcqVh889DTQL3dTq4842Xll
/C1D8Orcc0XWNPx4z+V4mXaI6PZMsFgwE1lG0LE4BKKSCKavlgRRAkJU/FcAbtwo1G1Dzq57xjvu
+QxbcFXhiI8SVceVQ+//RHEPl0MP9FBwc8+i5dk6V2XK0Ry6JGiOZl5tdBNHN6kTz0CdD+PoQLoJ
UrrceeT8QanSFEXLOqH68M9pQp/INn+dLQH6tMy3X9Oben8sxVuMqrxuu/SjEJpIorO6qK+5oUtT
0WMdZcnMQ7XxByiSWv1iXQYgkbfaWYKBrZs9aIkr8gTRIWF6uPN5EGAMZKPC+rBiK08AbT2n0VgE
n0atupvi+M7clUL0svXtun9eXqgFGLZaVdAADrT0l0xxo8Wi2Q4nmrjK43WBD/pUjE8xjB1CrJLO
ScWVcaZN5PXROcJLIXfWpEVRdwPf89n2R0BWxi9w7eVFtCLwIEcrfKiZwGnanu8C7WGTeEfk/aS+
xSH/bahmBE3RhjPrh8nHntRAoMoxFBB+jgwllXRDcUWQdSaj64TqvInFJ1ZwapcUY08xo7ZNopqe
JAxUJVmFAmss0PrVoeZsCzAlJD8bc7uzyJLJsa/bqSelCMvhDHwvwFAHLRkLMk+zdlPmmh7sE6Cx
t57u6qVWhT1N59RhAJPU6U9S15rjVKG8WpaiP5aeikZH9NKnBn4doEqSq5ZMrZxGSqB4UELNVeE7
D4qdcahJMfPW0MMkatk5Ka98RfPfU2DzYYjxw/04m1Wmo6mlmB1NFR9DEQ/hQpS6F8F5e6iz19Qx
HhdswPCUKv1c0xF+6AXAsrEHUpoqRP5Tf7oir2oJLnnhQ/rJ1PAhIeUFM4h/kydsmW+lWPl7osNS
jg/KlEnR5WY+VFM6PAfpG/4nP+oYlUWDLTH+2A/DVGmtB4Lg/B0qtv7rOnJkQziEidLzy9713mKQ
bXr7CSIbAU5e9cvg5ulOQudbk1DOYNpx/bsngI0UfTbevVJOCTjrSsm0BcOk0iOBfxkKKmyrYCMg
+T/rwdSiHLGqed/RQRttFopPqJ0sPbHEGiv95hjthFBsp8TOi2roR3l3jnMeVTYEPYMty7B0u5xt
y86vAcoGpck+8AnU3ZxoaoshMXLvissS8AY6oqa3rW7C9Zenbo6d19Z+rKedgi8TRmAQi5FLrAht
kG14bAQYeeHxlOxU8slzcKTuGFMv/SEwGvzMgC2zoubzdfOAyH6u1QEqW//guOOX4m65fh9LOvMa
RGjYPYZRa5ommhAX/ddx+zEDYz0xl6wxR7aw9v3g32f5ygKeJhkm53YbdRYjO8M5RuErvLVrn7M2
PytdWb5gm9TbZuucWKWh9gyOaiLm9UruTnyID6g4lvsou+90jc3ar9atCjL1WmlJyqLROE3kHYkB
oPSDL48eDZKTaQYYCj6SS4JIzLEf+FucyLKB3JMp9x/kb1dSImaLD0ZmrvmXQahv67j/gytrywjm
EVC6Iq7sgJ9gdf1hiSkZ3AJY3b0tsaGJ4atIT7IG3BhW5JH3/xv0MjBA9Z5H0mtsc0bZMxkH1Rdx
uH21BcG4ycUhEYWzSIiwaa17ZkJCauL8FJXwoeYEMwG/mN45Z0Dumku+eKDtRwUJ3ElbsMZPVYpC
aajuE9bxYkR1Cu+kIT8P5Pa6eNgqTJvHYs0WHLep1Ok2FVxzGhmGgUaQSqVOR2Mi5fFqs8uFyAgb
65lrJF/EKhpOPk9jOjMkE/V48RKgrwDwyDgZtIslH2xasxvEVYlly2g7Bw27iTqRmW8ra58e61br
pJ11LbXa6WbRf2UrIj/bDAt4uOSHheH+o/IJHWf/AGaPli5XxHy5pAGP7wAEki3kb3H5izMVtfls
52zUx9uouPfp4fQF9h5XiQjt+4XEbaFwcVhAZOuLE4fok205gEQvskhiS4J0XgwyGC41dIYqf7pw
fD5+VDXz8EF7bpAb0X+6LiXEf9oLG9V4Qih5Ue5Ed0Hv9mNzzrGdMkj3vYtR++SfoO1ucfkQrL5Q
LvJWHHMLP2Jy5Ds2oG28d+kNmd3vewWJiy0JtIqtTFnM7uZ+6jLSz8LwLoHSRrKdqMNo14wiUhMD
HtWJC9ndhFYAjQlMyaQ8jm5/DY8kyk9bsDM21P+WrgWZk1M6HdsbUySe2MMXQ3+RZiNedZ/JkpgT
yZtkI/c7fNjJJlSxxFnNN4/aNiH24L+kSJjgDfxPrAbjf2mPgplkhXmJvSMQ2CLkUGVH+xFgznnb
npyKDn8TyoXWpNm53/49WcD33FYG7lhnge45+NGzvD9Y/k2LSuZykuL4NjiISOURqqOkjxOvEhKF
TB1D5ijZ9WAkrvTa0w+zpvsyU/Z74fMmOyTbS7ngMs7Gvfjj9V/+LSGcU93Pa9Ut6QHJG+/9v6QN
ByJgI4fOKOlQkQc9R1AKm9GOx63jDA4VQ3T6W5tDWAm6EhhUw6f1EtHsF8XjYE+RWGZO5WB/uVbF
Bf220vv9yWGt4q6J+ebFkJsShBWXgRFwJVZQtGsN53vYigZ0mLqj6MwKs2ecHTTP5UNyb9d4vNyD
wzgchg7DXLa3tZrgMJV9tqHu7o+aMWTvgz8hj5cqU9PxJbgFwh7cM79dRvc95Fc42YWz1N815O4t
1A1BlhmZ9hjPz3utUwa1Wbh8rs8UnGvB/89z6PNzYhsBwrumsBwe/q9FWPk13yZuLnwaEAgtUxiA
nFIYkb/ChTSlIUGF9moKtkQ0n8NOb9ota/wSrfWJopuKzkuUmXs0bFsfMSKoKo4tPpN60xyH8pA/
EGMg2y3loLkmNHBlRyJu9sjWd0oJ8lIRlLbunOSRrTcCuagR7Vxb0LrfhxH+1ZlfFweylJ7IUe30
CN4spx0LCNNGAWrL24y60/+qC6Cz4liNVYySLRabxdwOs+NdsiAhi8J6QBnfYQfmuwt2LERX+WYo
Mr79EgOVzxBpvK3fnrhmA8uYq1y3AEFD6XJ5hv8JiFuQMEoGGT7v1jTR3gUS6QC3/GecmnMmSYDM
ocusL3LOTguwK8+VYyA/cFFU+ARfMS8kvRUjqShMAAhvCafhgeyxHG9X9spHmA/VP3GdNTec+eU7
heqPnBCWrjQ6SY5+CjYc7Bapt6BFPSSuQE8JzE/BWK+fQHfogieyw3q52HbxS10RpfuGGoSyAk2l
ufFPtWYm+cKoaxe+yvuNg5SqCLSKSeiOnJNT3wufJHCxyKnXj2l4ZU92VHL+wHrPKatUX+C5peZZ
kvKRYiN0ILSMXH8H0XvOoZcvW0Rx0TLt7dZ4LRJvvN6eqdX+s2rVESnWErwn0e2hjEJ/AdpnPyFg
sNaQYMwMwZ/jlWk9aHq8BAl+twLm/ydMF+h64geO0ksTc7ouCAlTxBsl0twDzU+LQWXWJi0F8eud
UlfYwi5IJWbaUULXOavQxddyTMdY/MXT+7OOcFznoOA1BtVjzv3Pd+QSOnxop9k64BOLkU/Uz2F1
Q1yoA0spDQHYHXoNo/S+v6tTm4Z7tc5mF9mlyFNoAQqeMGKLvH9YVR3pE17dd+i4XlOGjs7a0dMk
VlqoA0GNrOAz0nI25fhr9157tMinHu73loUdMJcGeDoXEaIdICAJ9l4bj+mTuhpD2iTNNAZ/rcdI
WZDrB1zT66Dr8KpAC0TKSzltiTad2Bc49GYrprapunRHOVYxl/df8fqrNlc9is4Ci+lq6zh3nolZ
mSV6EaksDZxIGJJpYh6LVjsO9pRT3daGl9cs/ehXeAP6g+rqsiHMMESB07A85BoHhF4r38ATlBic
P4BECkTf68a2iwFkL1Rei5QKmaFQ8WllwmX2Wk4Bq/voVWSAk6/0G7nclCeRzoIUN8lXYdszbBIm
a0aa5H1rA+NQkg5Squuvowz2auzhdPSMDAfbICojLqYt47kriLtm+URtf2pjzSu7eUxrCJBrTyBZ
qMcmgZEmi0r+wdb+eDLZqDLeK+fEsqWXGH5soOgNB1Uo2pCvyu0iYIa/NmjApz33o0N2tq9oypQu
791X5KJKw9aXypWbfFLVzvmVtygkuHUnFuRwFf+p5g/LAka1mqxhwqHhy45tgI8Uc8fs7BDkTsUC
a2V9+2IAl4nFxFWDYYIB4l5r38dNCulB/4kXkhiePG9cLMJpzuPwsaTfQP9due7CDdKBxnkGK6jz
JszcZW9P6+ObgF+4NbLlCtjZFk2bo8M0t/psNff+7cZv9oC4QBV1RsFn2ayFLMMZFBNLdwQLxFXy
Q2u2o7eAwakWTGNZXAvTyDmFUwJliDhcPtlt5r5eltki7kdKoSuUineoHHLr5tf17U1wGf/tghPg
R3mEWjc84Y3x6xneEOSbbuNol/wtzJLXJ0/DaQNzbfXSYKhinNTcVBoqz/AH2lU09776/iCvUkLm
xbhEfVdAvS+hwM+YsDMWJy3F5D078iCViW5E1qkI35/jd9yN56fLU7bsCGRyYwRY1IX+Q84p0Df7
jmcuvAhRAmnVqjRG+noJ+hEp/JHuuRyBCFdPI8lyi7OjZkGcyjXjWrRHMP2C0/yVrVw0AE90fAgG
OyTEZ6pOJ1f2OPzZOrPqJpFY7ko+Nqqo1w7s2jHEj4OhHnx/2t1WqtsSUshVaFUQRjeaPnBqzStl
C6oy2BoTMqx46Gskth6bu8hoj/xK9cLYFYmCY4/gzDJ0rk7D+e2DokDu29axgQp/G91NXyHwqqtW
YNMqscbI0orGC4DOKWD3jYQ/6rJ5/skLWt0XoRHll7z8DUkrP5c7SI5V19avGv+Zl6mJzgszZdP0
phP3EpqmU2++BBcyqArLc6HCQrDU4o3N2iSi8lChA+WVAQlBNWHx1zsk3TTkx5VwqODshz1kcdqX
dXBuqx9Yx/g4HMfB86Qd4BDcu7VjmQjol9tgC6dLaH09mXKCbkfp6N3NQ5OYKuHldcZTxsEmGwPd
6+yiBzg2w+KmRNC5OKR5tsUUhyFUZkmMTPKSQszX8ExXbdVJxteuSEyfCkpn9vvI/HQXuYRnd1OM
U4KhET1HHoNhK65cx4p1kzv2sBWv9NrTNjPYdn/DDBJXv1n7M0fw4ntz4WLmddvDLMRxmMdbU8a7
yK7Q0pncTUQbYFY9G3KRtcbgnlfD13lYcxZvjd8fKtKw7F7UPYosKNzCi7r1+cyRbKxAgpIwi68l
SGQwkOL/8omOPpl3eRU5mX29bnit+cT8Z4PhHijuOw0GIF4/uN0/nPGVrLNTIAmw48LqtSe3LyQq
UXe1fokNLr/PmYfYPgUONs66cxsCdIDMIGtXjrrkn8KkWvrhg0AWKdRxtuMFCtLDN6nhy2tIxxsV
hLipm4zIdTy5/A+9r2okwgd33AzUsE38DXxXDDdUM+NSqUAOQBWO+Z+r5MEh/A2ys84XGUg1/qn3
ptHtlu3tuR0SPbHOW+uN6XvNcAwhF99RdDcGjpd8GVdOIzpUgDdl52gcT4XYA8+GUgWjWJUe0Qaw
9tdKHtip7P9mvlHaezswLSejgAaexjv/6i9aq0oIM1S+uqtPxnFo22VgZc9lJXxuM/xXeq0tGQOn
ICB2TrimpPxoefl7ZS2j9wRxEs6WvFR1D7ba/Ze3rUYXCTr6Rb6lXda6SA1BVA/4YAwgVIZqga28
EhSDuLEFXWdqzvfoNK1wkrWDWpasZB2bvCKQ/hzI3Ha/HWH7hgfHPhq7ZlAPuEryo1cjYQtQQAVF
MH2Vj+JRgtgh4qqMECp/fyyWwMDJI1hTc/uju2dcpIvkz8ZiHexYbbDtktJjUo7HHUX/9jF97Da4
3p1/Jz57u93QZgRVXejsSs7PJIx/84o9K1gM6++po4nyih1CALsQf72ECOTtqGbichZvTOZwU81k
sPT7kukoyr2EnyWBq2qCqgb3NaTH0kHMtD6NTZCWGSzGSvRvaXLTXhLn3DgiEu5LYeLwY+xJPKav
sUx+vGsiQul+mpTgGwsrzWuZJ8yR96LuhYk4ihU9kosmqRj3rmTDK7mzgFywPkPkhvE213CQ7Wy3
aFtglKPdcqnwYZs2zrtYx+9ZkpYOT4y4cj2uXb3LM2rQbCaLkJm/vY+quVOvP37MjqEs9Kp6HZON
BL8wKUGa+oLhq7apEPFPDZQuBlQBuU1wY90VNzHcj/3Cm8cdZecujgFC2KK2w487gvmVkPEbVn7/
Nu9bWkcN2yB8swfwsPtk2BnlVmt4W6mvoSSFZAcpL69j7iY7FRseORFfIl4+U2rXZNVLaGQE7ELr
OPzlaFqn71APiFPX7ncW/7RRGd8Y9KHJ0+S1jegvD22L1G2YCN19v9JUR1GgpeW13/4fOvTylf9i
BSGC8Zr4BwvlmfB4pYx+EKTTzFd2ZUfXWPP87RCqdxehcTpkGGdy5MIL0ljg+gteOxW+uq/esA7c
CL3eenw9wV7N/MLsVE8yKPc1PPARvgljRxg7ChCX5fZcknNdTqkKIExoYdm5hkxwKK39/7ge7OAy
s5RqzNRgl5FmSmoh8Rd/k/jWizdtdGTTF62l8wIKOX8nPxcCavRimp20AOB7eqp+jcI3qM0MSrv7
eRVkTKL6pQSQnDPqZYQP9WZntgul/pko51pNcQBc3xOrv40TyxPs4LLXLxP2+Uwjgj7g1oLk7tMP
njPOySmjRNIwafksmgJCTvq8/UTmtgy0Hpdv99S7ZNVdMciXQzPRhOHCxXasdkL8MxaMKX/vuQxO
/3vyXy0DqRgso8lJB+7tAox9WF0AV4yimWQBZ8z6hjQQEWSBIPKWdfpfJU75h9fAyKZ0JLFCgp+j
/0XSxpPL4ehxNRhr4G7lcMaKNg3gzA5+i3Skya+Jn/q/Hsn1ct6RteYJZfYXAkti1hOM8QmpgH0g
BuiHCdFlYxW6ThPOGevug7QSdPscjU+6TUobJIzTyr/FfShX0l8S905hKskZdfV8YvijPPU2D3LV
uZC/Q48BlmlgPyyvLlcfH+1lr/aIfo1Df1dGo3ffjrU72//TUUpskOZWLQHOl2Vue5U+CgRIq5U2
Woa75Tofau3B5dxlM3D7U0FLtSa1aNJfG34G/1Ox2xOD8lKLlGUr6N+a3WZay1aOWtcWReFxor9G
W/dsj17p0r1DkHKGkib57n2FMJIo1RguPA6l4ubz6HWbIUpO1RU/Y1ztF1zEOQ9vuwUa+kCY626c
AoEyQdIG9T0xhIyZdendxaFhaQ1wm0cedQOeu2TNfpjZnWui74+HQmU3I+3+3dBzlsutNoa1ieiW
aQ7Y4/yr1ep8g4LRgVruZRgTpEAPaEGG7hB04lP4B7IvRqcJ3OJ7KykP3JziEm556v0CgiwZeCP9
q3K6OFGQ4bOzT3b/Dy0rPLElyQ5wByMClV5VwgNVh6GMMn5AOuby5TaUhfQBMHUDRsCKogJgNuZV
L8SnCNxVRPhwFDilJ+qsYn+fnfzW65JqIvdDUEqYaz/wgxqrIWTLL1OGCh7UR6f+RRQTpwQqyBuV
aBEzf7Lu+7rgNRJE+cymDOPlst8bB+epbj19EyzumuczbWimVEv43+gUCdHd56+xkdl1q4oUvqoM
TqpI1VSa1FT7ZNBpz+uWcVrATmJHcHCLurJL0urHmMabck75+4ZbbsdSi/BFTulYEyIkIVCxPJtY
RCVC5RFxIP73qNNXRYMA0xh0ref+j/TC3HInHE4Y3Qk4UW7W4RZA6QqeRACDDJzTZvQxcRYitEYc
qnRR2KbFL9zMgOG3C2c9wW/By8wI2Lww2n2eKuWlojRgU8JqyoR3XM0LtPR01nwnOb0iEIwJiQVu
FKC99mie5LIChC8LUI8yYylz/LEqUcNPycHzKdxiphdl0ltBRdvTjYseXU6F+n1Ev/eyRLWVWPAf
yEjFyHFcpukdWE9xTZqPTuuSsmavZ3++W70QUG5eN60g8F7IVlvXqZk39F3ZsW0zmJ7AMvy8Oy0E
97SoV+BqLxwL+pUPf62o2b1WVCW03lIZjsLF6GXsYjBvEBlK4aQ1436GLZP6ueVc1aXYW+1QxW7m
xdUzm8aT7mmoEuERlYpyKdSQQMGQfZLk3vCjqlXA1r/NT7e8gvkFCNoCNn7Efj73k9/iC508Dzei
kM/aI1dVAME0syuS8nazikPNJ0iAUnd450L856uvf1Sh6vxMTGkfrMVZ4X4VlnqvVGI2RbV2IyVF
QX58n/5gl37w7RvS8Z9Yi96zjdFlj9MxZAdAAvjDMHZpyIdytOjlEfXtirY4NDLKU0RTngTUPCo5
AA/7k86B6qhdY026kqUXPriYve7w3PSRYDWCJcLXjbmJAxsPlrcC2tWLnztNS3bKkztxy2UNfi8/
7mt6/KGOl++upQ/4vXotIjAhxwWWdfVdI3ESZERrqlUMaKdvs/cglSw31OPNegEm1owPfJUJDWqK
xFzSEjzrq9LjynnuKPBvzuFtW3SGl62vgdYNhIBmxO89eI3DBryCFovmT41InjSfxUf8DCRBCb6U
yF7ln+znAWrBfmWdc0Mw8VsF7ewSRu7bSIOO2bxqM1uNgPWUWovfmorzAP6nDQmSVHGfYGCr0fH+
DyZv0ruF7sXXVKgLHVkaf3ZMmfb4e1+ihA874RIR8yxWPbW+ax/cxbJOOWwQM4+rPF25IVL1OpL3
ezFC8M/Czgp6Zoyf39xODKuRFho0NgzKtWvbHVUan974uwBA4ibKD8hna4/A6jW3Uc+eUxhtVwqB
KPzQOMTLrDNwGMXfFPQ74n0eO6KD8oa8hzLwfohE3NP8ewhB2DWRa1UXMp4Ie7X+z2CFepgB6IeI
UhRV1/O6V5K/PcEklJq9H30m42UAlvJkXI8A/C5JaWOGaSnkNMM7yP6Vue/BtnBSuX0saphpcLor
2kFit/aHRRnuz6Jv51MzJQHp5pGB16c+Qg1xxFmOlhz4ATGEzFa9KIJu06FHR0UM6Qf+nTHl9PKl
4SeLTAKVQP6QJFv1rWDCNMdIR9HTd1yuIaE8yoDAXTDHzC0FDVmDn7U1CeJYoAtx5aNgs9g3JATI
Wa9ofgGonzmR3jZjDta7Q3RNP7e282DxGWEbm+zXgZJ9p7cmWYY2TicB1HQ+v0ACU6au7Fw6QMOy
QJ3sacg+h637oGQ+BsjDij76k0MkABtgH6OlYvg6B5RGEp9vtv+Doax8m4qjU72oKcTHVbgvuzZK
N/eo0uy08zWf0Da6NzSdiPYs3HeZLiR5jx1J1IaizG4O+BTI2rDc6XZSwiv9fAxR5tNmwqgi4QBl
qPFHK4BfWICqC4MGwN7hYm7Zq+/1RDxZGxsrLUOka7DJZRTD4zXx9WFEcPZFUZL58Mt3Hbm2NVXZ
fulq52d4LcmAIv1TQ9iep1g6t1oFmG8Qa+I0H//3HQqz7rQbj9RuO13Ir9GCDc+dK/970idRigAm
gKeAkY+3ov85d1TP+Dop0oE2dQrVgYQNp7Elvp9ZLp5oTzn27XO3O2HiVKXDDjIuhIpgmFYVo5Jd
cilQTTar/n9+E1XmVGJUAGdmuITCmqYp/9ToCIOnPI6wVvd8Py+NHvuyyobZ0TPTyjnXQkc5p565
S+/PdVW2sMRMrnSpH7WTfaDfyxviSX0YJQ9rPcvqwas4PAugfOjfB/2fugh6WX7XIFLlo5vHkTwq
SUFP20KVAi1tIertjkh8X2ZiSdGJe+rK8VKcJ63v7lTxqJT6b5uodWstuyWPh3tKbhdD8h3DxVKS
85zj2sEsxtdxj3BAZr7jVCVXCfC7T5uhxtuyqMdb3OtXWdZeHhiHuCNgfEh3fSc2I6Nay3WI2kSp
TVoTvJRL7+FWX2J5MxB4PrJOgR2IMbjMcDR8pQWxofzWH9K1dMItwPvEhqspK0057sVleon/Mjd0
kpfLZCmt+p5muP1xZpbKSYQLVt/u64SVvmaGP5qf6LMgQOZGO1R/gJu1qkhjEH2P/jrCqCsUJUoM
rxaEg4xnkRjfdYMqzsqbRXAzQ+9XULPYXXiEDXzWuhsQ2t2ozjNQWGBtCY/3oFVYEtZ5mI/OwWMZ
FR95n2pMbOKKW+aD20qhs77affrt27+TcWgKocO65CqubRNIMwuS9tUZIO2o6FPrzt0wBU5VR4lB
rMNJR+kOpcK9wAV/6kKy6nuk6ksXQ+f4UXK8rMz69ghyyKIneP7OiW6f8Xl6aaCI8Tqg+BLB4PXv
2ikKb7nWbhWoo1G63j2bekwMHrlwJSwQlRGi+9T0Y/6+zsCOXAVM2IorKCtepYfQqyZMVXtmGPfE
osOqTAyR2RXaAX3/22py+xK+HuKOtMktFo0IsAnLIg/R1ir0U7naEmlz0GPISCcPltAH438YiOkp
k2oq12ZbN/37POfn68WAGTsYC2JLRAFsMxW9SYuzg76z6fTdRj8bIVunsFJjdk15AekKtLp/Hdhk
7/l4omezr2MeFr8yZs8AwmNJ4M4Nv5CvA5yTQBvjgOn0OAgaGFXWjsbYTklbkzRFm6MUBBcmsgBE
y+kttKfd93FIa1f9yYvRF59MSL6uEwCRBK9LwzRowE8SW19NibR8k5xd3JHyytrBkqAh+ZesZezH
HoLLEV1LrfKZwb8vqGrUFyNUFSJBztIuAarhHg+Y6PXw8tJRTFXzI4S7X6ABuwAVI8SLEUNUEiw/
ewDDmvwkotcOYf/kd6AffR2y6Z/ywZUFys2XVJZff/XrH5a7X6JDfMvGUwLvuG6VkK1SWYOWXZQj
6Cbxz76PDTUoJ3F/I4dfWGjl5/aDgP0mIJtpmeq0ey9Yc2E/o3Q9tyyiheLsPoQPpJBikKWz/oJI
VcNfSO0IsfD9Ko9Ar4vcI0rLnk8ksE+1lzMDO3w6D9O4/FAlaIeDWwDvDHK0Fceu6s1Bh9KB0hb0
E9DHi3sNOGysh6MJ3oRkx1rpAzYXip4fy3sV1tZFt/yZ7d8QRl8Oj5D+dPMP/8L7mj8VvuBmm3ZO
MahHJCEyChcFpBsxCdsPYR/dtyqFTdVbHfXXD+BYRcakhbkc7XrAu9b2QenEnB1GOswFrnpjuFXP
sDcs4Aj39WAa19yGMj30keeFj6FeoahYvJSRBR6W30xjY2W29y+cOFZcSYfNl1zTSbiBv2wgz3nW
PXLa7+bcRXz6sJq1B09fiGy5JNCF4cYe47WTi7OFDKAJC9Fg/3f3IOUjxlCFTOYXaBgjXHRirZSJ
5fxPYyJZ+ta+T6XV1zxaChvyjOLBiYb4w0stow1k5fMDPJT9m3GabiZ4QuLpM91CCjQxXEf84FpU
0QcxDBIg8eiIk07WhjUuwMI1VYEonHrStPGckZaBJKZmrqHRbg3tA6hePzDiMSH/87PysKo2oDdx
DBnpdM5+DaelUTnDkjweePzJ1fWV4/jKteThUmDOllkOhjB4+KbLP2EDVPyipAQElDU6YBxsL03r
Aj8e/S4QWFIb5KwZccspkq2TKFEMF1a+0WoCLp56C3CHFEiF2YmGifsOq9FXfQ2nXEaw5C9rUVB+
gjesVSKKQ56UwMj0S2IL45DZduQ966flHe6TA+RXcAlki72UWpjHPCsHcKUMbXlaX4342nx5Xoet
gJBHymqz8HwArszuaQ7Dq6YtG4K6wT3oGzcbDHmzaGu9VuB0v1xq4pzDN41PJ+77euR9KkcyY2D9
NqZUl29oKK+5tKjhmCeXViPudP+TwkvFgqHzRXh5ht2ZKLSTeB5fBmEs26Edjp9oNHEJTuPLZCDn
wrvOyvan4lLqJGdh88X3i01nAdIVdM3N1/Ttj+HNI7qQowQIZg/gR0NrMdv4llUH4YSyw8wzRtBN
rBS+6gOaojOHVcrmLkb8NOZwsF/w64LN/dzlt7DRCQRL0gDnmrWhYGpbgYE1vxYksvZBsSox0QEt
fI4yPeTGDIpnNf8HlEH/J1ExC2pbHrLKeumELwy4NZtgvUiphImrlU2LBBYm1aJWpiIXlzQ4sMU/
NiX/WrSLA8o88X/cMwUMCU+3UMS0W6ZpBSXxYYPrEXy9sx4FH/Lf0gta71TJX25sC8Cw3LbC2/Rf
4GCnqnvU9Oj5ZlLl6moEXju5RI6F5oj7/Spn6NEW4o/TrZ9l6F+N637c7+Xq2jTHbxbXNLdbQBzc
Wk2tgZzVOqL3cQoTXZovEWqexmwcytaeRaAeV7qk7HqxLeqgpx3OYm3fJ6SgXVmJrYuazErCg5Dk
kwNIxGyPd4TrMqHMVq7j6dZuJfblMxih2xcTufz69Pfyovwg2NkmdKiHEm/E0F0iEoQweF8k/YRP
XiODDj4WDgAf39J0eTPba63GcaMxDzdahnGSJpJoPt2gP1IiSUOKk9lthpf2XS7KWe4rdB5gHA+a
1qeXzdqsbhK1xYi/9yj83GAsPBaXX1XlZHWvG8iHQlcqG93UWsr/Ld1w8bBn+dL7Qj+PgZv+6Gmr
2LthjYQEdxp43fPSz2XPrJ1SR7Qi3/o/FtZWhA4reqliV9vsiCb8U8Ay7nnoqG7eZatATV0PMU0v
niwxfoGYQeRlb7ypD1TH/gDFpvKtsv2xP/eRliH8PxTIN+yDOxnC5VZ4/yZLjXUeZIBj2pL5NJq4
S41kJObQ0QjPnWtUp2aQHnS1IYHmS4VrQ5SPKPbqvVU30GKC3SHDAYBgVp5NLT1syigBKOSz4zka
/ohLopRHLfjwrIvs1WH4pgJCasENV3Xlg2ZmMqjFcEPtzY6rz7lXXLebRybKokcbOOt253nQaTiD
7XqsQTvSliJPKHBW3SIJPg16ho4pMw9bpjQTByapyi3BuuNovGDevP6AifMsdnNpO05MET4BFKr1
vXJgrvHk4ZEYtUpQh/+iYrffHmHhatp359ph8eMDVghLvYn2lsI7rTlonguq/6yzkdi7MJDbhCMr
S1Hx5vAPtR5hSMQTDB5MNEBuaJOA/5nXKyjJkqsOr8U/ciT56GEz9qspWx8W/FnMSy2HMBJH5KdE
AcJJBuHOiuzJss0Xg4kGQuGn9aOTqAOgXnbH1g1T4HwHlvx9ehw1qF6bybk4Ei4Y3WwA3+XMyBAo
0xzkQcnWxobompJHojYour3wUJ11HM9f4EcUX3dxogyJM/y11ffTrhOgn/3H27GS3U9wxdL/GZrW
iEOgsc+bxjkQ0XbCze7HK/qUgzkiR+XIEshajkDOvq47OgTSvl5JEQjLUKlmi+okAbDN5975NVK5
NkWjJk9KIf+Mmrle4SUSeLVPv+MrtNBTv+54DdYJ3B4epXumXAFkOTYsM0RkX0qMxxmCwIc55E/e
KpiuKmzFK75Wwlq/qRlkRt+bEf0aqqS2HPsTTUb55E877syWJXwfz3CqeE9yM6iLfdkcve/CQb/O
aV+Jwy1Rwc2VNnse+rcG2Ke+0w8TratqGZCsSd/eyJUHHweTvy74BnpsN0CdrYIFhci2mcibA3GD
MwnZ1VK+imekWNweIf7V2TInwWhSnOY5/x2K3PcFJF2c6GPmVnjDyeE7KJjnCaU1e6TEsKBniRnl
RGrXTOPp/ghNdByL/Ct731/EaChJza2/KNZOkPKr0Bsfm5lSovLBQSQVmgrp3Mr3bIgrENhaaDc2
K2sdYbwiMgqxSuIyxqPwIynz/liLRitQ6aitv+fjt8UZU6E35LuoT7cSnYd17UtmEZV5dA7E9IXz
fMUQZMlG4JEIfBZgt1e586RjcrGDCyPVP9xRSuNGlaTuMGpzJ1VCh/aWbuinRuHudXegS7MvR+/o
gGsyU87gdvChVO7NIXB9fj8X2qPoRHJYiSOTpDtNZ7dE5JQxA2iMr5AlxmeTtXGbPAdqJu/VqYO0
ZwByH+hkJ2jve+FSO67qLz4ykCE+Z/HtTk8AeJe1eerrBCutwc2tOwcg/fchglwQMoVEabydmakJ
1e3ysxtEHDkNwC8R6tkAjB3CnPtHH1QlLO7F61sTqSStAwAZVcheyO7hV1tm2hKwDvH40Z96/n5g
kBlLd2+vaPMQi6xF1f8sDBB0u4EhdFyUOHwuf8hZL8z3OVCkB7Wf6JoVmhCWFug7s6eSWjwbyE3n
KDlWo8L/oRCQR2sZPno156VH50ZcqI0j5czJDgm3RE56TqFlikCxodhMErI/nKoZbidRowGlZRzQ
ylIXFzVRB4R+nt5g1sFKAm96aDVuDnXIj9IgAfI68rEjAxqe2e48lh4dgcgbhZZS1Jki5DagC2vE
M7BEmE9DF2vUKWIeU8webAS1B9vS/r8eJC0PqvNJYlkBsN7ge6TQTYm+kIQwEn6pCFzBJf16TmK/
PdemikBva44yy62L9vdjCXWBo1maeju6SSAvFxJE8tLWM1Wa1UVdMaqlf8q2FwEfRG/kfkUq1eFX
jSZVMIj/rjq/ge/hNzppK2H+3zCy2/JfpMMOqvrAwil0bAj+LRduXTAj0T3zYVIXafQIHfH56F/r
hPCMfDELNzQumTfcpvBAw5I8Om5ivOmVo3Zb23fP1A/HHmA9eCIafYx+1AlHOXBHVWBVSKjir4Fn
FDH+RrGDNNoxp9rh45136MxLCxtM1bne/7r5CsfnCN4sKRIyBdpz0Aj90O2s61czTeh+NI6DvO52
mVzUy3IEGfVooARcDfdW8FiPACFvmtwKO0uJI1Mm4wPNWcB72Qc5S+nwEfi5BakFBBpYKrNKSHj8
2r+sJH5IIr9KSsV341MownUNmdIK3zFd6BUYBB3YbOJ2Z2y/Xg4OnsmBsMmTe9P+mW8wLsMB5EBo
8MT+NIj366aiBmLTSdMkiadC6ZBmMlPjsIIBbZMzf88ovsE5FyGQ2NfewldPrU41tcaT2asqybcH
mb9t1798d1VwyrziYORubMdqqPoUTYSbBLhoi6Dnliyj+4iP/FhT4cZ+MbmAWlYLFMEizgAiMvx9
ZYCSg1KozQzdGVLr8bRUH3jhukkd9qA1MmpnT1uwvC+oQeHgz+Tagt6I8LFB+hqF8ru93cSutknt
5cMJuKnhOUWf1K0FCY+tmpbP4mAs/pZxby0N1f5iW0qrmzYLzCfj6+RMmRKSM+b49a/Vj9kjeASR
x3NNyRGL20JCQZOK7uL0z6lkHtgG7dtk2/S6aWiV/147qbpGRF+EXGwwD2MVRm0M40biTfrB58x5
n3YvePBLYDO64lJIkMPFqcDFYMPPa12XyqW0YppM2qT1rwv9GzQnjBRZhxZmyDrvfeNGRg3GgCKg
aJau+WTv5vhP0M+0WyxxOVsNeg1pC5mvF4sLPn28IgAAsIE1XmnKD0nZyHwUS/FQdxCkP4FLH5Gh
P1EkJ1EZ0VD4/wGR678l/hPNaSKPlCpLQzA7XkEcU/cHiKdeLcglDIkNvGyybSTnBXD//XlsYmfP
Upu7gOa5aKRRTfEacSEDI0zRFEDW122IMmRQe0iybwIl6l/HjRj/BXGf6MBdUBPiGKhj1GVVQPFq
BduSx/+0BZjTq+GViOmbgpxJZ18KJwIe1f/iRDBzDFJ2V8hGzHdQJuWhsGpdPvwbcZQCiraNjNjs
dIdLnWX0J24Tyvel0Y8/hSbzmBrJUdzUrQE8q+xQaqEWrEsJNnhcQPPtDOgSjqtOsfzwox5ilfRB
xh+JHqKuKAzguAwMwlHZ3ACuOKwrHJjaw2Kh9NLix35al45uA38Snso+0vuVPfPz07NMqrnCiVA3
Fc2o2+btJhxVHuB5Ak8DikLSTP6wBbkSfi/h2mqn5/py6gnsnrxQA5oilZEbmX0p0j+0S/1IbEjD
Z3CuvB8nX+GSqddxOn9c3QKue7c14E2imRMHdotFTZFlwJZYyX0cmKVu/GF1v97CHf/j0WiYQvw/
2CQ5YIcWncsZPIVtNYrHsedEvkFSj5WIhS9a2KEkejRmtrj+Omf3tvTZ5Cu/yGsQUy3irId0vUbG
KeNWJ8q9GBBMNI8DyhHMnlN7zxCu8J11P9gBl9GWumnSFJzSL5GfyJN/HrVG5J+xCKLGM6V2ZfB8
zRjT8PDDNT4M7oXOAYU3Y6UMfIAkk+vMA3XTOxelTzvgUDMNrLF9zS7ao9ZrWNS6wvUf8bA5mrHh
n+TNpLuhgkwohIfV3JccLt0VcN2ybS4K/DsvAD/FaO89Q3B7ULsZfhNGgYLx7Lc7Af5N3OLmd36A
pf/XzmEJdxVmrJNabA351w7En4ONM93sp8jBnenC/XPZunLRmxFGvWKovD/r3wrLR6tjZOvkFfi9
BOmCmY6O77IDKGcW+ShKAQMLXA/xNxQ7MIr+wL/NXPtgQ2kJuld4sGVkZ8IlGxefsnMFFT7Mehuy
30APNQfmGLi5U59aCUNyrRDFdVw/mV/6wBD6a5kMlnVtpBwKRN1DkPk9hD1Naws0x2yNxrotjrfZ
5350mDntDIonrp8mAScw9aIAR72eJ/n+6asLaDHiaLlaSzXLAVAtNBmv/8i7U8N47fbH8PqyekfO
VOAc0yJyleqFChqinY/tQr5aj9tseDdAn1Ou7ekiHXo4XWLt73i5qfdQVIkFOgGICZEI1PsIlD8S
z4X1bF4TJq57usktz2GvGTDlAyQlNkI3MpJzBO6rVxanjACFP6bOsnaDmEQA3EMd04aZ4y0UCiT9
TNIOgn1SfWov0LWzdxnq5xcXr562vTVgxb1aSZBRpHSwcznHDt2LZhMHngOObWVuoNtK7pa/WJM3
OIAdOi+qcsp7CaM1sYYhR+0mzcbdbgJeAid7r6kUNFZfcfipZ1vAYd4le49Bqrrc8VFWcdOzPbPR
lUOUwZw2aJVDD+eJ6915L7Id6+yAGmYVx0pjaDrx2yQtCRJAzwo76+YgqVnjR8r1hZi8gvgfOT9x
sP9HP2304ZhSLgrzDVNnKoR351u69F28dOMsDkGavsOlNfnRbgS6R2yoqZCQK1fwAi5aolklmn0C
a0sVAJ3z1lsodYmILqSMdfRAMSnJd8/0e3lChsjwdDeMFsTS4Bm68kXBICygRo243zMxcgmjiH4v
ewijlyFIFrjPEVDYpquuleZ33rg7vOILHyFFEes77OmWpiwxcVIIPC/a+8ZPKgncUz4rsi0dR65G
Ghn/2IoJLxgS3xwfjJsCr/NMLEt+X3mx/TDX3TWksXYGEXnuwKrQ1zZpN+AHKyIpUoWArWuA4wPA
CPhfLnrRLgHz5mzrZSz6+Km2/dd3gWNhUJHtYHYONWpI6lHnMuIDe86hF8Zo/ELAnIWK4askfkwE
QlRYr1SNwNcUJSygJNJCBPL7E5StDl4s/E1yADABJLGzNmHMOYqa1ZEwPq5RdHOVo55ectmZGgKF
ZC9+T9c8DgqOjlcLrCe7dL0JormULToVp5/qNt4KZQ2mX1EGbAWQyHDKi3MLLxKKuvZPkn+6ecxD
O9589hOIwJZwHwDg27zDCoZiUUJ1HtspiixpQMMUcEKkb74wF4Zb0S1YH0TG7fBOLdLXukchapCz
gSJTxENW2PPdvRoqfVEZm9w5SlkJF7AGF0QwoJwbSQ7M/rMH/URK3NRDMuZsnOriAHdPlzGenu3y
mh4y/QtXM+3asS531fQuC3dkSqnogf+sILQCRhTmVH9qwvrUBBOoALbT53x7J24egecNwrnBowpk
EOfSx1bK6ZESpxvQ7CcsjXPkSRgcD3Sr6v7XfvcWLtcSKYCnS3+x+QffIKnNvnfepi5Sqtf5p/G5
3hTtDOA+BC0UCqtiYG0ui+/kKGunZ1wa/inmEidw4WSox/zOArBDBqKVhK11/3yAMLtfytdFBEGJ
5EBUw1Igft9eFpwXX7kY1aYhY4QrJRsxRHouCb9BLtMSKNODtFn9m46+I3ZCd3MdgK13DqJApAH0
oxB2EvAyFdfIt/EeL6hVX5d4hCX5sVQKI9PbMNcN7mBYMvBAQ+HWPVyMiYvUxZ/J2y3JBwQWOFUC
o1hyiTSZKf4qL5IlYB8uSX7T3D6Ovix4WTkwqMfHsDgcYr+OdhuSH7KJI2OX5N69U2Gnl0KH6VXL
aIILCAYr8LkCaLodOF55bwH4Vq3W0SsxKTw2S6BFalWvo5wys+9547ChYecgvwLBIo4SyiKz0MEA
8r4Fxd9yVzz6L8QOcrw4njBoJFMZcu2pFuAWosTZ5ucRxRNAc7GopSjtNKgri+ocAFZ8WG9YJdsR
6f22vSfVGmD+pFvrThZ7kwQxj9EcrI60MINj47Wc1ER/pBUiH/lY5zCLbo0ga1HfpmBjO92yRjY3
pdRSkNzYVbUAsyru9u9Ys/q9fahxpWMMvZ+4gR371KYhUj3/JO2/RcBYEd3xqn0Y0OJg8Rp/A368
Mhgq3PrpC5igilBbsSs+Ly/ymX+ZmO+60UDaKq5eNwaUucIblGwpDshhk1eoz46+ycZhS76h0256
4VBLSCYPrOTBlhqiYns1rHW/+teinoxHjKGkkyDV9/ixjNVyWUJLPD+jjP/+YC+sVkopkxQ12gAU
54i8B7TVcxoOZrQ3Xcr0nGvx+Mpp9bt09lWjqVb6788jvCKwfij1XSOUw5uOgWYZLdhCOrDdzhI3
cL5Pa/yuaFg/7aWQMQsqUYh9QJtjsyc83ulKxI6lz2rjPdWqCzw46nK3DCncRLR1neW/7G4mYl6y
fJ1aHMZ7cNJ2Ms1uIXMOjCJ9032RgOzcc81+WLjC9Qph5hmF5kWIPhbOGwvCdRui0W4/zSfCQrFr
bQs0412qlMqV4fR4SiYh8CEsh53U33EtRgh3Ka3BGnT70/FMfpfA00go6kLyY0E7XsuO3pqK0e5s
1HEK5X6H1Mc/bmyIgAqAksN4hjdWXCNnkh/0sSjsS+fhsIDUFbGylz9w7OmA7W9NiF+a31ohDhQF
UllcsXnT6WRugRjtRrgSwYN8JTzw6uxRmwVzoXl0YoLrE7irw2YzaE37egs/IST/ToRcj9ChOAzz
gM+ZlyIxm8YWeZ0Lbj2zsGXYnWdKnLsNRUa7Zw29Or5VN8NPiscvShBCEIBAY7hu9KUsyaQ5Aj+N
mShVd9XO0H1ME2okarS3HGUnMgecMkJ7dHvcvYyy4T1s31PVlwpppq5Qz1BFrpkkkA0NRGrWF9c3
H9uyNKP2EQOPKWgPG2+rczQ2KGsbRcK26bTRcckEjblrylye3aj1RwRCJaaoM0TEk9sTRoCPdmL5
Iq+BBNf5+suHQaiS4aTTjDEaSl/HHoyLkSWkiSDFO+8T1uF7AukeTsHQd71AixbbPEmVlAAuYSrC
n5ee5ao1hXLcyTxYFUOFL2luRt1YWv4/086GR1cDr77ys4iZMIdVVq4Mjkp5NWG+uD5fLFpllTl6
x6CSZ5eN67Uhs8up1ifa01/snrldlb5Lq4Yj+PrUGG+pnpAXoeIJ+nJs6ZG5b36ydpItBcfuEz7y
8G6syfEta46qxUdDMsiG5JuCs4mERI7+Rm0GWVd2QooJhfgYeoAcqTKrxCNe9zTFYlpNNZ8hclfm
Pn5OApvIJw87I8wWrVebA4cRat2FH5JFnYhkUeYSMsnLQgEyqyDfw+1i9FjY5N1VV8Sbf+yi41uz
JwJdJDWL5IzoW7akE5UOtt4Qxhw+8b+2uRqWuV8kNKf8/6drHR/lNCebNgKYfDZDlvSvS4ZaNGU2
mYE+M67T7qXqS+adxWoVTZy9wMsoxViKp2lfsUGBqxHuVZr2Oif5FnEWU/QDWkwscxTWjXygB9Ak
MyENnv8yvrTU6eBp87uC0y9jzRgSUbyZqa3AFDsnC/Frr4CVndd5jnHgw3v6N8N9p8lvYexPwmxB
BZDjpxxUIJGsmriMXShY5S8ik43R0uHss1XyMgclhfvlAlCnTrgE2iW4sUROw7JowyS1PXgMlUeU
WlfPltizpT08L6/MoioHQhYd74ILUMpxFNm0zSsILj/zSauAFJ04tEZZ+iDLUZB+tU63z5zUsoB6
8xWfaWTOBzJgGvBbexO9ybtBnT3j/Kr9YffrrWC1J+6/eYy4FSfew9uuJLCJVqfecjf2tF2MH1vY
rDEeU1dYjd2JVlKTI+jV/bxapjHKut7u64MJc5p58E6lGF1QUIsK5qnKzxwQfMcZCErKgI1pnZB4
M3UkEamPsLTPu00SrqIwgvOE8mGw4WBRpr2QYpYzcObC1o9mCsaVU0FKWjHosIAXfMZV+b4OLVRP
WE9chmk9OOp8v5cN6tzfvXXNKtmfSy5+sFztBjUUUB6G1qfzVzONIyPx/y001p+u4533XcrE0Sfs
3nocAscFKFGPzQlcb9fZcmLB3lTPz/8iY23i9d6j69Vq6Q1SEPr88H5hoP7Yeim8S0pwJEuL1USG
uRvSaIUf+4009W8EE9jzq1ZZAPhpboz0nIirRzaa92BQwAt9/7BOwX1EZCjhFHKNy2LdrH3a8xwm
z2JwfBaiE3Ypsvusrilj37s8dv71y0e2wzhhE2BpfyD0k55MEPRaZXdv3hRH+HfQjDHjP11MHmys
4tThPrIphAxrZOhPxi4RusLbQi1hOMipjOi1jGd5rjN5+HQjCeOGAQAqVzn5muQhicf87qwNvg2U
iSeF1drsC8DFJ//RnXK3C2/mQt5Ut8okmHs/Q8qpV/+ekER3ZbaF+GoywBzJrWYQtWU7gtjSJ+x1
S0ziX7VEYx+JZ/qbHPGaNP9IaPiUWaYzpuh+HX5Io8OggVdjHWzP86JGCdaEyMmCRRDshmeyGRBx
wSp8KEFIYo1LEV5BKzYFuDCSM6svD1fcETKAEdNktuKittQi7mhjz0RvuoYS1vN6tnBqVBSrtkjj
cwIRn1csoUVvr38OSSjw508qnaU1Gs6/ia3SNGFp4QQvS5Fqkbq6nsGPDTTOF82/xvcgJivlqSQF
ET4iZtUdx5RiWbLOTzZR6I2lGF+f37DDtRJqGbHs0quGQN4XEI3EYGBc3q98wrvxVgR3Gw/tgjfK
UD/qt/rmANKYtEp2MFONNX5POWkYC/da2z9+Cgs0ZRpdc3ef9GvfcEJa3L78kpwKFgKcyXxTyhP5
C+maGEjfQtH1qpqiNvERPXZ0haqf2wczg6CwsB1O1NXgrSug70aoAWIJHe6mtSLjxWMnqA5z8/jn
pokoK4cxcceNjKqbPp2oFKlM8XFMpG5UkHoVrNls65OuSfUA9r1uFZqQ6Yk/CayjSfsSrJOi/TwB
lnCqB7hblB4NvTWIQrS1nwjWXzSe1Bcvuy4odla1BnXqx6QgRHI/HwUrY04xhtKJ18idhBmSoGUN
DkYW/uEWGdU42jhb7BLHnCx5dBwV9Q4Bc2NWMf6q34oDBdA93pM9VgD99LnxueMDr7BBDZvM0+1Q
Ou6OKllvrjM5Rh752mdPmrRDZ2eTBwVPVpVA9X7nT/+HSTTFbV125t/tQgAibtX7q1kroWaoDIHa
nMIONEJKs5uluC+667/BqkjXoeaLShPL5TZWHHEddKq4LgQh2arkpGF97EMtWF7l9mLItCkoWlYM
RDa0mpXxM0IioeVhi3m/0ikT+SBklMgXqCfai2l+bgzMNrNASEiEDG/TcJpMHUENbR7B0BbUL7/l
62ZSymJttvOs7Uot7GIPhMB/Vda4n84wS1JMMREzlly0tRo3RnD05QPWyhouWxxylM5Uq/7hkvYa
vOxWCTzyUvTQ9BI99VH1Em9uC/SjUDP1Ol/b7ePcjGDKTJZoC5mTRAxXUHYRnNnCaHBWows5oHsk
5c1KkRlOZXR7cNihid3+BtMiGS7U+F/Tk6R0I52rXEWDM9V5SlHJZBw9mvudIZvH4OcWtCCutkrX
c73xL3m3IQ2yFFxhI/YCsFMmCNv06vQFBbfTHfEVuKhdF9dUqS94xh7TXITBfUufTXmJQMbPMHcs
hIBRyRThin3OJJ5gpnO1pyz2KInqBcQlVpP6RVfE7ADDD5HR1ZBEKVrbAQ9UM0bJuEPlBt2QERMb
E3sBmXOogGKCEFGH+stx+Rn6q2vyUnKHqEVbnEFvqPxbrBIvvufXuYbIJB1MEIy5CKprgaCNNdNT
bbV4Axh3NoIP6y6xUVzrzrByX0E32aBNAd2tlc8BJ2ZFCMOvJ8cMtAUgrsSe0k46ehhT084h0X7J
v2qGJw8m+ycQEAgOvEVuIUeRksIhWDGVBL7oNtSxF8nRQOvjsUJpD/p+YuhV44bsIaBKssiHuhu5
pGJd/UOl54Hcvjy9g0dq8328beColutZB6RQTwILhiCMhwfKEa45ap9jJQ06gQe/OkiOSkgqOk9p
26hHVvdbTEkRAApIA9T9gpxhJTZKTHXBPDAiY5JwbhmGVg/N5P3Aczue+hcaq490Gr1mwlpctXJg
fHM5PrHrMV4oCHAWEiFpT4D2jCLqOsQoHBA1fGnhWw9Xtbu1FXXMXXm/d+swShIgwRA0dL2E/T8K
Wq0JZwUffYiwq1aeW+CFOkbOcJ/P9l2153b01AQ1+gTXXjHMk8jymsTl9aq74Q7dmezM/LfJ+BtM
ttmDyhngNN4Zs3dZZg35Jfyr8nGGBagJBsPYokQI4dHUYm5fgCC0C59/LsOWn8YS940fvLlOkCF6
2Il8qvBgvJAEq3ml6pOCki0WEyKvVO3t0DDqpvxBoJfqYY7laYsgqBDHI2zC/j2RhovLxzDhOAaM
TfgCcCcPpLJ3lnYpVUsypsWxvL2dYwDwUAEXnZmfHn1uX6+8GIGfFTTPrP+0uyBcY09wZiC9+D0G
HB8gEhFe7JnVQIb27ThsNXCsJlujSD9GOFW7FVHGKN/fMnCkUBzsFk4ElKpgkYlIBNdLyzA/wjP4
lhuYZMmOZuv8F6KKbuqPWc/ev/P5y/peiP0sxfFJQRYtUaFFMWWx2Ie+9U2puxeJ8NPwAmkvAt2y
PxGT6y4ZNgZHygXbwwwe16dvciCv0c6PiTv1OqISEGvO0KG8a6FeT45S4MgNSerp8jD3bq2G+ZRw
g8j1Ju+jctBKSnCzAF2InFyRuAXuCUkmGqz1v0f3294qvDO0y5m/DUdKoTZaq/8v/JtvtepSMZVD
ewv+6sF2HXucVn9omN/9ASPVgrqnGz1Y1pVu9D/Xg1HrOzpLFj9hZvzlbguh/h26Ra27XzA3q1Nu
0ZTovtJgd/eXBteoVoYL5Mzx+6ZRDUwFX1yGDX6TkTRHktteCLqSk1CRs4UHUnNXD80O9rNszlkt
aaQVjAJtryxV9Vl+dr7umGQwrnhU1c9+2M6Px4EI5/Hwow3VtgDw5/cLzG0AWbKi2GQGkaieWi1O
CoJJ1jUrtegwEeXtLwW6/qzugXWn64gyZwum/UL54ulvAeMOjre+nebHVG62kXQ5VOBxy6OoGH4N
IeenmhCI8K6VbVMAlv9EA0msPVB97i+dU3zt/x/hCn/2WCtOMrZf13WTbqvvLYKR/VGDwjg6Rr/F
5LJNLjDWVv/CfMp4f+Fp6uVo5RKTspOs4a/QcrsGdlegF+VngNSrLsSkOlukeeUTna+WoXcVG4rK
m0E6ccTQESIzNO/tSlZlvKdfAOsF5ELDH5RtZoCRXpxnngDWF4+iDosUVmLzsSwIfNU7rqgFSvpL
rC4tgrk06BMLerWnBb+FFIhw3HAPm4boUq5MjGBDnXq4B+NlJ3mMWjlFImlBtIyx0acXous3U5JN
kw+gpsrzo1SczSbxbUkXZXex90wPFCu79pb3EXClrGNYc97J4mjLJMkGkDptWDkYzYb080Ta01aL
/oxrWWExICs4ZOw5FL4AXyKJcn566zKXWEw1iltMy1uLlCMBZBH1GbZ1GcM3JtuuWEOXAf69oFqX
UAq/Gs9t0OPeDil1lGnGIs5zUMCJcMiKizFHmOaITgy7DHZ2Tr7hha9fZY7LtF8ob+flA10NDaCv
ucTEpp/HhaxAaVwBus66DlpDCheiMge3pb73NnTNYhgeP793UzpfFxlbEWvl++tw2zkQCF1u+Zar
rwPV0SXM3saW4W4xDk88wLb1fYQIMNbN/sdBJVHXnEMIF3/5xE/3vL9bzfPmpe0m97LMC7RlDxRT
/jLT25BSavCIHqhsgVH1QYn5bM1V33+FBucC8a+XJGYeLPPltY1zWUH2G9u0NRMqz64jRl4p2fab
n0r2m2aoTVl6pqL/XO60KGTNioBbQGw/wk+ivmsY+fORnDSYNSyptFUvjsmCxNsxCPeFduD8FiZs
cvDMuzUawuxB9ZhCwQCLDtcvkCdUWQqE/lSr5j+UipiRB/oJhw7SdmtaPLPfqTeEiNY3QijQQfgq
gcAfcGRigRJImzrz1EpD3J0B0lXb2c97CmRd1ZhqrZ637ipyngkzpZ8SoiXzbUGP5eamedW+ubHl
eJsFT2Ptr/8HsD23XbTfhGvEaiHLOXvBWPjilZK1HvqmGlS/kdtENmNbNeD84JybUTRhr2nuyKlD
I916c1g4CDybKtpxHaHLLV9HNPc/YSQ1a7VpbQHqEDilqCO11DeFhIxDeWaFVhia2kmd/j8J8O5n
nyMDCBYmtMHbXUfJE5oxqS0Gtcn1vM37p7M/vft1C7+r8zgNW8ZOp1iva/ctcNk8Y5dvGxaO6hdU
JZ2MKXBK0Xa6AXmu3hQuB6lI1FxP/ZL1spe6U/1Oo1wJnKWyj5Oq2qcM/IR8d9U4yEghYAQy2XAc
QzG1/tvfFBdWAQ8U9R/N0+zYmvv7OkYHU4lMuQXv1ysIEpB4BhSiezMe2fdtOv804VUxZ+tHJo/U
pE9dJr+IC+zCqOQsniBO0BHAue3qu4/m01lXgC+n/vKZcSwz8Wi30dVR3vMohspcuZ29inKY1Xuj
QainP7UehnYIwx0X7wkWAQdbyyh4ZbBgF7A0J1g2CLPDZ3FZpP7unBQ+YNo+t4O8L5PBR++14BDO
5kH9Aybd1aVml3MHz//o7bCu7H/qsR9dsqSVDvs6FXL7T8Rmi1uZznAOcveBtr3/LFQhbEDF3qP6
Ees/k93qvdq1HKdYAyN/d+rIEbS/szO5l5tI33IiRtBNZsB/RPNv5X0LCMcnOD7aLw3vSvAL5LTc
pRaWuafFveGLHqggHjmRMADNwnpKI9JiDzFUsKCIWdRz0B4K51hxhDHn9uWJVy6Qxwtq0t/K8eev
6danoFvltxI/pSZsBx98MKSsMCWhZflrryx55cUkL4U61rTaINeCOsN4RRF6h3EpXPxmiZwbFjaf
ylH8gl2n+RL/CEGZXwiXfzm1U38AC3gQabHkEdQkj3TYntB2rONIyc9V6ZqbdUATmJKMGDF6T2Rk
nDp+jhDVrLqYyIayQeVDic3vdVu8CQjqC8IxyW5EkBitDtuizi0Oex+EsoHeww2nnD9oX090Vxyv
klv4thK+CvWZWRNR1WIV2DSg+oz4Aencseyk1jZXTY2lJk5WLfpVp9McCUf+Y6vpQL0QIthaoL/C
z6NUJyK1U5V8x3oJe8qK0z6ZiQ69H1tON+LwA9pphmTqsxPAZXEesMlqdyOIr+csVGsgNtQdxsos
6tTJpqtnRIllN/H0YvCgiZQJ8luJjl0JaGEVInZill/EYZFt7iHKAYcN8/uwqa6Vilf92l7INDtH
m/Bwzb0HR3SfVLQ0e5JoXKrBWJM0sqrwVQ4R+2fPvrL+Tw4rGHojKRsFhvSliwvWWLcivbj4P2tk
sbDQ+C5ro1XChYlNshzN7Hny/bxwEhN/c5E5NgKk9dfAyH6I86aKty5p4IBnxfaqNOHdjuc+dtbn
0K2W1oh1qFS2PU3N63rtMYvhJiLk/xtfzOaCKC9q2BSvyfDl/09ZnsR/n7avbpG0WfL2sAhJ2IGt
6cBq6P04grQJY1N49+obaFb5N8laQyvn39BvvLSEkWWgbVnwoEswv0M9LaLifpuGSHibtc+dWv7E
yvOLDnaEvPvxYKKglijG24cXQpxnXDwczP8DmR9lNqu97dilpzRY/G5e/y3aXPPm3un5W7XY8gxB
WprHHRwLPJ6G/Lp8lHVLo6v9UVsLVOHjIqUAgdI3vT5y5eN36ptb7XizxMxQFkfjGqw22xR4RYm9
EsmHf7MN7YFDIr25O1UOczYvzobUvaRAZn0N17vYfG8Al7MS2gSUmzcvSfxFv2/ugCS5AxQ/IR7q
RXzAVcNG69mdWcalmOyBTjqHAwygZAbO0cdf+XwoYS3Dhm/6Iyuq6UTBiiPOE8DYpIOiD34XfXLk
dka7dqGLe/xRMy5WvwAYxRr2ewJL1j1oWi7D7GTA3tk6pYODb3w9+xVG6Z6vpecZ8TymO2nQW419
0bjIe2heuZkSAIq5SC1QriOvPMir6uh9Tj7sDZR8mIMie3ULOjD81v2Hd3geqYw9KDi8iDT+b/Sz
7Ku0yUUpcI5tEw3AUO5QzpMn8VUE1FDAD2GGgH9O7SgK0n8gO2gByg6mS18Nt7VDF1NnuGl5XBho
azBAk2vyqjyxeWqTtFW4l5vFnJm5j4atCHIVd55v9G0mC+Yf5KRMFC+oxTRlqN7T/HEsP5xqnxER
LGSQgTgnzQpHI6JYxcAWgGXMOOXo/KRkvNe3YycEZ2ozM4mjBGeA3fKmWjw9BtOBSq6yqihnI3Mu
p7bFvsO2PgYPqxa3GPB4ax3MvQpG2xJ2fkcuru/tqfNaY9tzFQp+r7iPH7lH5m7SyGg7CNeBcCRb
dxJjKwwUEcJEM3NZNM5N474go/SadpXZplLiMnuPKE70wOO5hpXvg601neuRw8QZORdStK/B+Sbi
qUwCwwE2IlkWetDT6fPssTGGqACNw7qKCZOOOTU4M+NF+Jv1LgCjVEWRI34Bq05vR46x9mvQxVa4
2R5um98jYrO21yQ5UdWOXc8RV7iaj7tpIeNiHoYKy02LrGDqzah8Nf+EdaLw6KVNBZ5pmW065IbU
2fHaJFDLhN9+Yf0YpNAybYiSeHWnQtNfaqkkHf/yTftsSorNQzDoquPezDnyE5vHhkxiVsKbTUOd
3wl0NxFq1HkE4iBpntiL5YnVVkA0t7SUbV8G6ACQvZuTasvy9cyuqH34zp1SNwqeJlxPwwiyr96m
TAyHvnk4hkKn/yTlmxmrtp07h3ApcZ/FICcDcTwSjJ46qKTMHUlblkbpESaLcToiAvZ1JB7g/63z
DyNolHOrasSEaaXH5Uc8OuCum6R9JS4abNhj621wmIbRjPlkvBZ3z5ULd0jhIc7xKlB9uBTZI174
U+4zePyXSHHYsXXPl81vOozSHldmdEv0LV3rxl06fvoArhW+Fvseg7ccwbrNwwVLPj210GU/hUyd
K0fBBtSF9iqCmeUzPiMKwL4Qtv5+mOJCTgUamW+fsxl2xhov/uaesCIbaMW6sGROecYhkQwR71nr
OaFeaCYCTZlzbzGNeu9NLz9xf+QDQmKkx38aERIOAxMeyTr31ZCeFKMuimtpZNL+eXnwZPGPrP65
yDZIXt4jPK95Xm4kXtXRmuMlgLB60uvZXy1VoqNP8FsqHoPFCC3ASdyVb3TGkG3+++h8wjE7wplQ
/UC1kkHY5GwRKFrVO5zgJ2/T15g5PriIb0Z7lpPGdaujbca0ZBRzVxp71gQZGqMFepPF2eDd7Wmi
MWUDCBifhK+FS6/KnztZlEW1O12u42Yjps7x9DHnWvbjHOykqNCGpqvi92FOxIlok9nt2dTqg1Xw
ki7Rhj3ZIxSpXzeBo/V6hznCTQ9lvg27bDtjSW9+gHqlyo6q4+pc0U301NNkFCVqKkOvBdpsPiKu
NYO67MfTSJrzo+elBxt6VCqhNEA92hepBFBkMpeJhEQGzehhDS8V225d71hXFS0A5q5uqYml83mw
ACiNTz0xAOLn5Br9jVV7FWZRhNYtgyyvmNR2mONBhIMkOb43uZZyyXu8Ljxxek4/g+7l8iZn065+
cmIHaAKpg69w56KWB1KYXQ7D9dN3+gxFkDO3btRDYOsZ4YNH1Y7p2JtSTzOxVS3sOKF7kS980K40
LLnMHfciTrKNiZFTfnU78OFXGDnGYet0jdyllQ8O+ohkXw8Yx4navmS3UEuZRCknsnB9G9LFfzBn
PYFeJP0FelES4Z+nj6TDKE0/N38mjXES+3cFM8hp/lrJK3q/DrHT86QLdGdHyN2OgZGIszk+t4ms
3eM0Uj0Ze028t1sIh1LirpTlmHf1EeFR2DTSdgDS+pBK78IIaIptiVUjv1yFnm7BPFDdAa3koMqm
0iTk/b645NPBs4sGh9tblISAgTEKdDMboEoJPfInO5tpt/yZM/vDUQyWnnv0vCdsejXs/QS1i15G
oB+fPNvxRqGoT2ydztmdt2u0fm16EcJ65INhGkQK6DLa6IDKb8aggqrYSgo8cG4RYyJj5EA5rVaM
LsqpfTq8ovDLNPBiN+PEcqQfrNITm+UytMddObDQq8daybuiYrUhc8WL4zQC0pwd9chMvL431WnE
87DTIkR/MYupxTwxFBDpETs8nxgR6s9ngqhDogMbfmEi01ldWrO1+lkOK0kbsxhkKMZZ+PLC1N19
XYPaKGQih9T4MALk2nPNWk+gqZ9VU0twWMmpZrgUBm5WJ+tZCOFM8wBzmzJ3DYHZeGUCnRT1fb84
GTkF6y/yR8Vhp0FGuiDVpuYCXvHpMorLqYA3Yej1K5rCPUSv6p1VmHLywAQvrLWjPjhx5I1SShfD
kHjVjBK0k82kIzr71xj0eR5iSp9roJemD+cxOoVuoaIHmm1yW9llHduX7QhZstpvsCHOOf2jTr+f
W4RY2aBxtGwJ4DgUmBTTTKcEvNEycMblNNoGVQHExRUukU1ee+JOj4O/iUPXiF173ppUbLiJ81+j
I63Lcw5UMPA7oKD7I3hItw6zs8WytYcvkcXym+9VVP+NDV5Q/sS6fTFecgH4H24+30AffiQQHSpk
OBXm26NH7BYDMz84KljHbDInaGS1/HQZsUIvQHSAsZRbVLIvVLts1X1GTOaFMZfQ5D+fKnlbeAVV
vIf8Js3fzhT2K5LYDrDPj2ggRTNMQHSM6+kn3jsRPFMqgy1BG1pQFZxjT1zrfWpcyKX0Egv8NK7V
ugvFrSmQgH53/zmrcq3ZEgIWDLpIaoHNGwxIGBe+lGFGqYRhFK2FLmEwBlBjqRrlMJR5hCukkcbX
4zOWo59RUdkWl3v5yxwOkSCtc6U8XllVKx/I9SHcJf/d7cMg6nXLljS+MULP4jleP7DKcME9xms1
hX7SMYfmih493vUUyPYsQz8so9m2yaBbCpxLsZ2V+nmDI4IXS/CRwGrHSeHCQ3E7NTglr5LYJpWi
gA/x1wze/V0ghNn67ba/7hORr83hU9vi/uyFTVk8J5wJTlWlCyYp5LSDLBlb+MNnFwdCZD6LNN/6
yqfT3XphwYDliVZxQ1TaJIjXy0CQYP6cFuEal8PRfpjg2Vf7JZO984szhEZWYfnM6ScbEjWAXolA
ywo0Bom0uIsOWfsE8GUvmzFsJq05UU0m4IC/4vQnXT1TBlwXqHapLLejorXHPx520cNhroqHtmJN
8OUQu+c5EFirx6Q0nFEG5Gi6739aLzB3Qz6K7ITEs8GBW4zstJbW1fUXIwa8eVxdynUaOUT13qfg
MwSIQ6DQVl1bkZnmxcNOcJmPbHwUeGFI4mzpK40VqFZmMc4P7nknjdFCtgyRd8bJ0rUZkNGJvciC
u4VOWIPP//JjwS+baCGUQRT8iJmWxVJEflBOKxTX9bPgd12s6XjM96QWvZcHQwc/eMaUuGjHJPjb
zJAPH0hfNFYFYe0DPYfDw5YVkWuSUzTO0JO7s5S630Njhc8z+GcdkS0A3nkfCTNP0gR95bBQlUgI
OFtwTjp1680LV96ccRQa09MwdovzgUI8P3yVEtVIsDW5zQcLZ1H6qwZ2dHJzxdwbGQTUVsuGzzxZ
Iui48B4kTEYlsTh/1sLSFkvgatw56dBLoxbWUbZSz5ABMvmPByWmzZdEzUOmyyhnc3uDCyO1ys5e
zhtVhgjDj1iEUskBfIijI96Y41cAUedIKUylrqcR+Tuauyf1EdTDdWpn2hg4wL2wMNzw5nJqw+XG
ULml8rjoIERX1CCxGqXTaUAsk+osBU86fq/Kp/NmKD22l4KqW+gwHGVXUHFYbpy9Ov2tbv3ch4HG
iOXKdGdiwdp+aQQEIUka1YG9HqwJTOwBuw1DzF6RT7gVJHb53JrP2iIZ5c/NUeFk9fm8mP2PtAc5
BMt1xKk+uFlbnSlxesU4LYMk7V9VrwCd7WMX+BK/fNSYLEaXe062Du4FvD1wJ8bi2JEd+lGVWQXu
udWonNZhGWQBmlFGf5kaQxvAaD3iMIpTgPQnYRXGZrlUCnp/oK5yOWG+MSZL8pTj7qAgMmjgQ1AJ
oRZZHVdVhh5P5WOkyvD89DuqtwtijgEZTld8TmWsICiHqRc4fithzPSJXa6TiFl1JCrulTQFlyRY
SmtUE4/ijb9rApDcGQC9QrJMmpJoXNxrwYR0fqXZkbyOHedjnRuYqESTF5bWzvQgNPQ431sk3Efx
qVpAkWh0CejVfWTlXJNCyuf7EsWR8ieUk6tPCbzdN0n3QC8LSfwVWpwtMP5Qj+qXEM8H4uBHYSw9
kvMW9xKRdNsSi+CHm43O5Bhx9eAd41nWKiZrJwBzl/0vmQUSayvNa1o+oVH8f5295r/UhfjMchGi
04CsNWB1ERCGWAJ5T6LpQOl7NIkJrTiRZ/Zd7XmrBPkfKNkkIeQ+jxQiixPdet4GIPfC7PeTe2nb
2OzBgocgNQeh+OnU6/gbLbn1Wi8GGOBDcGs1YeLFlTOn6Vd4DZyZ/pKxuJVE4BiMUeia0IJAKN0N
0HSOqZeQhL3nKfzw0z0yMdBQkK+x0lmdEhI0DJpdLgXa/KWUf7Z/N4eyWK9ylXjAJDSgshycReq9
NEAA6+qnE9SnrsUETdyHa0haGRaGpNK46+GFRaruZ85MDzM66nY0I7XA/9z4/U5Dolkj/f+AQSx7
kLRi3h+qr6ID/DLpqZdDKtlzbkyKnDTmFBDYXvF+kNpRD1gokK7KQ6iZOVp1mnTZyn52FVV8Fp/U
O8KxKzlUyI8sEgB4HWdLJNL7gsB0dAxhp7mtzkQ5Mzg3DX9wJE3LMVgaxCfaL8PFar/AicBobHvn
sXEsiWDnew+Vs9INajiQ5hyS2KsjGiq37lRsNDODMfhFcXZujrUjMOK4u0bnfTem80gSGPOC2mZj
ZCpF3MtunhdB2eCXq4h8KZPliy0P+6jfY/GrFHibyi6JUVrC2pqQWGsMN/REY3fGC4UguQXDsoqN
w2hj117dFbpkQTdmhT3HM29rC6CVOh/s+I/0qzerQ22gDpYVFRzvAuWcaj5Cz6T8t2+7lPCRnJnk
XUlZscn5G7larHV3r6bbQzWqzkIScNpwNPVSmlwuB1rIFUx2IDSpHwaQJz8pP1JSzi5dmerrNVgQ
EZ8oa2rCmoxWQsVd05v18Qd2iYeFHVx+NNcltvHcqd13hyNhvXL59HPVkDxdRa4f30Zn+LOIa9nv
KKBhQVku2hRfX4oMiHOzIw1rArmhdNiMIrqS35wJLYJfqGd6z/QNNhOO9EP+UOUvakp5Pob3/QTF
evBfalp2gDkY5Fm9PPzO24e5Cj+IXp1iRxZkZ7+Sniregv3GRTl+neVRZTPQP7FKugP456Z7C3zA
cnSWDpwyRKbJ/hTOG1J2xKb1lp56MldQ+Ke5Nc1vi3YtbpNJwb0oFWdchkVd/zJuGcQhJBig9QYS
fJE/kPBtSPLCFBPkEjFk5BNKeXAGP1yixE42H83Ja2MF1AJ9G1PFa26sH7BO3Odc9sL6aGiuW56q
X+5OgeS2pkH1ZDE6XlV8fioCa6aOcOfc5R26U8n1ERQZGsWBvOp7eM6DtdnhfDVB3C99+GKf07U3
idIIJAB5ep64fLJ3PnfusWyi7hzyMeyn/J8/+MRfheFymNdsRiVTfdg/B04LoJjjENj8ydASjBJ6
RTUV9YAX/Ndh4T6JXHxnF2ge82AQYuw3n80cRp5BSUvAMUDc+Pk+qaTU4upESMqJQ1VlrB5S/tG/
qfmGxGM6qcyGIJ4twliRMhy9aYw0Hz1cFlnpa1rnlj29PNbVmRci9/QZwDMcXc/RfKf+weo9Reoq
v7l2jAL+9tT7K4g0+P28PLncUp919x0+/UHePoQ9O/Tu0dBBIJP51z6PlTfpvp74au67F/Zup76T
M85Ji/W1ui3iAEW332Fuh/JeU7v6Zix6N6z93fjfyRmNAD44g1vtsT6rAaSlOtKzGw73g/f8u5R9
YUapL/H0P7p+ZVjq4+JnfdvXNPBUzD2TwabCYGNT6/VwotOtaHxatGGozbRK9x9lSlIm9gjVwLOG
WsNTn66NO6i/2/ytpUE8W3omWwkZh2H4Ny8BoGNdbPZ7Nt8j0jF9BboLpxu/+XOhf2PgQyF5Y67P
Wa/iwYaJvg4LM+LHa7XDZvNDv/EMQd6wbi/q8sYnX2nrYBCHcRkMMVEhBvZmNF3dGY4qDKr/cFpb
eMKOzlH/i2F/6glOPK3i0kTUwjRK7ZpsY1mnF1IOxb9aFMYUHrrkfamfyVwpvAQr7aUsZJnLUrgj
eAMonMGfvXI5b3Q5mOlBsMOaHoPyusqtbNMU7wnGtBFR7RmwDofAJsd+X6Yq8maV13iTpSRXgr4g
w9Vt8ug0o2VV5R4FhX1gEclFoqLZYSEyE2xj97P3ohVmtb7VtzG0Pukbi/HMWoap6nAe4kPj6FMN
e7aANJ1pzPYP6lbi883DDmBYsK2KDWF8qsb9fywkG9LZ0wNwNh3qVyrda11jR3TP9NTyuzOom9Hx
9FsZ8e7S8VGhx9Je2hBf8A39+QrcdKSXvfSj9vCHG9x+IcK4bhz96bMvqLl87SkIer+EbqpOO2JC
EF8SbONILMc0pdeskH4A8c49oKPAJz1lC8/irpU0MDjAS3yKQTNJQId1rn4Wb3yyk/hNYA1jOv3U
uc2AW2l6gTF/zCW1nMVdreQQ1RFZte3hkFjo/UpnaSG1sJl1dICXQF9XZ8gAyYAS5Fv0oZDdfsLj
Cqgb3jQlkb4NlfcFIVQ2+9B8mq63jt1wiA+SWSOmUAgIZUTd2UPh4LUIPK0Wh05BsmSq5TryEbca
bJbbA8uLAGYA8zPQ/gUm01VD6XbgUezwrVwAd/DI3+5ok5OMgBSab3YFjZwhv1Rk/7ht93NlBuf7
PA9A7N86HekvQyBwQiCn70M0MCCFLh/JEe4rej4n6pPQULYxUJDqxBA2ER958TuQcfpFbK+3avga
XuiGFtKemHYAWSlaoHPpBCV0d2w1Q6Hed4ppmj/AO93hY5ZIJGdCpIxxqXOv0qYdQg98tasZzhrs
eAGnppSoc1ssnPe2VH2ZIQn8L8Eh7OCHTreO6WLLlEfMQm8UkWIMuo/cqEbGxUnhnlsr/dDcEdxU
1zibq5PuHkCscbglRXwaEfbjJ6e+ZG/NGp9M2y7r4cajFhbrHGPTpZTUaVW4WMdcAWgkbrpAnQqa
spmGmcOuEKclUJ2P86pSAAON2i9Hqos2d7mbzYpGXQ2FHueG/aCyPXxuOnyN8Fytx62hZ23UiZ4j
Xnsog775hd1aGgNKl+A0fg/lX2rKBwlYaU+KlXoJxx+z/mPWJXSnydkWq46njrfJi9UdPw+bkI+D
7K2wdvPloMWbR5E6qbKzAtUdZw45Z5dc2i4s0ygSg35DQ7beQmm7m5Y86uCvLAPADKz4ftHWoBmV
ajPpUansG32NGAjKivfGMKJ31Z1m+YyfYOBb/o7jt0grV87tH81PxM1dFsaMdjFcSnEKeejEZeG3
/ZjaYgJ+VNwtwqTatRDycPFuVPDkIbVTDHe4a8TW3BGH/wnLAGoukg9tTIrL1jOo+VI/lCIlwThq
M1E75fMBHFldnBNnBUfWQCZZiEYHsXXlF7dlOcdng1kj5GgdNDopjrKttAbMwPT6ZdAFA+oPvvPT
yHg7oC8XQYu6p4NJbeXxga+b24F2FQxdvGaibn8eKbCy6+7IoL7cmUX/Wo3FTDnsOOyuDkQ8qXQF
eCGtJRcX9XKL1AtS7FDuX1dWv/2uKsd8sbTsTsZOrCFgjz51Qb2uHKbRt6K7x+W52ECFM1Hjvasg
X6YAC3if8J44oJVLg9BhIzlPJteS93oECgbtyppnOmyqQ1hLJHyGgDj98ipnUONtJ7Tfm0zZUC7t
hHqRH6EeruC6Kc8OvJTWh8YPROnAgbNvGiKw/9eCaoKz7Icv6mipdFEkP/GG4pe8XISgQWT6MLwa
6s0ljtmjL0anSkon2dmgb+VJjl93s+If9EoX3fqEqRkdq48vu8iT7cNuP5fL3nVvUpuOApHxKj3a
Ck3RCK8pRnTVYXF/lmNHioKAOqD2J4rN3Hv394zA6H9ioXI9js9g3Cffl2xH+mG+AL5TaFo6Elgs
66+5XW8uXxyBTiCWf0h4YCYyzHFyyyOtGUdElyZPX5xCgcnCz438xCbNQeM3vNZfEDnLJOzILZjs
uoOhj15fvXDQ2N9enzry9jyng2mYSVeesMDPCoZQkPltA3aGxHQJdUQl3B5geQy5w0ynNFEdpVpd
L0mlgbykZ6MmxBNjLvFc73MfexX0avibSDo/bjhSQ0T1p4oI9NSSg1JPW3rI7bXc/F+IKA9qRX8A
XeggP+9xKOPC/XJp3hYTq0hYYugM4vM3NvZQ1u0zGs72xYuxAu61ExnM42zvkzRNqmllAPF3Xwib
khl6NOESO68zlDWq3dhji8Oqjpw/gMlJ2akfRK5jw6y55mvqtu5L7wPDB/U6E2f1IoAPbZ4yNscS
dR3cwnWdgZ92/ELJROQHgnd7woGbpyOKwjcwYPAr1nxf7dLDCxVmQZ8swhfMbAQLOW8Vi8I8TXXn
7SCP8A32GnF/YgcWveopqhS051oLtQGMwTG+wxQloouf4VObAEzaZ+ed1oxE5KATTDMCp6Z+37D1
fcZKJibRqJoUWY1wdv4CkTHsZNxokbcVMsGyZNuX54JqUfzshIovhzzj6mY8yoAeCKfYQa4Nq9wy
XmgP4Bx6S4fBSMVN9m5K654Bc5uSygLq2/MdU1XYcz31y3bZ/tgGXJWfj0D+SuirfEX/3SGaTGFv
5oTKmzRnZ6XyIX6fSz2hzyyshQGte9DHW5fEkaqaGkQZdU3YVIjRhzd3IMoRWi9+gIzNsNcQ/Pn1
wNSSa+Sia6RtdG2uLQp/JnZET9lVp68qxLQt1jkRh5Y5taytkDFmEN7JyfG/91n0OViLUk8y1mHs
cqT6BnV/KX5e3fo4dvhVFPxoBNDRccDQ6yRvgb74vA7VgennGqtu5wRuc96CrBUksG+iipjGHHXX
UZWRLyvj4wF7lUWRaVdira88v+iNHE8naMu7Q0ebF+LlbeZcKrN6m0Km+E+jNRmRfQST+tqB//A2
zc3mogF55jgvC8A16ONbE4YbdD7AQxysasTmY1gYnGhKI3n2vgxgam25r0jde1pFiekWehRydmS1
zB2nZDZoZtrRTu+S2hsvtn3vMzie8okUcxrimGqgbFgcdrx2K3N/Bsm0R+UeXEpSiMAzLyx9vWke
m/SPZuzU/cJKhYdrV+S2Hlf492NxgHP3E4KNpcDCND/UGohArRAS1hv/G6zxMggOFtbSLyQrTiBf
OZrGmMNgA9vs5NuZPwGNkZQJY65xtP14uYiHyuyfJzNeifxSp6tmXA4RMO0n50CUhiaZQQPAaPfb
4W43aKrBV2zse2YHYxgH6aggQ0U7i0DnMXDG7ftmyuD1XzMirLejlolCsaBXvxO3RREeX4W+PyCx
RdFpANM6b/yICw8LRUSvDSJMG1YyHGkAzcHDcTNOMT4irbBWuns8LwB1vrtsZdBgfPgStwVJ3wLU
kf0t+j0/N5eWmixD8iolmEEb7Ui/aWwxzSDaJyzEwyCb7+pcScvYPaZaf9bTNy7YJvEIkM7majg8
TXuBAcYXOBJCw4gOKgViFAaInba97lNsCxWJpmxpm3KjOAPsnwdrxBy/d+HkRZTr3Nv4ZSXzngg3
PaQPdqwB7uurLYOvPjvl9DTohSNO9b8xeo9STBGlXM2nzBCrp7mwpY2Ta6qGrkT6j2xgRKT+vwXT
TEAPuBuOK716TxNg4V9QpNTGe5qkf3N4VdSlERo7TF1n3IlDC+2A2BnAWP+LyES1MkcRltUcFP1u
dPx+v4Pv6Q46sR69v+lz+CsbKoK3F3XGzPieOkUOHJ+7tPmZNB7o0foikLuBKzHXkqxiyjvrkOtB
bAUY/rmCXWMwGwV5Pwc0JIW+/02dbZuL6WPEuGQEMQp/7OvmUy7+BwnsCK1o4m77dtt5vWUlJmml
Jv8eSGbfFlP9op+WXVD/vVHAJzPgIKwb+8tSFomJ7ZnGBV9SqJBuz5OACQokV6PX9bZ5NfMU0az4
IDJFDlA9Zz3Jxv0TiqdniQG+/+rto9XMw2ZrsRgZLY1C7JnMhLB/Gqmfvj/FjcabiAjvQmYQ43Af
iVY5Q8LPXqXw796aHypfDkSP8SOTWuQknhizTIWAgpr0e/hUjVgUMVl0Fodu/OuQQ4bI8tzmA80/
Pgceb51nTDFjDFzWWPsylrcoPhgu1IXWDH//OAQ/XEaIvxw6awNiDc2PmGGnB70Ju2oqVZBUFFjE
SeMR9yjXtWx5gSqXVutuFkwfAI86ObwOloyhIH5lBGW85zYplvjEuIoZt8rCr03dA1fIgFhcMJ8t
iBdr6OPxTCDRd9G2Q+c3LZCgxu3C9R1XC/ZzE7h9/j6NyKU4xNxT+Y4JzvFdtpEu8CAKn7NgU5Wk
4kQtr2oxKOEriqU9rLggKJ/L5doD1oP2SeuvRxBPk5YcIlz3Q5xU51exGcLCkVylx3wqJZxJYQ11
kB7JPJOwudvD4wUgeoNWxCJCmUGCHgY+BZfIqSQxHG03xGopSC6+e9TSFh1GMVLfKHT482/I71PR
xfoe4wqoNRWxmuTFkikQ4Tf5PwsCJW3BGK/GxxXgqCBpZjbimtIL/JgxhTU/O9kFtHYsqi9s8qJA
01VGpPeGfRv9X/CP/Gro7LZ7D+HmKOpfAI3DlIc3myxiH8mAkqp7VBtubWt/IQVt9BF4Qjbi1PBG
GRPMXGGTZkL0DdfJgCduRbGmH8EwDMlcpI0RxmIrQv43mgO3sUZvhQJqGHCooks4R8LoZfJswaiJ
KOKer1Fo9/svkJf8V3wItBwMabNOphHDoP6vF2htH4UAUcegm0SToUafswgq9L+rIgc+Uq3kZ05T
cc5bUBJxxuv7zp60rWCKcMmUHtodMxosW7O+OmzUPsZEII6UBxeGC+Py7hYaEqr113QIDFeY+5nW
qHfJcCEkXToWBFRpM37cRmycSWb4tvVT6c/YUfJp81f1G7pqnOyupeWXb95R0drP9CnQqTVX2Tgz
yhyHS9vFcZVL+TSGrMX8zKRLgXIbguzzWIJrbLntaJn4ZgzDfNDcXns0nHLML6mVO8VnwMftrwxL
SEWKYVTqMsIlcycuxqts0L1VRNMxXQ0oT88cx84QJL4GM41wIZzCzQS//G1D+J6f4m71D8Y66bkD
MgVoumDdzZL2YsjCMqIeL2cjS1ZLJuOtFttwDdH89BrBxgMYe3V/gzczFWgIqx++3vqUExMqBCi5
Ogu/d0aHlkIY71qB7hMPKorBg2pBmOx1x1EN4jdsh5hk1iUA6jKuk6jP4bTRcmIKJGPSXn0uEBk9
5h1+Rilbe6GBxA+Uj+OXodz/ad3uDz9DWBYzGTTLSVNyAtydDDhWKrx0o7kO7u0qk7oi/D8M4s9P
kKKzeMQXCDgQYAGFnZe8gFTm7+89mOJMF2CNIFFK8AXu4vXvNdneuO2iV7QGWN3wedUqTlgXd2Et
V660z48+gGeIpzP/RQrgvhvWAnm0l2CRTEUmDvFJEPNXlmjwbfymZWHWlwdL5dNg0xj/hBbb0dfp
eHjQJfK5tFYv0sWBSJpuiLdNW8ar7yH9L/IradjIzOqBQRei+2xOVGMwou/xA1zxzmWrgW4j3/1t
d0JnnM1jx0PW4V9StiJEuIZriBQ47SgAHysLddaeE2FyxYUS47TkJyyOyTbEGfNTYWEr53728TLv
qDZP4CyLHnT7iAD/r4WnH4iSCStDMWteGh75bVAk8Jca4PbMm6ObcZlrDcNV5Y4C0vaIGFCbXzRd
tKR02BUSKBWQ+M6PQRVBZNVCOSPIoulofXW5iR3YY+S1Zn/rMEc7QibpKRb/fNwxiGNqlmiwoqxk
iOlFHbgQ+WrKKDgZ/I3wCklf8SOVrpGacFnpLltnSsFdJCaA45P8cQ7u7fVnq0h4DX/DJqEOM3pi
PNNrDPZfV/zyxSd5DqFIQiVnAQeQKfQzh8z58ZvjyfWHtf05fFzvNjH0ucGLNrVtp7n2BZ8p007o
Q6TS/k0BXgGIv0yJF9PvTgTGt/215HaUkeKciDg/RCIusNvtTNt+apgwgSN5q7l9J4QGPRPDQawR
PMj4wh7EZeAg5igtxlwChjs8hzi0g+VayKBA79VMBW+76ip5xJ5EJri9nZMMnBEdoalQxK3HFwlj
/rGMCo/K+sMwDVnmMqa17sA4+H7SXJwcdMT3F9nGeIVGFOHHxl+IEzBgpjQJSGnzobNhJfegrbdq
iO4PwC/gQMqMAHGNW4I2FnEbU1SVq9GMoRmo3jIdvB70cSw6ycDdgakMcSYkRWw9Dxlx4jeqUSbm
L0HR8ljd+rkm7wNI/+yj1LSsTiJE1BnNQuWICmkbOq1syYzYSZRuf8hp2oal66Y00uJRO5T58LDS
AkzMPpxhAiSI1cD0yaDq7TI0Uxej+sXV9vOZ2wumUQFhbaY+9YvA+ujC7K6HCdQIFJ4rO7Ee8Gye
+XzvMjTOgD5uucGSGVb3umd/hH++45cVUThoGBsqyU6vcVWxRLsGmhfhGLFkFJv59LirmucNAFsO
ZN8vfgoYQ0YxADsvIcxxetzlKC77yTlQZO1wHsIzhNR0pUbbOvQxoDMVUckpGCnoVxyPNKcaXRs4
JPUcyzlwv0U/suak1+5tnjIwnHl4SkEL00N2rEqPpLqKcqqS4l/Ks/1kMj4VJRrXfNNyTzWe3E3z
B39HsLKmYls+B2xQukmv01zPwnt5boc8fogwyQCX4lJAtEyDsnzS3eM7IdSnIw6Z6QlB5mtohR/K
7BV841p54FnAdXiNyyxKZzUnN97vqrUx0SfWDM9YDJ8KJ9+9aduBLEQfcZyc2azQvRzlAu+8e4Hv
5TuSVp/E4xs/lZdb9nm8RgdP8c+jcg5L/D5PwXH/PzV1DXFLS2Yymww2yQ9SrWYyb3xlOYsxMiyX
Vkq+QwOwahvNsni7ISMntOS33jZ2bJah0JV2eJyTZO5lJr2Dv63NjyWJwthRbqV+YshA/YS1Mk99
LgcGiOOMugr3G8gjAFRkc8OKbt8gNUXkdSOjQ6V/pv9zyrdAF9mubdLqxcUIOYhn6s4M6FhbMS6f
dFSgzO6XFJJND86GwZ3K8CSuY20WVJtslk8YVfLlOWgj9Unwp/dVbrbLTc0NWdKlr/kVC1NFDNxU
fD+417AP0I9FTEyRslGdZm0SbpVRkE7bXnoDrf0KBkGieuyySrS11HUZYP+LL3+r3x96buNeKmol
QCYhFlbOEDfjV3BSvYpgpvknZxNM8waYp8tHTcN1sE17OyAwbC6CF4bsFagW4MzUQF6zgzml4VDZ
YPBZxxH0zIYuKRMoGxTCmVSusdLhaHWtIaOlczfQlty6B0SxvQ0+r1xpwIVLmoo0k8q1dz/w0rbc
b6VpILEwkpKtGU19akoZLsd/GHACksqCVUTjb81iSRNeA2sUb4iSygRVweN75Bsag0AvvLaeqiIR
/ytRBxM+uslgyY6j7SnuFnDBSbC/qURCbUarlRvMvM0CwWhniVPs8v2686U9dAPJLkIAouqU8CjV
mtCVS8mQWgL7ROAOVSz/t2ENyMqq0aVPXRuOs12s9xSYRPTIRzM1pAdziiqibGc0TRhp9ZW4YDwH
rKgUH/0yIeGaihK/NsIJUyFiHvhu6OaU/436EMfHKAnIuaE0spXyTCaNbjKTw5sps2MMLpJr1Tky
2pySJ355xw6VaRvbuoeHgyLtDjN2f0jMWNqYfkC6uNu76jiynJU9oURXURvAELFcj5xWzXMo5pat
X8aino5e+HPLLC1PYCWQsgS4hmGr7/eHKwzUQxMBIkrJiY26L2l91B/3JvXFc1F60LAgTvCRzlt1
CqnwtDNm+un+VYYQpNilgtvhb/Z0UfeLNto7luelX9Xztw1U1QwjP2LS73BNNWJ2fpXdtL6FCE/o
b5jLZnfXF8yCX17r8S4SNlwmA5lXZQnk122C3ZqaYZW73aI/i8Npc2m96iwgjibuyUfgoOniTnkW
XN1IfEi/2lhclHJt/GR2h8duzD3Xz0xu0zaBqU9glYsmn2OwVm2p8om0HziQQ8YAwmO+m2dW7PiJ
GRcK6VfkfFaOBWAnWE0cRDFWB09dsQ4k0hiBorQ5i0D79tpRLo+6QRkZESrOlnCepoRBaR/kL3I6
IRNiG3uLQrKeeGxS4E/s0e+xAfBkJn6miLMVWzNQJIOaRItYYAaGpGrUft1zGUB1pogoFAmcWgGg
NHQvJsLAuRrXZfJVLJ58/S07us+9iZ3cWYBEcF9ZZIzzgKjW3+3RruXMypS7whKh4xW0vg0DyXNY
mZcBt8oDDZRgSpb7kwnQmlcSsGhadDNx6Y4gJn1UxKomgmhxeBTr8E8K5Q560e2nr5HdXvipoJN4
RpTiDW2iCzyEHKbJP3a8qFawd759vXOppGMhpTxq4UjO+dvG8yFzwzBdO0a1A/8O/Z2Pu4ECbafz
UYrLh4LAc7OCCv0YntiOSWgD0gKFB9rP5Yj+Pa3hKkltNDS/48tYu4vZmQt24qbb/Gm26L7tVR1C
k3EOLGZ+CiVchQIJkdSpFwjU/gjG4lQnJEVnoVEG5cZO10+pBhCqsmIfexiPmFcNrJ86OJ/BGT2J
bPgkrt2P+spFyfAuKQ+gFILTYqTNbwFPC6bE1GLwJ1yB1UmKzqJvL3egkPd70nU3wQn6ANkIeU8q
/KuQQlYOGNPiVWf7Z8SuHbaH/nv5ucbfr1Po/BP8MW0krpsAZxRVz1fjDVP73f820S+IxA17Ev3w
ut89yrMihZ/Wku8vssZEY1PCImtWEzss0Pt09i4ckYhJjWsp5ctOwH8FJrwct/5em0ZkyBRRe3uF
asXGxVn7/IrY6EPe7sXiIH1ZK55XqphMCeTI3O16Fs2SHcI75VO+fQlWqH2bfYh88oaBl/qTfNhZ
Y2rR0dyQ5OGlO4wPKhl25tXN47KTT92OTfndM0XC7sYJ4ee8r0XKEDlUxmE5vis1IMvxzUCob4gu
VvCun/ldnpN3QAzsNvz5vELF7XYufvT0PrjA8TTwb3dOXY/Yb9/NpNVlGwRroDudFrQvPizkqLW+
K0uSqz6/1Z7h424DHeQppZkznHU5X6Ly4s6VwacdvkLK4DlivFRnG8CZCaWyHfyvptgL6nLyDKMy
12fjg1GCTdTHMeOHDY3fkEgo/iZ9+P4oMKXkbdwVftVk9OgdtKTldKJWXO8E2rSQX5ZxjVQAqA8v
tKsTk70CIt7DbvdqpC6bntYcNBcLVY+uGYkpiVwR1yeYBL1jaucMasrlge272H9Bm6Tgf8/p1D8Q
Qhy9ZDQKUmrMqfm/vt4hdAzacYYx7Y2Ux6DC9xlp1mXiuBcxSuaHTEgJMPPP2vGEa1Ui6MI4/SOZ
tvnjP/gpAfNf2hFByHVPEW73FSdaPzeVEDqWhjAWOaGQeWhgGDSUqVUvuAvs+ARUJIrbPDGO0o5b
v3eDfqmdDpJvDAvG1alXIe1bhI6qyBgFMtzT8M9pRLMKnuRoJfURybn6BvGBji2eEbbBJ9HXQ7Uj
DurPwg11poaFXNZw2m+1l2xVHLVV6Pk3Ub2nhCupKe/6xqJc6IqehEdo7l8sjE6+kkDRBSssxh3n
iiKBN9BANfnlEG3ED9C0ITCWwQMfRd86WWeBnxvpWKJ6KSObZSG7KWmhoq8u6IdzaZyJRL8gTDLx
ybMZgj7QedPLP1Tw9BjOI0zNp/5YXs1vAAn5Jv9ARu+zq+gQK8DmhuggrrhjcskD/BnRKxODwdp5
MufOq+ZKYqCHaNtlMa9LMHVilmJm+rtMxVAEN6Xtq9ao9GuPFKlFTjhI7XdGKrxU03EBK03jA4U5
91RGAI7cDX9OlYG7oGIBZZwI9ISZ5s0+yGxAwQRcttFXq4AK1HvJEcnTsPGA60ZWnwpB23OM1EKj
3xIPVZazzmLvycktPPv4u+PmUNlsOoEI2X5xCIv4s+AlhjcEWXmTv+qfTT3ALxIVQ4T790TnPhlu
MxHXgCF6iP076F5D3maAhGj6QuUJ/XSJC+5IeDlRWNt6ymGmZgkVbHYjXlC3cvD9glYt853Orryh
T9AfRwSbeJ5ia46HJee8thgLISM3NQnoVjhEHSRy/l+NEuD1PqfJ+hNaDWmg88CHCzvaQ3lQmJ1l
/eLlkUggl5DTU1pqwRnPyN/bDKp7VD3pdJXQV5Q27hAA5qr8VR4U5Os9ljFIMDFAcU2euMEzVegA
yV2alHyqYDzBuFC0Ww7E4GOrZK1kklJyO0WoboN7p/6i2nEivzoL9ivlTKeeWBsXSLiUEmNqgdK6
5jEFIMw98VDxzAyRjI5WxXIY2RhiqMk9eFdmLGLxaz0YrVka02VNDRZFqIfnq0kZwvmUsFv1UZrZ
zQFzXYTFSIuh2PIf/z9vWjKsvAtu166KqgIMTfbm6tXQ6vVjSLGlPUJMfDBoHD/zwTFqQvqWn/IR
9tz329j3ejArBGu4LIivLQAbFapEnm3wP+yvCbCywJ3vvNhFDqBjPYNkAGGfvaGUHP2V2V/PPP+x
ew0lj4/L2MAUowRfHa0iMxZhdGBhF44wcSq3tcf8vUfEH5MAgahAu+zxIL44U74LzNdZkvvWONP+
COsuIyAyZ5qdSjFynP7vVMUOhTguA2P8Yq2XozHpndfYLPceY5lnrsfEQ1zBw7YXLHrW0QFM7npO
TI6GB6flqwpBxTf6lr11DRkXJ2eaEoQ879bxqLOJXHjznsyanFPZHINSyABWFkH/Qc921+KTW7W/
drFyLsJObbhi3kNAf6XhH7B2YVILM3OkY96fzFMqUtomjtF0WC1zYV4VYlBR2aTUhzUJFIhvjcnJ
6OJPnweuTQHabo0QPbMKskZ7xJB7olSH3hzgHnUkX8dyc6n4iumS6B+GmFdXBh7OjfuSPeagH0x1
55Q0yPGNUxQicFUeq1i6Zl/vO8Cdqgx0NOjqEl6TIwMmSwKJ7XNbpZHzo87lJpzYc0AKjjmtScJU
TVA+aAF8kE0sDORUl60nwN3zYZ2gIhFASXSdEKWd+4XP5J8pBWyLcNjiAFJA/JBn/OmqnnWklj4L
xnB8T6HFvl7mipexw5PMUHwSfxRNAuRI/Vte4mSv0XoHIEe9uOZlv4FsZI73hzeCw06QQRPM/awS
4oxvQGiOG3viaZQj/RRENjSwnncKGi+9SD3m7Lgxfx4pBdwbFjvd/Yx4PedczYVuuUTBC483+p4p
f7DWCKkLn+k5IYVLtum7iE2fIjl32tCMkEXW8DpCRx6CQ+3NLjUfgZZfYM/SKPVJb5IK+HAnORnA
D76IEQ/IHi25bD+0cAuxtfp1oTe1HMVaIS4z6NVLRcPOsDTgdCYs2b+lls1QNWVvWlenPFT/q16t
pCqNzNQXi1GXZVGcqC59NyKIErw0TiRB+8TVyjBOFcyDVggPFy+r/HQ6PbSLBBiR0QNKo69EFxjU
kucJtQK6one6HitfuWvooriDC5oJzrSn5XQzbVfLnTh7Vl4pSrWxdHRSiJty9O2yloD3F3o4DHyZ
fRkHrH/4WhceHwPVMnsU4lfnZzVqG3fYARcfxUthR8gxJD2xjtu2j8tRv4KAj67fWJTo0UrNJB3I
ya/LzQwiWtI4C7VjGvZx8B/EH6fenYhyIV3Pvo1+338y2A9kaC/n1oezKR1Kn4Wbx2oIljwNnYcN
2fxRof77sxwlZppb6z5hUudydk3+nWDzxH3LneYDihSae4r0D/CPmaisV8ZwrqgkYMTyEv0v/SLe
WNB8X2FApsEo/dcbM7Y7jS06wWDPZHNzahcvJt15BaTugYCyGofkhj8iDZOSfU28qqN7B7RqPw4s
nIt0NFdryi29MpxUTF43BJU6UUut4Lv/0KaRd+7EVq1xoMv8iF1TXxGHOdR7ghLHof0ZDY2Fg090
y3b2fLzeybktbmJE8GDT5QS0SJQXkB+1UZF2VBgitydsso3l2aJw5zH2Nv0xBZ4ImvuXKDqQDCqV
fvxtYr5WVKTxGKfUybkr48qjgtsrlMKNG7rDD0BOTDXDA6k84F7cyzMDL7m72SnKllDrbgZVXzku
QKdz39VclTZRG+MW7HZL0Xz1zBLoG/jDj8rxQbWe2aGOKkJD+JROWY+1ROvLITd88b54CBRh6ckx
o/+oGQJRRc1QjisZZg/8GUBerdrbxLsN5q/Une0lDB6PFkEDaL+ziwXu8NUrAd8qqpXqLSgytyn5
ZpiEnfI5Lf2HAyxwiLPHt2MUuFdPSH+6jID/whkAoUiYkQ1c8rQVarPRKmIxTdrajktzhABiG2GL
DNHinCx9GJTeOaRFHizMsbtgnTN+b0ws9aZtmHb+XW66/5si+OqWWoFqs261W8H98HtWQ0xogADa
O+nOcFmP0xjfsdnpCePf2JGGSgMnL69p2ZEYi60RGE/dnAdBXbee8bfePge6aq5GHgEUkf/w5Qt1
tQdqio4F7l/03N5Yu/96CkiWUv1QZEND+z/QlC1XiE6ODeEjMHvzTgW9qr8Nem6v3to/brVt0P/6
kbndufHMQPjyvLzV+q27+h7a2VGo74n5HcWWUlYowAvS/PHkNnvfiOqADhSoBfkKkb4kgz2pMSX7
eM/H6WeV4lBkx3v9lRo+NPsLcJn4lu1gzKpI2lFS980CEnZawUwCd9qkuqeAUugSJjcX7kQS4v3h
HERMEPdDCarEjL+yXOr0zt2YxnFyhPDZOWKLBDqegMMP9XWvgDAuLd/SDSQmoiYr7aZqKtTRzp8g
FRh25/WIszUMeH4cT3XooTlO1NCJDKt37l2cHNvXp2LYTs8AjtagieiwKuu8J8G8BI26evVrjQjV
HEGQyjlr534X357uk9mQdDLOQO8yp9+42JaPx3LjsOectHCETyweCAumE2biYMAsFqzs84bRKw4l
byhdhLReRIg3ra7OR/tZHakDmVcAhPX+OzgxlscIbNgVMi0Bk0OmnZ1HNuSA7FhAUEFUSsVelfc1
ibBqc360/MxSwZrNbklvoIUyH7V+yLpfNV44TXH9888z/TXVrHK3+t0U97QyDdDoAGxMynhQ5Cws
jFMvvhrVGkpp7gW6QBHIk4mqPdHHJV6enl3zhC/e62wPEZMp6U74+VPIo7ceP1h0UBvni4DLPF79
bxUqWNb1HUw5fu9wVRQfxaFdnEGLftG3RmQeNwcpJNbiAq0js7wZBV9N4q57e6KcAeJRMI/77Wgc
MBvGO+1xEPeoMOE4ek3F0uzvF4NOGsRU3bu7ZoFxic2baPZF02OUY0MULgQkOLTrSI7EiWDJgflV
vFNgMdURolQeB79lXbnddb9P5NUMBzEguRIl6Yv+a/sMDdm43MI09rFHJcLkEVlFE4EJ+jn1U8O5
8qYuK5KNDvsTW7Zdwi/1CQfNEvhIejXb7nTGP/zIhPeQPIk34RwqkN0e//m6hGeKNkjM9lm2I1Jc
1rrRwqVdLtqQ4Gx3rF2DxMIvp+L2y5E2duW4eQsdvTqCkhCFn+zdN9bu9R8fj4FW/LjC0vZ4Hssv
DPTa4+TkX5EZuzBTVrue+PJX+gs+1w6X3Qx5h2fToYW574e9P8R2CKy4ApY+L3Cm+SvdvWvgZLW4
XhrJTjqk/t52I5A7jagodYNLJaiPdDQTD+kr6CCA66NnLD5L/dRFdhajiIS0iwubI00rNfmIpIx5
TD8uakqkrmJOthN9YjKW3LFdbZodP0y2u4/wEx5WTDlDy2MsNrX/iHnB+MyKAMYBb1ZXg32CFbT4
W8sLqNW8Z5nRv7uOx4fi1Rj1GguDJRUQujxvnMBSh8THVfY6nBYElqXslPEXr2WdpfY1s9GYg8YJ
lnWrpTnR+E0U5dSjCjJlGz7YjOa1PjkGxrTdyalamxx9R3xDIv2hd0lGbD5/GWJ13N2jx0/t05M3
YzCUCK5Iwmgc7pqQLEcbRjS34e/MM83xN8ZgSOJRJkzHZ90nquhXftq0oh3EOIOwtMEFqKiENpby
xDU06ynDiVGuGbnqDGadf9YHBhSR8FgLCSpq8PTD5k8fyTpAwZDytgFBr0bAw4AWYbVqEheoMtog
E/w1Wh1jT1qjESD8ZuUL72LzSnYTdgByIklGEc+FWJEasBtLmaO2wb8Kjrset+t5VOALgOyxQAkP
4Z1P+lzyHtsvhk+cjI9EjjJOLHtf0dRbWws6rmFZPTf8NQBfTiOIEoSTjBMolcbbADGutmDMk1Mz
PRwrFRex3jReo9/WJTtDdZmIeVp9h7bOHWiidHL8YsBx+31Z9o7VbhOBiNzVo8CgDTe+FSAsKO81
bKL/EmGnWFuC0MMrrsLBqd0vkOHeyZ9PXjMwKHCiBjVGy/l5cCnvojqAiUpGVaSdCJq4NiU5e5+l
Ibp2Wdyit1jYMXCAuIMjUf9TkRevlKJR7q0aL7crvyifebf6jEz3JIvt4epXPpvFlQrHF3oH++/R
JJs+FmBWIWDSZNYusdtX3Ene60kcq4U2X0A2/mH1/VcyfEqKdNbs7Et/AfbaqtH9D1AJw5H2PM9g
m0P6XwRRAw5B5va1BHor7J/rCDDFSeRgTntib1cbIB2jU3BU4gU4PUMtwny8POn8m8K9JaYJ6Miq
RlkhfwRCeL1wcdiJ3aqdrzO8TsuztiTYgb2HU9BRqEDdOlocZgctdd0zoRLGsJ6mWuGMWgl1BYKh
5By2Psv4h4+CRq1QZjehBWQwAaNSQNjq9I3ULih/9vtLMMcBr5gAsirWRV6Q7SgAzhxFcuuQU3ND
Q10ElN6dmfKECBwaJ46UMf/5PbsElhzb/70eQmV5Lz+dRu2Cnadtj8NjA9wnCBxnx37hwpzfoa4R
epSBFl0+1wmWJqwI5eAiIdqq4E+LCfw/Nj+re/98mqLGrqvcCcykrG4U9UdcGnocSGF5ajdJAAWG
zUJTAFGV6f0jazrnH5/ytXEUNETDjj55C/pMlUQzm8M0Wi7N3i85rdyLbApBD5rXx606W51Q+dQJ
a58XC5GDl6BqCYKgICwcl8siLSIBrvtH18MXK2g2PbLD+F4TiZBLVrHrmJt2LQe/poL9rsGpetde
gV8PXmQ7pf0a0M4GXpxC8YkZguUeC9bAQxLt0gguPGgq8bcia+ogIVFiMwu/Qqa/7vNQrKy8dqeQ
prcD2xK/UEGUW57SybgFXWz71Mif+Isq8Vza5SYbm8nyxcQoaOeaGcu774IiFQufPcx0FJuz7ElA
yd1kmKv16l6XKVdrbds+8F9Fsnt69MO3Ts+m0BApmH1MWGOuWcP/ZbW0uQOUYSAu9xmnuredH+Gv
wyPDWRGIsgsXLWPFHKt47CHYNxmcdKY1OokwmOO5bv65NWVdgOaQTMjpBxbUoZYu3ON0S4y4SNBk
u+jTmzPctobl0IE/Tl8UF7VbX2SpdTYiqeOzrrnFXWd65nb0/+Q2JwQG3Mt7u+FZnUw6Y0HhPGJ9
hL/vdCnJNbqKBZqsvTbN/9yyXFK2wv95RGYAylIziCZZvhJKdyoAdLdKvpORYI26ObH+zEEPPpyC
tQpjYWOO/lyYPU294BYevYaj9fQnTuo8ekeOQGLKrk2he4J/tswwaW+csNzpLe0aockNO4OG54qa
8gAHT2ItswDC+Ai6mqLN1LSh/4Eqwy9eWfD/6yP02SZVsOOwFOkfuP7pEcl9UCu1IPW10NzYn3SH
EbG1MjXkQQ/C0S51SLmey6A+6yEkyfZfltrUT6SQmEaSPDbqxGnr8JfJNAsPNE7t2hLwtUd/ASuf
XHOarhrqbPSl4Oyzf0aFfGjVM3EDfwbIb5j1JsvFb/HWr4+9QUqrxT5i4ScZ73HK1EnoyVIzlaXh
tZYbXzPTEvxbhxTYIxofpqB3Dyvn+RO1k4mWZflE6xPjyD8yUMBjdynxYylf9HNSKeQzfeaSP3hu
DtzTD2LB8PKJ9JTzerkmHfPiEwG6rd1StgCXv4kJrPaqXQoO/ArqEjmmAekYAjWNHyJzXbOVuAo3
MDbt8JzX8v1eughrd5AAX5GhNJcTLBP3T3ATvlI5PJALqhQRhNwqYfEtPbferd3HWyj3v46j1qcg
QeIF8/6kFvmfIw5iLw2etCnVgOIoFjySxCayqOoZ3Teh5z8EtpV600XXABr4cZAp3PQz4FQz/T2h
R3skNSY73aq2deNvVVhbCTGqNV94Llak0MJ9zVynhosTr1GgHqzYyaOEoKXfEYct+f418L5kNY78
9/ctMmaD357gGXeNqYtynM1W26qZHVby7uRpMQyGXd+OrdS4B0USfHjLIJ1OirZmX+G/q4aMdWMu
hf6vvCM3QnExfgmmzxKleC0aV+6J7994//dVC3wlx8FXfIGvrMWcM8wYuSnikfnuQMRrRa5SNCFh
vl5yfFS4gpmPNAYdGA59ZwVjKYbUDzSCAYRBk3QnRzFOn2B6NhObAMspYlAhappN24sxOHdt/oeV
lxGEwYRwgeIx3NsEiV5iSABaj5PgZ+fpHtUFWrYFgHlur4+VZ+4AJBvpH45fc9ilnQjputpWXRO/
NLJVTXRbDxPivOQTILeA6eJf21+LGZHiFS+jO0dWzAYv2asiSiE4Sbrf0vWkb7OjJauIcPpU7upX
MI7mzceVdnewF5UM54o6z3c9Sj6LjY7RLsq1gFTDengzLqpfMmK2R79vruIW/BcNmb3Z7NaEWcL9
M8jehfORdVKYLxtXUwbj3PrdnYj5MOjklnLeUjxnS2Z1/zYim+PkZCBG6OwOnJxpR9iMh5RR70dJ
CW8mA+M2IDfPOxIUMfK8EugLsp/NKe8HAIJgcC2a2Ae8G4zK/sClUy/1wZlgLj1BksILl4iuhJfK
SHCpbCwmrOu+akoc1gsPMUV7VuxYUnkin7CjM9lGMRJp86/d4/zAl/8gXsKIEeD/aQdWz8IeKno5
PkLVNZ53WbQMEVgtbSxt1UuX+U7u9yUfaOZzz52clHjtbh5hRAAmMIGsWs6BGu15kAopb3A3CHPu
APsn1sOLu4Gfwromoq8IQhEg5XA1HXf77nkcb0Pi3ERhnOwD/oFfALkXN9HxMRbv6vDWj7xFiKQu
rBITfQQ01PLEuRll0i5SmfgQjac5FIpi8JCr1jLcwhMXMMnEA34ybWWHrxeAjwlZ8VltstQ6kMz9
MJwlTos+cC+OWLzzC2Qzk8+uq3YjIOWW/f1A6D6eYbfyyH9HqNti9con0XWOcc28JAf6W0YHjo/b
mYG/n1HX3gxPTvDa8V4YPVSaW2U0FA09lh9XXwEQDlTiRDAwJ7+igMUL6SGPbfb5fro87RIOTu45
WTSOBcyO8TatZoJX8S6D8CJfZ0pkldQLRynMECTfzFVMRvAptLbxN+wbkSIGBZ+DfnEXVYh2MrR3
3WJ3dqIcuu17WGeA0SWIxPPd0AgOOkp6QS35s7541WoAAiaUJSCrNM/yA6pwaUZAS0kMiYEvvLJI
ZRHYYZCulc+q1GEkEEbI3uGsUjVuX0L9yOjy9yeGoIJnII1lL6QidVDLC6nPpAjEe+B2bS7x7el+
bsE33J/Hn0t4nRuqGcM4KD9+VbFHBzyekQ76TAi57Mj4wcXXJ+hK1gw1ckbn0LfqgM/UMHBsreTh
XRpPMT77X6Yl1PeapCR9Tkzm1s+lXRxr8mLxT+Ba9m1hwQOju27xEhy3wXnZ1scRAF+yjNxiVKqw
4XX+QqNcScE+lihVZKnqQwAv6f9d6I1SwKHkd87WCchZJdO1NAvoDMxwdBaWmM84212cYJ87dkoK
AHNvU4SAY2TKdPm7h9XmU7MrFLeIeFEqRM7GZkfO491AMSafDAWy03AiopXFuWvP/Vggoe3iabMR
mrv31T0tBaTLQK18MDJ/LIbUDHGUeZsAl/sRoQNn9utH1ZyiXbIKO94vCjyAEtROFk2vS0D3a8K4
mx8HxCeX1jCi8bIEqhyccVTGnJhHSW90nqujISFXH25xCqjY9AHl4R4jJUilm1V2iipB5v7jtKQH
sYwVe6i+Jh/pnGw3Xx+1aHNh03ModlB21NDgZgLh1KBs9NPg4vICUN3m3YBv3M6UF+9xtIvLXzXe
DtsEF5sHPHz1d7oR9C2GrviRfDD+Gq+4aQqVb7HWIcyglVyowjmBgdivStklUYWjeQvpGsE8Bis7
WlUtmOr9jv/j2ugyL/yF9GZS46DKi2BRDZk0M1nHPG6nAhsxLJKILHj1uvS8qGiBqQVGOafCjHmi
qxjNSlH5bt/f3WKxOy5uTzFBedyqSFnpyOMatWp7jh3Y4oZz77RDSrywcNzagAf7fBEFLfoBE9V7
FYJ4HoRt7+Mb6xnjpEhzGqhOjlmw+qwrFePlHgnTEtNpqrtxQCewweNxUfmWNHyEmqVh9nCgJ0UP
VQBAcDHgFhVJ8VYQs+egJzUvN2XZj9cuBQgde+5Q3AJz44/QWkgqdaiC5BVn2Y/ZaHlML6a9pVjj
8XbF31KRJl2LRoZg473BbSn2XNbiChxBZDKEesbCmGy62s0O6s8qThqKRlxxJbVzfqTRu7YBTw+T
RCXqDDgTnLCk9yAkGmATnj7HNXEKS/p2WcmN0OVmEKOt5cMILjhAxcftU1F/Lxu0cMP1mpCRHTPL
FKTvHDEeXKdyylkI400YYYYAyJFci+VVbx3YqqBfuQ2Ei46TA0q2gUGUAWb+c5czzPdVxyZ1v1AJ
ZHDNGFIfif/z0I4QUXT0SVh362w7SpGSAQ37BkMrybaZ7h0wpGFzWYZWkMwvhcdFelGQ1Q+eBUEs
pBnUfSbjLcDF7XMBUkywEzKgAXl1LDspNp7l41TPjZgx/x97ZEl1qxe/+ozmOCRvVIhkEOH4xGIe
7f68Y9B9TX3okaJWS55wslLGXjvewjf/zlBlu0eOntl9OwfR9hxmF+h3uIafPt9wgj4a9/dmv7L7
/+kvVM8Yzs9GLqdyThJDPdN3/YvCZZ4+OTIC5ZBtOJ6Fo9MIMb9eVxYyygyk8Q5Iil19WCoYlppQ
PmauagVmzLqx2uE5FVZxIR91Klc9wcZ9eJBbMb5AakIEnTENeKu56fso83/BPXOFIIE4XOcQz7Uu
90USGcT4uBBsAVjbTeFT55dM7uSM+LmDzW77G4JnTZ6B/7s1bv2DhE+Hvd+v79AyeIrIxwtyTPBe
HznxrpFbpcT8L+1+Ge3npT2I7S2obS1ZNrzzZzFa3bP2CMkAZH0hrfDEXpB+f87mBM6VFyBsVgao
Ntf+AHdpSGzfjguBgohHUokP7O7omo/iJkHNlpJGqFLjr+gigzoT9XiRW4YF968lcRaSlG/cUu7q
163wg3tIR2QwCxpE9AIWgpX4YAmixXt7ssWO8zkkGg721xhZilN1TNHCTcN5lbyEQABozJxnCn57
Hih6SxboZcOlFrwtlSeiAzuiK8RcOTro5pFSkQKJzIsG72UpzbrJGhPQ27DLrsZZS4Ouv/AMW237
REFXGxzkK0Q0UqrA5VViqqgC3zcD0fzvzsRgEcP1Hckd8G2Aq12pCeMkBorkJTgO8WUEQ2ZkrXnX
UC11JuBL2XtqUjNm1ZnMnukhci3C2Lv0cEm3e0YZnlU9yA5CKmZGrDbbpETGncqJUlVvaJklbX3x
0gd9/L37eq/rrrNvTkraqBCtlZsYa1Qm1cw7f6jXOVyWz7y08lSfuIBgFPNqAfYrQ9dZWpJETDSN
rX7Y42BIwrzzT7bpZlaYybQuOvF4bL0/4d6Os09dpkcMeznQEl/wxOqRaNPmPKtYvJj8YofuM65t
ifZ/V/3j/MnJrWE82GoYJ3QhzLLOgTAihdNEG//oeBmb25iWscF1Un4OXXhS58Pewz/IB8mqYc7c
kDgsAO0f2OJZbYsnaHIFvE2rQytRy0wfrTzyt6ZKBsAf4RjxzPtZ8Bj4SbhHxf3COl1x1xpJipAw
4pJqEPIPOxOHIc++tub8R+WLRDuIPLKkiilXYrlb0V/ITPbxpiQsr3qFQuI7ywgpVyaiONcuL2N4
M2CK/QKZsxPpnrQen79eqAOl78eGVpVBoDN4el1+hPFE0sDz1iU3lRE12proVHPb7NI+xhr4/zrp
hJ8AJPWsZPi0My44/mA/WehbwhXIlXqc1YWfvvE7eWx4JcjM0EEDLtL4GqPF5Jhtdv8ZkK8Dmh7w
Xf5wcHBYG7jPjIqUnBtgRRtT+BBSTj+3kHk1gUk8MyAsKVHKzINniV8010P0JVOMJOtJdhcD2XCj
OPnyKsXaC/7heqSs7KKTtAKWRtT9LgZQ5LEM2onKnp/CUa+pbIMy9j4P2W0sKVOqb1wobxSxtFiK
UHY7pytGVp4jLknlz5quwrDZwqicQs9Shu6QKhPU4h1zmwLQy59JMC5UuGuwtJ6C/DqqSzV4tO70
hZIugSxyD+1zqHaOwxHkmDqrVFbJCVOXBCiwlIdwMKHrx4Y7VTM//BatlIhQfyrwToGLZGWonvhS
U6b+jaP0Mhl7rM7077QGXY9Vl6om9C5Gyds5dZTX/t6hklW1VUGGBoKzkJ9xWMhJrbKLmYRtYOSy
mfwC+D0qzMusNISt1JI8z02vjlpejv7tepK83EQJRawaPj2XBWTBIDEj/ppMGO5PO2vpkLgzSS3a
Iifd3Jojdyekusw/Q3kFvd4XMyMbDWeaCIBtGNZ/ST5SK8hMqKUQ+m5EID8OURDLW25o32QD9P/U
miKglglcl0vfHYDRB6rt0/9S7VTligvZDZ25gkgfIAkB8YGQ0G0HzTwOY5vGuKZAU4IdUoVF5PGU
N3Ja4rkFFrI27kKIDyINNstsXWE4DfYpyZg5q0v8jHTNMAYpojRVym2tu8nI1KKKmcYGEhFoIdJm
FMfvYES1i3kK8r6fAEJls0EvE2sJVwDNk2Ynn3L8kVxfytvGxPmY+G9qn+hSpE3w7RSndNvUbdFU
ckqZPMs2ztzBjxWvmcxONVlUHZMjyW8dFlw8ogLwczATzSSPRHlD6Dqzj3us6l/bXrOEWcz/Cnqz
8WqChKil0uJ93ogESApfmGIXFQnp7n9HfZYK5MgwYKa6nKqMlgl7vpNFL7+BSr1s0MzbOn6QRkoT
LasDXi6/9YuY7qYZZi3s0DXekKUNMToNv4+zk44R5L4QOAXxvR5haW7Udjybl06ZmgddRJSIqedC
BkZiKvfWtp1C/iX0qrQiiOqamSIoTX8JiU+5zqbt7dRUlIgPte3r6+GQD/DS3Orr1NH6Tc4BfZtw
OtDY9UAoLAgsH3gj0eV1n+tMVidVd99xbxZDXsMYpvXGdcRAe24zPqUvYqK6Q0NhyxDWg49iB4dL
b6Kzmc91iBojIz0QNeheYTvceE9Z2lwwpP0sSj9DSDXsZ97EFIMZBbpnqMvqiALqVcTS7pj2oLU2
E/Iq+BxC00cjw4xz3RsUMk3xjcvZ08fhoTut8cTWQumk37p/Xbg1ESiwdYCkIGqx1fBvhaRGpvoG
Cjgple3cgz5ossVvWlPlwzDPZ5kFE29drHSAOrLOM7YEMzyjYsPYJuxj9WS6opZ/QzC/cHI4Zu7Z
iuXU33DONv58voU/2e31zhjw0Vl+NOesBbpzn88QqHqbuqGVHg0fxdxP18vp1iCpONq/jE+zMn9j
lQqOk8ku/qLSRrMj5yzfGtT/AKCpH1jQSQj7/pAIh57bZA0ZQajmnz2ewuGQ3JeHeQjAKLl/Kv6Q
tfSss/kjQlW0NVu+lcOU/BcMWfw4KQ9yeLRh6u2p+KzHMdXwAh7HF4P33PnOi/3ghRwz+fX5DF1s
fKPh+ami2J7JW3iBfUop6kToGDa9PHYS2JBohKnC8aSLOuqaGqTJMEm3MevZg+1Piw+25y47OMn8
Q85SpEGTgq246LdK0c3Bj5zIzDfYZnEf6PVg1eI+qrZhse6zF5/HMcHVVHyz62k5udgpDfUp4+wJ
pvxsqby2Uroo58jMlr2Xvm1TqYHTzXWWr5mWfQckBRT/HNHATTfZjmqTfnBOrPsRoJx0K4U+K37m
zXOtwpiAhmrb6K9DvRAV2faTMEbV8sYNY+EIPWceujygTdncHUVJxqso1/GV14cz9a2ZWqtI4h6C
jVyIVm2tuf/QPVtocakmM162rcUcz6HdiFiw+Sq+fYgEpr3iks6ic44qV+AXw5gWz/xnysECY+la
YJZ1NaQbKVpDOPQvHXS99VsBUJOaiM0XJxn7MY1O87WqtQvosyZn6yu2LUfmHN21Jab7pW0/mCtC
JFwtSKXaaZzlBuj9sAmtZ21NO8C3vV6pY8MR8dINj7HUZJlcp69uRB/aA/KW9HOppoLpVkouAyBO
pYY8y2x4zLomASuSKjlw4SjyQaTq6N76g6Fd+hDfBUZIOW0TK+D4lLQGxKLCMndYK1Im7MVqWGJF
fbfHq6gi9kkiZR9pnFvrDhOtYkMpsxWmWmmH5f33fYZaag+PHiaFoQ/91Il8MXWzhKInqvndrBJ5
j4vg7ncXujmqhgqPQxtCQabMrlHMXz+VNxsEgh4ftn37Apu5AXujcjBqh1PdZTJOB/W5z/eOPWIc
BP+DAyu7AmSjiONZFyFFItPcGynOXwcDK4OyPEQINiXQwzTEXnbtBuaPli0oVQQfbyRGTRyShrcB
vDCjyM99GSPm7x7WYYTEob/q5/7Qa5l2Dn6UAb56XYXMX9UHoclifQ57ES22guKRaOwVV63t4EW8
Y+uJiEXTGmy3YTzgeZHz/UvkoO7FWRqRPa0Wq1HXCv9703eVN7ZGH/sQKrQUR5evqF90/NoTjQ1F
kPOu19TAA8reQrOrVR9GXTY6qECNyVjNH1JYa3uxBk8LH1qxm6H06Xd7GLHQowcsOuzgkS1kW8nG
jHphDdZySxsmaamGqGC3ld42SkKXYA/94xSoldZZyu44SDutx1llF6smEwZLduUITmHoiBZzqs0r
e5oVrK8vhkx+b+8KLWgSmwc2kPA9yvLfJUSNj69AN8zr0c8VyHWhWq35XzEm6PtHKBp8gaxRw5wB
oysr7/gFve9Pjsq9lh9cCc7AZrWM9041OKgt2gDRbWQG30s++NWrejDnUO+sV+YIQskh1J59D1Ep
87k1ub/WOOos8AS1g+zXs9IrA97M94k+yPiewrVye44+DXRQ4VkpGQs9loGcmD5b5Vr5iheIzv+h
tIElYFPc/f/w4lOQy3/MvkQjoART+RaS2YWagBGL49KN1dX5t4/ymNsusihJCTMWSFm83z8/nyUV
2PSdx/3/oNZ2TD8e+/kAE3DAJd1XrA0xXP5OirrD5dcIbMBZk2RZ+RoIKKqkXpLazlpd2eRMtcTO
C8Aa2bpWmFyuiA9e9QeeUpIuiMjM2kzia/EIYsrxjRRne1WZjHz5MMINACczESZc1nZ0FtZLmQoK
lFy+72TJhI18AA2j7LrY3QQgl/VvtPkcnZD1PB11huDvWdSbSFH1gAxf7WYcYD8Z9SPCxUjZdLpb
hGPhQiyWMwnzIDJRgc6UTIShIKHUngOvk4gIPJQPvl7IwGsibSkwyRdSj3fPZuWKHYFx7rRvtXJR
2tdNX1f5yBN1fT/DRKnayuzSdNRJ4MGL+ZfYhEwrd4XKtkiyx3JTTSZtSALs6VfkH00jWDOgkYvA
QZzsvA7N5S15Ty/XbzMsyxydQyWoa35/zerLtvUWknbB+SxqDy7xz5fX+awGVH7afrk0xo7d27pJ
U4+q06JUQdAp1q9OZ4UEQK/doyq3uU+PDIyrIvqYqM+Tu4RoAz+4TdaXz1u44mQpCI/IyRGGCMOq
6zfWaTeFSDp4ddE33whk+OcruDqzXsKkWIjutjjdktQq/IghCbiVXGeKAyIgUCD1R/NvouxHU2LT
Ant4TwsHSKhl0JhJmmrjGGd4NJ5K3rFKL1ByyBZLJurWJWKkUg+Kx9l1y+IDckWOugIIE0KhHGGH
u4HcM8nlN3DpICWQhRvDpBR5ARqbRIPKJtCKTlCibZoxC7+eFzWP+80gq2gstjkfjO6fQhg833WM
NDO49i8ElIIbzIF0+itHRAUR70whMeijoIIIA1s6vma4kUPRIhuFshyXCsvtcGBFCbop1fJYlHaE
xX0LbkMTApgeagU8HtXYoNl3SNnb830dPDgQSQ+8b8eHAq0o0+dsMYbfKoWYe6RIyxjNz0VnLDqL
F/yXC1t00oPlrFQUwO0hwa73TBkU9KgJ7ydwUVb3jDgtQCRuf/UIniDAN/p6Kvrg82SSxX3BjhaK
fQ7KOea4rW815BouV7I+TOc8srs5v51sh2m/a0/u5Edu1uIMEpUtZzfQY+KCFu0raL+uTXgiRKuA
WqqYH10olMN+in49zJRKw7EH5HdY1Tvtm2z6hr+FhGFPwxE7spJElebYkX+z1Y2snDFAgG9R4g8D
2dC574Na85sGDv2/ltZSX71lGyfn1xfbfj/XRgloTbgppRNZDUo7KqtIejVMB2RoM2OsC2WnuBTe
OE3e84GV7tRuZOanb/CzXo+4PZ+tau1ElWSkfKd8wPwzg+0XEG4v7UNpwe+Z2aBGI91syg2CLyeG
ptJxyPcO9KtYEyFr8o4/BEZWOBp6tA+RZOKwL/+1KH9+QUqZ+kPb+ZVCFQUtNA5pGPq4ilniby+t
ketG5COWXbMiorwf2yEdN7hCvPd1a9MbQZF/lU4zmi7oPJtJDmgjqH/8uBZs/w2QeoQOHy0cn1cr
1+VMLN5KNHRPjeXHa+T7CcmVew6EAkm3ZbCRi/Vjw+QIUA3+t8+JQ3fIy1dnVSGlUQbMcRXCavss
8kEabj/f8Cj3EPn0DON0Ev3joXaJW8mLh04+gSlHJHYRW3qqTxrYzBbMFOtTSQ366V7SK9RHI5GY
Mmc6QaYa6QhiAsziPRwTWWoFm/ZR8hkeLInaDTTDor6A59kfIbKczytR3sOyf2iD8c6dfT61QmVA
09RUH7suBtDiq4JJh5wllfCe/8N2lKJi8+aVzyeZ/0paVACu+Ljx4X6SvWcBRiVVPXpOPFugxEFb
Qs4z46mz98wlQK7rICiw+PQ01pDpvE1D7uNEG1kEF9vTQjcnuinpZm8tllFIOE15FVfjVcwWL+AR
TEcEUaI/hym76/6G3Zjskgslc0AopkUkGxcsoxZuvcWBR7dTzQZLnpIQ4I5REmRbGQnCFXrn/huL
yhTANbwfGhti0IHC3lOzEOEpP1qDuHlNTpRfKuOSFGgjuWLjBVoGu7m+jWfQ2vcey36UG1z/eCwC
FuyWn9DTH5updJaXsndGp1OWx30JuoTINN++ToREwtpZVqSo9JRet+MjHvv5UxB+CRVP4aI4GEjO
nrMHtIGL3t9pQot8MIJGLj7JvCMACwUFjslbdjW/7UTGtfURUm8iF2fdv8vj4434ZQ5WmerKrr18
gXkINFfL7L9yWcLVrJeNnQQ9ZRCHWl+LbbSerZkXTTka9MBjY94q+nQ5mu8jLwe/inzP4UKHGXWm
JRHnDKAvr61AOjjeWKuvidDvBbvoROFhb3q6/vgJZlP005VZhbRcOGrar1O7MO1qFQnHde8aAkga
StcA+21jqCEEBmDm3nTtfr7WM4X7alhtHkbzZ/XZDJcqPUrSZdM2RyqAY/N7b4HFiVfywXsIuDFG
mYwEO3NXAlOp6KNioRsukAf4e24+gMVWOKLTuNg6R91Lpa3Njmt+z5eSnm4AC8yTWxVENLLfls5V
Pjh950DYS7SEb9Rg3DdUXcVXan++3jBTOm1s25IPX/EDmmFZ36xAOhoYOivjkJ00ycXL91ShfcFU
jUduc4mINJixBdogE8gZj3nZNzP8F9GNik7Hbo2SF9pTP7W7KfB3kj6RUzkb2AmUUeVJ2pLY024U
2ZWkSds1lTrRmMGl4xrub7nc7fFdpuB9M7yrfHDH5Dr++nSreGi7OmaVLLtJJC3eaeuTufzfs7LJ
wI3+qLQ6Unvlzf/GfTOyoD4scLOgBA3+WkIFgrejzj72J+6wRwgyiRaCOUbrKbIycmldRoCTZgdQ
kwlUurBtCWyFvA4qnXhQirxGfVv3dEh9YzotJyaxVQ7bjhN0WjktUHduavRWtpy26539FqpFHW52
05FD9ECytpHMlzCVbtGcN/QZLRAtK8238xkxR6TdyteIOeyiop+pVkwR28TCmE21Ns4kWpkHsB7Z
TXd5VPxZBGsq70f8RvQrb8FaJh2v/WZbmdzcts8nSSvkHVH+i4zFkx7LsrTYllAJN4b03Dua0+zU
8rkjXZ1pItZF/rDqEWZPzNmF1CYjUlauKTOxJJbAWrWI1ED373jUgmly3M0diwI2VZFnJN135amt
A1skxHIFcKr8SzwqRi6eODHhbGst9vaEsOemOb+k9P60HAmXg2ocNu90Kjp9LCiTCdfpu89rxv7+
sGxAH0mjkMf6zHWRyxxukp9Rw0CYTJNtNwANnfaq2XY0tE4B6ZmA0vRdd5tn8k+6F1mmxUKl4gD5
2X02hS1vdIyOeWBrStBEAwGYHHbmcbF4ip8Z2jvow9q7TcdiwGGHzSCm49woR+vrlUY2uHMAWPdQ
bGWOykDT7jZs0q3uAaYv9FFjgPvj9ADXrgWTOAHFg/aqJeEqXBQpsCS4wW1OcMs3jQkZeyyekpME
nJhCKyjZkssd369Kg9YuAg7r7lEc93W6taMSVHPkIKQ35dOBqNNX1dVzuYAVTxM53k0VMNm+mb4Z
HnHHNQsX1HBfUvLMsrg/TKdRmWhBafvP4luOS2iL4meWMgHm7zu15VVW/i0QmdnFT5R69AxMSwCg
bW8X+oM9TnEPc3ayn+znSngR8lM3D04g11Qew9j5WBD/wMzs3d0wbatN71bP50YBZ5rRaOZ4gZOQ
kA/E1FSc2JLh5iOFStn9onkArNbYHm+HhWZH21dmLFvu+3rWLJLn9wbba1dJPbHmUlHmI4nHdrlo
dTQTJshBX/RM2dPI/s61T645dZiA2hEL4QYEVRWF+OkUyQtZBJM5gqVGT09cUQZ4mO/eUrpbYhv9
180QZk845eeAYgQRZc/YqY7VkYANDB5ow3sOLSSukMpxoYPWdX+V9tUOqMDyOZZJyj95uzBgPncA
IPMPIz11g2f8v/7C+R6F55hU5aSQkU+eLiJC4AcJInY9YW3rYwWIxtfzYpHVOj1pM0PWHBK6DUm/
NtJqTyJXDjmWQjhHlG0SoZugrZXfG5WffrNNxac1slC+zDFS1fdgFvcPU8PEr552AhxndBMhNaj4
DY8Eo+cji5+7aaHhr7aJ+HEvDYl/cQHqTt76IW/xQPOUrJ6lk+HBFS+2Cpb7OypZGB/HhuFRDirP
LQxGian8WBidC1O/pgz5AiKw6+RufzQXireWZRhti92KsiC1Mg/B3btaQN9Tmo758pO9K6dVeGFG
0m+cvmpYyr2u5Gy0pUIatYKcQEXIaq/598SkbfL0BKF1zLE5o8xSPRLPjsLh13fCcmclgJCqNCp+
cAQwlOnsRmKy/8vevcDHvyu6KBizf09ptv/Gt7S2qFi4KGR72KyV5RDGMP/psY22Cz2mOO9MAWYe
e+zXWeqzRH9DeMTCcVgTaZohrjc2BdM1NdVC2zQyjbnxgqpmySCkvfNT8Seb3XnvHPM3yEHdIopw
WNj1NXcbBUm+EcPAQrhe85LNIC/ku9zory08S+tgSKWLi/elmGtNRa6KRGNn2PUdOi5UipKpiXqj
gZ4aYlfJ1ZFBsOxY+YlCRz9WKXoTwOAdT8JLII2YgI5Vs7NG66x16MMJyeMChTt48+JCrhJZpIMX
AbI13Z+hYyGvVAI6pGL+R5q0ktPSb1XBnpzUoDIKL4TSc7tj+sl8AkSFfqoqbeyy4grlm3HvdT3x
ZVHS/p3UG/C2hPtPqf11igJNonQ2DWiQ4Vw5P+vDjcjA5wegZbJqOdAbKfgvwEsUg30XZfq0lXFh
rX/16ruzGBYp5aCyKWjVm/oukq9qCf1yvnqe8kuLbrzmidJSPfxbjEFFL567JzRZ48gilSmvDKoQ
uT6Um6DEySZM4TAWrrPqSGbkBgep1/c/d9xtO3HyeKFi+Kxxq9EYqdqUaQGV6Djtxa12rrgvDXgV
fmEc97EtUFtLc9DuJf6Or53RQhe+eqtridiqPGhGUYhnjG09CvvxecvsA7Jyah+uhdP/6W2dt1sC
Pho/KYAci7lggFRsyKqBYeiQkBlXRvQd1gOx8+lxHbzIX6+dFK2BigX0jFOiFReeF4wSHhSbeDqg
OePJ840lchAU1g4vBKvTkD63Ri4QaI/+0gx5s1/9+iIJWzfoB7G4w4yWBA5c331Kuner807px3sr
yzcLEmyk2IDPpEUtwnmBdfUeoXGR0CH2EVm84qiB83xhNdacQaG+bIFSivnKiQp7EqlKPjte0R+r
bGKM2kyHQEnJz8EiiBiLxsWBv8+J7gfg1/vAxNG6UPKZDaQq5rdYByaOOq00BmWk/XuEtB/xPSwn
4Z8xxJdvKZ+rw8NnNXi8d+SHr6EWp2Lvq5UmXdFp7GdX7k8OxsDckfkjq1qFOtuGaJHbPT8gERwY
uDMTGpUReUjzD/VLnUvpOg/MknmDLJhWQ4g8exQa7jgkSSeEhfRwJ35G1XQXaw1sgyiHCAf4TOQn
zJLlUcXY9xNKJDwx2DB57QjPzpvvXGFpP3KnQcapCk+JNG96wqlxQP52RRgoWX0PduUEEQRRe4Hz
QYEW9p8JgJElO2JcsehrGZPakUAklHiWfg5UW1cXoBHZoddhE7aO6vhyo9WOzz5lnSvnROZZoZIG
OIRyoWAfBwv1gZ2AMLtHb1fVPa/TZnNYu5mQBk1+1LACcomKTk87lP8r/q/nLbGM52WMqKA7JiAB
rKHbIB3gT00Mp3IAsAo9CZ37Ofq6e6vI2FcKinu7q+tvXpi/iSnczVU5EGNbsYP1bIrCoduc48QH
5hJqaj+0atwjV2AgNUb3OYfEYHTLHELVqQlZJneQA0xhI/cZ1GdNH3o+IAVZe1MJ/P/xKkJT8CGW
zjWqJwGOSiU16cM2JxCEJWkq53CXNfHuQD3kT4gk3XC6Dc7I3XBuo/sIEQsY3IcQxqJUzCIiRQcH
qt1UBi4exokeO5tfAzDEIgdtIQTqKXhU4zYCqyGJCHQrbGlJ2sk0trddjY403E6JI/8bI1iaPe10
9NnAwqDq0PjOFJfe0oCgeoAfIwHzzTBIAvw60WEuil6adOeLafu9r8qoJecrdh0Vjrg2/aJTTJhd
v/0ao1g7i57Be6JdbyBhKCDEhlcMuoKbgpz7O1pFFOhc3TuENMB73Tf9JwkWm0FOog6Zoda/KZ3b
6j/wzr9LGbdDE2z49ytNjkiZfGtCs76u1/n7XYweqMirSuvztZTfyMXjF7LuMSVthd3h9x/cZAWv
zdHJ085HcW7vZmYw3qHUfEz+Y1z5wleupgpnCxfxf52nRnSxYe6Jymbd9olwhv3pHe6uUSDIoOSd
gkDxmII8k+MFGvM5BKEqbf689MQO+LRrLMnDzGB6VbwJlmBcxZWk/doTwYFOn4kYfJGB3SMcMQKG
v1lO5jqL1gYPdzgTP4yIJQPqhkdFChqZsB7ZsYZ8P8Ki79GBMK02YKfC+KjWc+uSb/a1Qf0iMen9
u119nKyK+OYhaJjW8UrZA5EtIFS33M/cFRBTyduMp50lcin6fIsNS/lXH8Rj6ZpXkTCVyRPQVJGI
yvc07m5YiqFIrnRZJFELSWmo0nICxsqwF6tdXFPvT18XH5eHOzh0hUyB7NyoZNXce8WcgUPG1Mx9
YWUgOY2aa+rjRiLcSKjGuq8DOA/dAaGVRTEbBdIfrCswLvd7+ngSHry0vbn38XTEVWnI5PR3FNEB
0iyANsw7eEq/MLNJKGyYzFJ2t6bkhU2uA0ge+TFWcNOri7RQG8BQt60ETaLDPfxbKBi7+Ji1rtkT
xxrTl5CH6pPAf825b6XDQLEXk6OpAjvq9F0E5lAHdtCpjLxmWmc+fv4WMMFZouE4LuJS1VxrGq1+
UB6qAhuAsayvm47c/XRH1FGb5Ld4iWYzcM/x7gIC+rcZIVWQdUb4ZawYBgflHXBEvPRK/9uCOGhx
VCdvKpFxWlVjec5X36yMfHPedgRlQ8krBygMO6fXo5P9g40sLCTbBhrbRMecCwq+Ggd/W8eMSPR1
qbb1dtTfE+W46tUFBBtT5e6WgH2UVNuCqT3Uw5KdVTHcRh9LmMxwt5QjJy10BqDJKxbk0PG3xCVP
cqLWkAohBfjXMlbXG9DAeMjyKrSEw2MRgIgSx44O7Bfd8I2c6YgdPsskiN0IHrRLdnm0DZd1eVsR
OumFKtnRmXAi/dPm7Bjppct91jOQJq1XgBPmjyyzkYilOcC/ynTL2ss0/s52k1o5F11QANJrcoXm
KgwtVt/njpTlUlWNKbdQxSS84RL/oCuj0MPx9KfBVI8DIW6sbEp2s9xzm2yJXMGv5J+ZZIuH0C8E
aMooRWfvlubfoEgpn/5WUmuEFSIGCGRsJnp8dJ+jiBegQHqnhWcOfb2OlsP3wF9ke4KystMS6KSv
SODKQXWGOt9uXr/kJvFSKsMlptdA3cYanacd+YOPlV7xi6xbvXOjGGxyYuJA/qh+I/48QAmEK/mb
hMMaMnm0kk0eiVNg7fqNZDI1swtX482LKZXjKhsjiHPUpr2VEA/iIZ4tRgqRNQ1CdDlLUHJ2lNcP
m/UR8Qoa7sok+h8rfovKS7gXOuskSWAL+sT9RRrqgHU2DDNabL8NN9QWHKiUhVOxI0ggKPsZsRQ6
bjHo/nX0rGojq8ZQCkGJFC4pFu7x0KCHzLwbskHNE6WPbb3BrLA3JjNG4exDZM0VA8RQ6HA2jIZR
BIZRmiMY2lLojnToKQVR7t8kUZotAFaCAF1uPyNeyZ9Qbv1teZQ0z5E/kn61gyPlOP+OeU7s+NAd
zgx0mmqy7CdbgZDnLnL1X1WC0ATi4+oSlINaZzCXVwcFcGyqSWr182xLOCtvZIGCxPe+77CuQ4RW
F/FCn2KOsxm5mYI6OvXdUkS61li2gAGcZjkzpOP2+WwYhxRaNgH4RIVcsyn95+4gKmaPbOA7FiDz
rkka1qslhrk3O9QdMxBaffysHs+w7OnbTlAqdOn0gWtEEEpqeY61KBlMR7/pKdNyQHZtJ44vPvdM
nUZ1BhcjAZS/6QUbeA/iN4v9llwhHXS8Sz+a6wQZ9pmXiLvjS6gJROXvI4u7dayQKasieOq0dFpW
fv3XhyAMC+Fh/dfkxu9S0zVtB9UTeRinyDU9Ru5HfWxN2QRR8H5Vw31BcBByeb/UL4uNCg7+ODXu
l/8OOxvJO3sbESvKToKJHK4fwr3RJG+rLXX4ACcb3I6oyUa3S4Ykc9SShjErft47mKAaQt2ylmAV
VYGCmrJK5KvQVLi3Tql1U00nrc9m/Of+YC4s3Ktsb+Cj7ZpLr7XmCQOukPRoW7unIeGfYkYIDonH
B5/N5V+Kwb89/NGNPA5RdcP1gJEMR6voU1I54RkcYLIDaCvO/gakgT+Yi4b9bYTkPa+NdUetUbcu
toR2Du9hZyEwU4Ar2gBfkpshnhuEU7ygfmVhQ+AJ1UlgyuPNQkQeA1Km6jcX4ELxWhppkZFXw+YS
3LJIKLjj6MvRBlCRFpi9L6I6uo60+922cPwl0XSh8rEyXxuAaNINDdUPatBAr6U3ZbGmzR5pTQ8A
Tq3nFz2AiQf5RoRKsQRvjiW3hyCOc2eDUOeybqPPYpcXsxoMABnQtF0jDcubSXUoshr/HdYux+DM
vq7UyDi9t1kry97MA0ND63Bh7A3t4yGmau7k2vzyLEiTvw+bvRd3GBe3NAkifa2UKrSJg3oupKQs
QqihENZFmfOTkzQuHZauvMAsR0qsIIwEFYQ3W4zSuN9xpgW/1Yzfl4GJi+Ht1SRr8ddCLGZKBZYO
o48vso6Cip87sa8g/kp1XDzoWNCgqfttMOgrq+dFOBDg/J6dRoNzwieqCNr7GYBCvZKxWaladHA6
in6/hgz3oDutOD/9EXiJfYJ3UFThAcMDtCOceEXv7j8boKkkXanRu3OvEAu/3Yj7JH9JEU/J26cG
xondQOCGNnlnaJz4/v956fpdjIYaCe2drnVNqOh8TsKfQ7y388mJYbdOK9Oai+L7q8Sa5oKA5ll9
myVtDRII1m9zMidpY/ZKEs3IMOTjYMsrJ9OihDRaa8KAzL3VuL+c/5G5XaVPrfsPT0K7LViu9x2h
egvWiQ4IImzmEI/ct4dynYqm2aSRw0hhCbq0Xy1nipJuwi09iO/E1Kdx61o1ItMnR4WO+gfAsjqt
wIXCG7TwkT+nooize97IQVkCi0MJkXvg6ccwRn9tUDOnsxTGGD7q+0thlkPZuh6FP/SMV/DLRbKm
d+nolfle1emOkWnZHqMHJWTW9qqkJu2avtFiycGxZuM54rPSJt+P5+BfAlNxKe0H4cDYgsBJmSFm
fp/eyuTyOisfyTK9sfl4SJWjjEwi6k8SAzkqgwUDEK/+ultC6AO8rIoJ5OsBy8VM3nz5EA3+Rt10
YqJFROKsZvAGXaTQGSv2uRDC9Ctssqt/pXDBEZDZ3JZhRXBs8xna4gbHTrwdvSM7mX4WAyOk3+F/
RvCVAYggjEyJL8Gcyf/ueprZr/f9Xmfey6QVViYuKkIWSLNDKtLTAIYP7mOkzuro748KhmzugV+B
ryowSiSgfrjKIS9ZQkNwKmhJEziYKjDbcCOkICVIloC2azydPazS8ZSFkgnzqcVAy71JCd1GxG52
YzLpP9dbGzh7w6VKfZwrah5TaNBEGYjQlzdvkNr40V0cZmAwhlLeQbhoO6NhRFKvDCX7XG6tvG+7
bscl0v5iuBe8uvHuWtUMJZJS9gwJyCKGvkIWbQyf4sTCXYNvg4ib8LgKxVev4RxqUlEy/V2UWGlH
FgFWnVvjQZzlcGem7Dmwvy6mvX3oaTInx2wL4fSsFY2Rnr6ZDFjZOtfnPvlL0CRfNeHUV4spLiO+
ZfQTnl/Vx/Sg/FnN1m55MeOd1X1IwEy/0KBl39MDsHzNbm1DUz0T8kH/19j39EHB6yXpRCKTthOx
5kUJO0GBrGBr1TyNuLRHGQh/3onAbyWzxnLoAArqH0Os9+lBIKlyx3u8Lwtk5ZmYizdCHgKI1IoQ
LvHEJLHtgl+dpZGMmwY57pXCPwXweQtrHMcsnl2jXO1bWB+ere9Df6A61VxAgHmi3GvzEO1hjdat
NF2cciIhqo9zEe8paafG9pqC2bvLGsogMqOJ3VBQcyxqB4DXUj9mFAGY4TnuWnlavgSR8gE/EXnC
pzkNvLddVoerexx5ZdxCHMtjXU0OL7BcwJyVMu/Bnzz7kI/6WPGe3S4GNn6bFoqkfi6Samcjp8+s
GiYXKM6k9GvuJMzAJC6ePCl2bRt/z9suPeDRN8gQmBts6fF27gkxLwK42VAra+T8sWFMuZc+GX3Q
Mz4Hb4V1epkUDhcyOsO5DE8Q3iroK2obqvmSWwNbSCy8swr55i1V9jRf53RhHDDyD/0siuHdctyH
hgn0kYOBLgxExHimrwIlYASqpWaIFzYtguen94vF2BUqmkMV3bj9/giHaWZgrM6++G7BIpcIJspP
ZPdo/GZVhqY6NZigniOmqdIAPw0F93BYfnj5d7qqLIg5Kxt/ZwaRUtBvy4zp/HXmYuT0O1FxEA5x
N5V5svzk/GDfXr18XQjbkST8FzXWeKAXuzKzKYKekwzgYvuhDwn76HZ/xQHwfuEJWXDmp9it5g9L
iTNclZiJIUbYhbLX4bvD3LiUiYrA26gZM0KxCibrsOkizkIi++o0T+1KTnI5JlfN+baRrZfJmZed
FovAbvCI9WNm3Q1k3XIDTgsfWIjpbH+dKNyvWadURWLM9oq+NvMH+4NS5BBIHIuwUvWYgZ1l0tXm
ekKCW5s5LEp+ljgLC5iBWgOcoC2Mv1CMrtDjLfA45gtkycI6FqtFS5qwvSYlqfyva08kqlDt7vfl
M0YyV409Sa9JhZHksIs4YYjnszrzSPjqk055LRA6R1ky0n8UwJOjADgRh1klG7fHnocwp/1Bdg73
TPs9cQODuoYtBQMHFGPzNtdNc5BluSq+LNYOrOYve8EJ9I26/czAQkeeIg5RJ2NeU9WdAtk3YZwC
8b75pbVtbIiOlZ+FpM2ooJyxJu+gDevFxm6a/wOGk3JapUT7vN7P6aQqXOVdZg0f9hKdvVMJBwQU
dA2WkJFtbhih53BE8XZvR/V2yeu+MwsEvF8MOg8qMUpm+hNckRyl/zbc2M17fkzmQCrwuUKDfuVb
QG3IXiO3uUO6n3ufV5q8ZUoSCk8pjfrlMWa1wkf/39VsT3mEoT6UjICzGVWu/ilozRnuZIVluGiB
sCyEaBmIVPbr+K19bwZK+SJb7FUwaL6G+scJyi6e73iN5lQjWQ74g9Hg908Bl28C4KXYGhfTC6gm
GMQHilYJPHRvi81qTEnhuD2gvcLIZH5plX98W/nhvrvRBsxK1kOhfVKh0B10+6nuAGRkZO8Ygg6G
IR/FeQWxjlDqbqfAGNFDBYXy6mr/1ytPo5UQ8yKsTlS9UMg62RMsfIh35RT+FS7cm4gndqyiVkx8
1GzDL13MQmPy0/AWDo3aG4gA8Eh890jtXIXkSnN+HRBnusg2Y4oyyJIDVuk/8Pv2j9xlwTL+z2iK
tqXOSBJ6iRk/hltBw5iHhAmkdm3sgIPRuVi95tq1YHyM6hROPswJwUU1bZiwbeaQ9f5FFdZowl54
RBzZ6Tuq3GjvzLq/lk62yeb5b3ueizbI/jDTKrNeMOIIoBKrPbuAMsfPrzndwD+AUXLW3lPl+OAj
qFy9jg7MUsbCFYabGpsFpfgKNLsz8FkDba4Rb48Y41ysF9/qtbgeMGCgb7DS3ZrGagoi/lhSK870
pA4mxnORj19W6+AHmTkqJXuJIV6+xL7dVfIgHv3lowICyyGz+dAHb1KxFCAlzL2YWJ8imgRySgC/
V6g6H8+MXTgEb7I79uWiMx/joGH+MexxWzbBCYwsg8d4GCCIgrTZv53JFKHk7oPhOOuhLz6+2goF
hUhCbtjZzio8A/I3vzQtp/R1PmV+rvnoR+VlfqFemjicWHhoX+CrRCZ/CvDG8+GPD6fiIav5Fp0n
1XZWfEvVPaui1x19yNrYAYyWDBVb8d9FWpSrTvcDFTEvHqxPnPCGvzH0vILLxxF87X2LCMWvjePP
JxRBTMKD+RbfscbCWZKPQbEYpXNJicSkdDQis6OAfRUq6pV/jm08JsqHYpC4C3dZ3YuXVSmfxupS
NwLBrVQw1wjc5R4pQ1lcXuNlu52zrDqWE0J0hUCDaNQO8fdFRM3WZ3hiNVS1nrD7juOR/FVymQHf
qWC9yb+uu6ok4olCJGrEzfyqZMlXoWlpKLjMHIalkh0Dbvl+R75HNstQV/ZuYuAIob0jb8mis1px
1JqhkvAMTl54fDEG52EBDoc3eTQ6EE7mJ8aqifEKRcTngzhv7rN0HqaBgz6vPIBX+3c48QM4EqUb
Py7b4vDt6rAhD4d7UNDTxS0yCDp92tDVaSecdwrVX3g1Q9iQZseeuKGwHOBywgGp+oXeitN3VFbA
4dN6JQZldICC4j19Wlppc8sMluvkmfAPG4O9RwVulJi2M7NydxZfdNYBrEEvATCl+YPpAFFgzZ0j
RKcnqYfeBHw4299DhXn/0wUTdO6rLkQkwmvVs5SZBuYvbXgCE8bY6EXjoUrHzjbvPFOCTecyftzb
kiign9cNN42KrOFiiO1QEJZ5vWlbbExdmPVMBJ/QqGLO45WsYk+XRpFzhE5+4QYWcUEVT/2eL38s
jl50nVyBjpfQuCW+IJZRGudj/aLl5ZFDMDj0avJezVqyBSTfKcmRLdQ/HtuYolMcyWxLtxLq0rE4
4VIp0ZmO6XVa5c56Fz5Yxq4HDNjxBgRbucUUicVqv4IOFCchIRg+VE7d0OO16mq4ONCT0ikw2lGz
g4vxHOh/wjkpFYPP/UFtfSz0bjoAH+B2fKsL4d/23MrwtOmetNFehITT7/3pcJ2kIVGP5/FX7yCk
9Za9Jza3XNo+4I5snF5aUXQFAXbVE0bWeoDAKXhGiNL03YQh7gsdkuzb9ajqAaAiSH9KFXRlnqa5
RuhQzvyVhtQ+RK4ly0Yyi0nO9eBHq13nomgNJR+bOSZM+HD5936PMQPd4gRvy5T57dYvZ2VoQOhA
kZSX61dfH6yRrlfwpVfombkxmnbGs8DA+ATFRtFoCQPiUFDcEfW5DZ0fUtkhck2jLtDBrkHz5Q5J
+tudw8Cda6+CC6iFNqfzPadVKBBnrDP1u9cZjPAwySf1wvqMVZ5GpXRYYpxiJ6anyjBHDHnuHtTB
uMFIs2a95uTeBUpkQUpmkbn8xi8sINOzH3Zz4zxGgMVbWaoyo2fzWjt2QQzABEStGzKFswJ7p9ms
fbWZxD0a66pRvVLV7nC7PDRidD+RwSFmp5qyQBxrnNhkKj1quu/Zua5eZYcwpJodqP2Jm2F0KC9K
D9EH/0/u0nc2sprW7PHEk80fNJzJPxPAo+5x1/azKdTQhONjWcJ4+4jNZ+n1lr/d+g8aULr+/ImO
h7k6etG2+hImvUhWS5Dcp+XPr3wvbxDJpt06R+gzQzNePdbBig1+1uOldPjqshaKgK7KyAUCCa3T
P5m7qkePd/acmzdc2wnF+zSVP+x5zrVZBpYWz8c8QTqLBtB6k2EFiK7ZPGeQ9LjEQ/YR2FEDoZqt
XPXn9TQ99YwHP2/HelZsNFhfKpYFtwlm8NJpFuMfRLSQc3AxDgukrBPnax8GqcPHNffsb6VTPwXz
gXkgTyLcE9FEHyObpoFZxp9/aJ8mmRloor3nqMwifVUebMbTYQeEGasnxbMQujhdvAKEw5FBOzHl
c4Cvv/BNFoDupG0DhqbZz4O40Q3kXvrP3Od3Xyc3qSLC4l84qlKf/EqlztRk2uoz5cTABmyhS4+w
XOjf8TF+J+MGmDLV7bwN43gqFiug7OccamQYHWAK9raGpIHkw+21f7QjWD4TR434UdY3NncOmJss
CYjT1DRRu7s0Bl6wgzkahiRii6KgUvxhlYOf5aFFyG56g2FyJsKTxqLyeGR153Auq9CKdMc/7eCH
cLOvngsNlAwhtQgNDIxvg9Zcj0zdzD/YCded+/bipmlPYwdSNWJq+NvQrj+FfH6HmZcKgHls8zrD
0Ip7TnEYTnmapnkkm36L0kU6Yv/uM8FTmA7oe8dl2Q49HNHpmJI626kLVA5QGFlik2RqE3hRZO6x
YtXSfLdRHQgr4Go6WeLkpkHL6Znmc3wPaoHvYt338Ub+LFVwlK3Q4brUurBdJt5dnKC0mVBNxyHr
UnWw35eooAS+52fmdcB7mnqFOm8c0vUR9Psb5dGo+WQIkhEmxyDCpvdz0cBjDejxru6yMOV9HCCn
qv7xxBUX7EveNC7A8zuTBhNtSLPhQBjqK175Vvj5TVjsdRgbSfZofdFltpYTWLd8RGF1TIL4v8Jv
fInaX7ING4uJipdQ/6d3sHHg8AI1xCdJdhWz2CEqSHnMtTR73lh0jqsQjMs1MbFJGeFjSMKpSiKJ
PwHl9Ch6aAuWKy89PqdNJND3CQ8g0LxPPEKFfV3GN/UlomwG7vPe30YEX7CzWg0ERKCtzvdy9p0w
tNclqYE6xRUVUh1OmKL4LqxytWn7RniPlTQ91cSikhlylSwV8FaaSL3+Bo9E7wLZ59/BU7lv7Dt3
G8rPWubYyYeEQo0eoMGbEF3KGbDUHCjxLFANavhSNMCSWJ5Balfafl8RZcTfr3YXiy6z7sDWj7jk
Rvbbwb54pBWq7EXyJRHWqNqUSOFiWh8UhLqFc2R7UlHqCPf4erWNpztgvGeQ83Qg/4Fz3APyLWPA
31ax1nl6DhGBmydUd7ppDYi3xL+cBjPBGHa+0RcMpkWar/fMtHKQvJKX5I0ZnyuwxuPhJy0Sd9In
iQ/tXucZ2Uo0T/QzY4wkbwwJPh4ttCnegwrEICu/4VzwbJccDDPqUOHTk+MqOyv8RUyPzeC3RbDC
U4qAmiwk9KN9LvsSykb347q7vl4fjafZsPPUqS6iCgj5UpbpAFZe+UCVPq7AMuIoGt7kBKahJNhs
qMmLXnen0S6B8GAMnZ+h4dq5vnoAtfgpmjzqZI08F+wsHyyiH2gHkuT2KDKwllUxXRNV+dt686j8
46WL+JJT4iIgNR+moT1IsQRrEs78pODS6d3FARhG6OM4VZLrMKNvvLjO01cl07JNJnOhesX+GCO2
0x71uf61kHBAkm7yyLyamASOSKQ49BFDhv5Li6Oj8idg4UHysUvTVET8jMz0frvZEMcGjFEN7e0X
ZriZESebtgGS/UVStYeLEhvWciyHTk6ZpjZKtBphVHz1QaQTF2YgZG2DR//cQZUl3tnudVzkhPYy
aBUbAEJ2Db0PPigrovCiTOlCWJ0gszft3AA6WmCmX3wt77OcpqI/EwXpouijG4pPhSwz46QIr3O8
uquVTHVhWaI1EQDvzpj+dNOpt1RqDKW315LxYMyqAd97a3chBiJ5WancyfIgy3tlJLOaIJB3cCF8
4dJ5xNpvMo1u8E7j/GzxYs40xjY3Vsp7O/CYZ7j0v4d3voQbwol9EsvydHaUba1qukP3DKWbplHJ
WNTkWIrdKo0+59QD1kL+18cXRBOQvtq8/0H5Oq1cimZcA8m1PYzyIcZOMv/3wWrdlbhd9Xx4QGLG
3lz2MsBw8UuwOxLKzVbyrH3upn3brpcKvAc/o5xaX3aEq8QnJiJVbF38u6K+Q8NC6uPf8KoMk50U
fOSGhM8uMF95AmrZO3R163PVuJNV3CnSsJ8mFY+YBL6ujkIHuWohykjxyGxQbFM4LM10sdB+bxi1
PLuOEi+N2pY/z8MtEaFLt0DW9fC/EXJActRoBmejDwbkAkXJWc/CjhBgGyDjFqaMitpWEAcIaDYZ
6D64oGA9q6OrW9eqOplZhPPn7jXMtYuZVJ4Fn2gjtmDX4E6DfbAFBxa0a7P1OP9qhVDCVYsQh+MH
bNB0aOiF3BYUSFnhEnhqAIgv3sgDyv0pE8IdQXUgihvvI2QW540GmMKFLO89+Al2fqNWSEKZsQxu
is/D6Y7lmka/B4aJRqZolBdOJeZzusFG3Qzg3+Ng/Xob4nwxPLklTlWgB1wHlgsko3kgFvdssxXj
V5zFlGBWdpGcjn3tVEq3kPmoU9bx+Uh1FRvDkenHN2FnKXZNVfy/HkIaU3nVrViU58DFXWeRypcm
kBctxK5Is4oSnzNF38ywFPEljQyO9SE1T1q4OdTMmLIGgEPtt+SRybod7Os9W4rZcaRnsQIXfLz9
VHuCLjKbp8xqa+ugS2eXKeM2kAS1kv47eVTDK1aS5lcrxyVc1ioMyatcbLPC7ptG15IzArPGmzK6
vjVGEGnrjk/HOYNZqDI/5AxvU5sI9cX7J4F1u+fuNFX7KeLCtcRoV0tU5u0kwbBDC73R/+WyCu6/
JvBA84mpFiWU9LPVucnUKQ/FWyzXS5Enxv+7F5f35710j32EA+9GKxUDOWGQnIc9Hr0DSgBqJR31
oSPzFM5KtJY/dM/wVUR6Bvapxvp4VQ8geq08riuwDtrICsiZxM6W/LzAqPC0cN4JSuFSELFTO/kT
4zAnIiaLv2Ld1aaKlRmQEYFTm0LdUYIqDMDGHUgZWZoorr/Js5p+r0vJl+Qhsib9Pg+kkuMQmyxx
Tdh5OGMyRC9nlEesxTfkhr2meQ/j3dKVlIT6ARbkVj6O1jVvn4f0BwQLnTxdP2ooPjNTWCmZk5pc
OyTL3olptYJjXsztBoBhly/+UjyndxBGkCENeZcCG+1JpeevuSPH+ShAd5onD4oMQdA5JKeIvr7Z
op02Rox3e58rMFJW8gH4fB/3R/zVi7F5pCt655HGarz6qfCRY2RNze8P/YfH8p3a4MvlYBeKMjNI
a4bQU85WEHEriixSMRkLkkP1EfP8Pqpy7qg902gPrSpjsfiSP1tmBML/e7s1MsocktDnLZssICX7
crGjI6bicq3z7vpIUlF9M/UTv+O7VCH4xj5/5NgvaG7KjPEQjvqvH33tjIc4clhzO7QjcbXlFBlI
k+fCPqbl5JgV7p70r9olvn9jApoyM7YeULMQtiJI0750sJeamAB+KZi26JkdD8zSA2Bfr0eed3hz
qIjOpgvHMV8MEpGiy0agxUodDXJ+KhIxJaOyXYsOqky8Xe/+rnqxwUP4f4lnOqKV6oTGk1zAtaId
51i9eNPRUM0g0Mcd5VqHelcefBvw7aZDB65511eAobjDsPc7jHl+1NMVIUoMTk7aGHscgoTA9eG3
n/m1PS9wD380S2YOkJwWk9PlQuZ56iROqCWa6KVNKE6UezBH4DIP/zjlECu1EPn7pjzC2yN2IY1U
WLKJXKLfPpJ3VvNhBjaEDKrC9jT+vU5OQ2wZ4uvvj1DYunCBWURfI1MxzF7qCyuHcNcjLwrorJqz
UXSkw9v3R2jSGNwKQAnZBc63TD0878VXGzOyl+vWN0YEQfggfSsPa4H9ExGYhNWsm0nNNU5j+Na1
vmtQnkkmpPXk3oewQ+CYhb58g5UKrWDgbdhs7R+CG3ADydUvstVYa5RzEBh9cgHXmSvs5bDvS+5G
bazXvSKy5JVDEwczLk0tlhu02viyqMELGriRuMYQtzicSJitUH/kiD1r++WcFtdtlH3078R1gQYf
Vooivtlq6E75Zov3BPBYNPPcByh17iQMIj8yQ2ZuzlusZDYOIcx+CTXaaf60Qk+G5PnsQhA2byUt
9337zLg2qRFnjjMbdZhMJeuTRjtAQwozm0y4JmTujxfTkPFnfBPHz6t+2D1RbwbEhtqzPCXduhP/
R/eRrOOmmjkevaEwYCQves3Yu5Nref+BC0vSGOl4d6NHIjmzFc1zIplIhcGNvs2GiwCWYWamKwrA
nYUwBn7G6mmZ2FFt0jCNuTtYw4QHYoZhb4Y/2yKLeVgSRYWKejKoaE/NlzHgd6CQNfDuKoq0zPOc
Ea12sq4Dfk+bxd6XdX6JILYGhhBLwRSZwFEJb+guA5mwekgfIWu5Y4exWzTcAHA+u5R66txw5MxC
QICoNb9z7svY8gtxJvHpQnAEcPdLP6+kV9mqQ0r+qqJ+yiqlW2D+Z9YO53oLkD9dEL4dD8ndEtXL
yrt5ytkO+jTlOjgKsHwUjED0Onr6ZvOkpjyZhPAyHExYw/y4Q05+nVDM3VRZ4anTbZh1n85jBsc7
n8ZoLJhKv/uz1+h/DsNYhxTk9jy9tY0Y0EjXpnXsUxpAzC69Lp2inFxt8ffq2rSSEwvVbBSqqTs5
Y03jcubPpgadd0BIruFJGQtuiy0JF7wYS6xR2WJVjuC18dlR9Pk5jwsI7vbkc1t0UxbXYKhhI0o0
uznNDC3cCuh8UWV7UUV6OzeKxZjsLcAVYJQJnrsDa5Gy6LRyGvSWPgW0cTE0BUGMsLvykr5WgI0H
aGwcIdaPA7mxjQZxkVdMNZ83SOCLFW/UEcrH1FkUBeYv57uWzWAkMLbizlaYx4JHAAdJsPFSNSG5
ednrAFmlxSbyHNEvKr/kx2tK2gyngXUZ/tQn/i6hCq8mt9Wl5BVcv9Yv7RnKlRmQDP0nLLs8GZ5H
B9D1RTlAxc5Q0N3bNpj7SY3WR3NYrwZQq9XCiQhPXrOfBIN4lsKbmsAEp0mmgUAXo3zKR5qDoyAq
Hj/+G9KFcLa9bGSHD4J1RXO71+frvmL2hWki0LKbqx5+UPtVHrUGH9tXQSt0j0acJ7/MOKEIFGnd
WEJvwfYQF1NS5yheRmpDEdnI9hVV8xyyB+fsJBUNAViYy3mlTkytaKQ1oCWWkd74tmP1QwKwOuqm
mC7+PNvjcOgsn4p5kfFCtEEZc4YQeBK3xLTo1IEUtKJBUlfUYt2Nz7qJQellrTmV30SuRF+JeQQ5
y6XbCglourLB0YR5ChWjMkC5RuTZqdcqFmEuf6zlLJoEQ8WhhjECCg9Ja9j7mL5WJ+wBl7/nH/km
/zc6a9xr+j6a7mht2QiYbh9Pxw9uAwq+xa8szmQALCgJtZOHqXGj85KQSLljFsS75rIO9Ni3ei+1
QjCmcR1foJJAXepGJ/h950ESMwBP1iWfQdo5u+JLQmF6S88UVbuV2+Or/k4BYNieXN/MfWdhhlVc
qPwo2Bz1gVRHwjYWBWoIQKBjr3E4vSSz5tDO5KAINT9MSdv6c1x77iZkQyejsms1pEakHyXSdrZl
WEvsB0uQ7tq43pFWBP8xOYnv/rvYfQ1mLYDXdgIAD8Gq/Fby+mtPFglyxLm82hszWtcgVxX6gKxY
Lgsk8E795I4kkX3GtM6e7JyKNiRBr9gWi0iYrMLYNHPE+HdYhBaPvEfT7wxmAI9konr+S2R1xCs4
QSRSPKgcT+4/rE0er+A7Erhi4FweLd6f3VHfGnpRL37L0zHF9T2UiZmKcQgqrIR2lmzhQb9d/AaI
TVZxHqXnMdT3a5YcimK2MJ8kseauQTlxzR2abXSaW8WL2DTGaQ4rzHRZTgBqIbAgLNdabO6d5eSs
ZXzuAlexwDj/ujksI9i5grIGQS8tqPF7uIgbT/dRplxS7RYV8aah2VADsgxDZhQsV7s+BZT3gVDG
ssTnAjcdzeCVnTgLA8hbO3+XAtbVEGD4bfqIiTWy1lqoj5Ndcm4PNqFlVLTprFCH2ake3ioXWQt6
XBG2PT2wopDvh4kXSCaVjhV+SJuFcRR+94NXQaC67xxbOr0+EUPWj9HdUxaxGuDnKd6RnkRi7AMp
t6uD/IM0Hj0HrxCAWP23VakYcD+4HmvaONk/i/rYwyCs/6RCA7olCWMmmOiZSCv/Wn/hbEcsWKuL
1VrcZiXcBwpT4aEIumFh9zlyoju4D2uRJYnavJXmWnmRA42T86zawmbj4al6VXcIF0xDJusXuOm6
B5mv9Ifci7zDI4K2XC0JxJm2Vyy30oOSgMbXSfRQXuGPXRLPD7iViYLA1Su05SU+WtjpBN+yXcn3
rnx0ZSlJ0jGcSa3qWK40QBb9LDnnIWcbiLd0Zc6gzpgun8jqGWwKDa94oMh7y8V2b0qVmBngTaEE
cNZMXNXVSkTuaKNwYfMQhjFjDoK3M/TFIXB+3JWZK3fhDzBYrMHhyaTxCr+im5i3UpNdlY8eAsmX
9McWw49OXPqE11Z04qfu8WtRe9hc4PnRzRZT5WiHUNRAJbsnwOgY+/frGR3GUrYntCRZ+ROjP3zK
1XqS6iky94S4P7+p0ZF75okX5l1YjmavM4pqcdEdyhsYoAi4z1NhpTjG4cFzaB09vL13EdbMsUQr
MdxrW5iMfqfVrub4GEqzrX1xtdGTxuItgM2LkPzAe2C55cV9wN4L4VC1wXwCHFoY/D4af4Atd9aG
4/6iXpVztmnzOO0WJwojW1eak3/kdDawsE7L03h6kXNFlWY2yIfWkd+r0eA/Z1BYvgom7jOvL+D6
9txmrykKDUQDRhHtJ5N/ZZIzbuFBI45QuA3rtBXwZwPd4AOR1lfnf8skDrTM1iFFwNcJ3LPBZavC
LHmf3nwZ0xDu6g78bTpcHgbMqPnWofgsqsvEcx3K/qhJaSKUyyBI7NI4LuqopdTeR7xwohVaXO70
8FMO8nauc9TNt0cTNXc799A9tfZ9XxZmJb5CmwWg5W6osW4PIql95RPPw4G4ZLz4sH8xl3CKKwtd
0nUvUA2PvKUYEO0gNYBIlXk4dbL5sgfdjqNUyTfRqNu035KVbUG8img8zHTX6lklLMpj5KI0vC7Q
5NeAMCFJXOl4NaxdrCE8v/gXJYob5siM/QxoKnsZsRV3CHHbdxUO52zkOfCbAvF+YM0LzSErMQ4w
hV1iVI5xG1+imbwDueBiIJUZ7NktTstQnloijwtwX/wdTanv1WAgzyRhrhXwPyaX5KnIocc3Cf4F
/tR4wwZHImnxeXc7uYVT0i0KYUqDQ10bBJGLDn7LtM7LK8lfTam70KGPZ6Zp3yICtVpBSjx96qAM
WIOYZ1MfhgrEiv3eMCdr0fRvJnS+dqkOIMWRYnGHuJnZV7ICZEasGh75zDHSN0udXIz9c72bvXIS
KBWFBR1ZC1hH6wHOdAP+7OdRwTx0Ru8X14WE6/UA362cAjxzWmVaJ2qi2JqU+Y2REgJeGBz65Icr
UtmzqrtsSlPqlaofaGKYN0suWKu4/gb8ab+yRPNvujmgci2QrvahNWEbgvKvqOYIwaBRcOCKbRQ7
Y02pfIREMZVyPKNANj9t7DZgb2ShtdFcLJ7ZIbw63d9pRW15GNDHEeg8k+ialJVeixiNCbINobBN
fPGVsKi09KjrIAtA5GMi/aN9PYDsH+xddmD3bsNKxXVW5PLPH4eAeuqYcrfMv5SzUgomXHtM//Nl
TqMbJ+OevY6dfYlcD1HOo3wQ1M1cDpx5SuLieU2d/LO4eu92f4NBJeiibZiM6+U6nNnPuOQFrENE
ng7m7TNaETuufKA3mMqra4Ze2PynudboOmvPUc0dN2hL1gF9wSLcU4qJDnVhE5AJaeCH9EXM4eXo
y1ZupVv5NvEf/POpIf/81YBSHwMy8Npm7OhguQoUsXjgHvVG363yJJcrXdsN0EN4MeHYk8lz4DZU
LCeKCylDyttnbBJT/jk2kg6Aj68JbfTqL4LNnXRX3AOCyZKJS3GNRW5kdHn0FBuS5HL3AIG26vQA
mwJu+Qdt9s+UKN50qiIwNNLWizTiQXNzVwckLIIjaP1aiRdSUFh2TtmFdnJ8jUvIWRyliMJJPd8V
S5/jmf6lR569QdCADx/v0Ya1VYSyFlkf7e4Z6n9doIwaj+PyjJ0YDXlmAjry5oVdw1jJWhYAX3p/
sd62Rwteb9bky6o4OdrCCATTy6NVco31wBcXqD14rJK3blwQ+t1bRxP1q3KlgdZknPFJFeb6ACUo
JpMGrhrCe2t0YjqZZPbi2YKgd84Wd8YHFe5DpGMItesIsMxN4GypX4+MH4/POzwkTV6Sw/F5mgUl
c9i61APreDGBjlHIBhC4Ed+LxYvQAcFiBZj4Cogx9j7VNrJ6l73ffadzMr4M1z9dpXLkNLrJ/7gk
WkAW4y1pnO/e9hUOmIo1PNJUb7KSZzsZGgVX/kopv385dXI4Blf0heGz6xOLBZrjreyIpfeQivzB
pUKx0QRqNqpfEyytkim4Dq/ltqB97BM1/FUVZixzOeVWnigcvnMoo4gLs4AsD1b2OXae7eps49TL
//rE5HQbutKwitpGOLIxg89hG3a8PKJVNn+jakQgHkhVKRV93WWh7Q3u2NiiNGHtxV/riRTukueo
ihJKrSq7L37JGgDhazOoHPXUSGT9B1TV4lNxTDZMx1+t2F5KgbqvbCluAV45VK7uhTs8CS/A92aT
5qAsNyC4YSSCP+tCl/U9OZOo7t5yt0jUgSkspTLoFAUnJ39B2gt3BKRNTErTDjlQFktr5BTSXvKJ
oQxYvwAhXDPpRztfpieTdRbZgPQlGOZjjM/3YhfHmldOZtguXmjxWV+eI6ggc6LGDRwW9ldD7rqQ
b6Z+r5GnEGJBq4LKPuLWsCcA0jns5+NYIyN2r52QRDri+kz31phlm23uHjuBgIhNzXiF4bMJo6Ed
mtJDh7ZQwfne/X9KiGt6BrVivPOD8hj1YLS92+5ZtyehQSQjTUaNz4pM0nXD9oFRI1G2/04EdgBd
L0feOOvDpxt3l9ZYdKyK73eV/tP76RJy0gr62BYPbi8OI9NrlV3Rqyyb0ELJVGbKVpnnBaxJs0mF
njpT9FIA7d1yAC1NS1XjMnuLuRIdBLui8MoU2xZdX4mRxhD63OQ5jNZBjJ6ijva8+2VCov78kAPL
gjFfRY8FRLm8NzBQpCya9enXemk49e1cb9VO+oi9KlUxwJMt4giBNMzryjmMjk3MR9JeJ77wFMCn
epxGb3huPT8UVDdPUfoQ2zVos/a1sx4kWVFdod9mESdfo6UoMjgUtLEQ1AMTimNCMjC9jW7Ee6dS
fQgiOHyZ4w5CbCTeGGyVqztVYsRkbPrUwp7iPQQRiZazi7s0T5AivaZx0+JbqVl7o+P+8krWkMia
n+T7HQELPEeBSXfU0IbDIUuuesZPiQgmJFaRoL/FoLQepyWPGyxhmplXvgpUjTItLA8yLNhspYXy
72xe8475BY/TirorvzxmOxWQm5B2ky4qohvQ8J847hffd7tB98ozewpyiDZTZwKuiUJJ3rFhMjiF
ZraURxmPtC/FbVKc46N6eSKybrHNMH9MYu4PsymQPjZxmzj/EgS9JMeNKu30+NBOT5ghEeicOif+
t1MVPXMo6kgMPnShw5uTblLPNLazIzlTmbpYgwo0hGcOQ9VEbiIAPHumXP95Z8v/CECzIfjZc1tm
JIrlShp3SW5B/YawGEfFhtWvRrfAjoGcr14a98EaRdrpYcPTlpZ25sMbg3cKMBPVyR+RutfOnFnk
mhH7JIjnvPGJ8lpZq/JAHtC+ZMBFKnr4S0wjthkZUAXMxqzw8oUM9dhREFn0+Vg5f+on82cFZctt
9plPO62sueVKIfQI343OKxtqDwjtAHCIuvNsMuPRPTDFc2vL9MSJZxP1pZFIu5JWtng5aEJ94F4S
zfhjPKqbcPaH8F02DwWM7MwImzOvpJGmfFz088a89CqMK8lV2DMLJyiy64EV6jKaYZj7omjIvZS/
psDO4UDIEJHcXxkKZf6hIJLI6CzfQUGpu9Wn+A8E4J6AP9fiqsGNE7EkXUxEK+ZlAVd4cTfDScGz
iUQgl+ectMZ4hT//TumkJSaRPKtUFtxtHJMOrRnNI/9TQq7KwNo8tia0ji0mqwylWU2vp3wNV8BN
BGr8pb86zinaEegRtnKXIripbSRehHa/rEudgkO1jUAe308wXsTmQs7bV1Zt3UA/QHFDKt8grsWM
hoUftrSEsCSOmhdXsMoyRQDJwWBM4SEWRo0Z4qfaRBd+rQmSaxorH/Umn76dsJr0K/g6g8Vzmkqn
7S6wcbYdV0716ekXbC8x4aDl3fHrhAXvR2d+TcFmJMI/kBSHRaT/4dLriahy/P4TJJXlUxH/Sig5
NBBHG8A84ddhbcl8flOJDUD4ZK1pI8fgGGjDlsMWemNx8OMkcSjXlwKN5WLhr87CVPHQP1TMZmWq
kvKU+nQ+TLjBgU3SCx1x0/p5TajBoCow0aGt78Q0Qe5NRllEgb+vT4XIa4dz73iSs5bJUKt1YtdH
vRTmv5SnBKG4evstBnPwrGhCLOYnj4bHcZAARkc0LnRU/EAgUkjwv5rLSvy5a9gvHqMhi6kDjYOZ
3hzSVk3QdMM1dIS5oYl4lhTW6vbba5kImL1UUVHLv0PJnaO/j9athsnqvFmf2nS3hb9kJdoKA0M1
8Wu7F4g4ZySvRVAXQibjo7lEFGQzX4ztMKhivdu42rwIglBNdQYqeCkIY0l5PiEhdnSnVPdAOb9A
ofS0ey+CRIpGewaCiDig43mHT3Utii3y/MXgt8gKNPL3j0EcgoplXUs8617xmOoas+n1dYRjxlBN
PspiS17uOsl2s7Mh9wV8t2dp6ATbEgM2tfCnLZFj/SptIEpLh1zhp+4ljancL9tu2Z/3g31kmmTR
DbjnalA4MNJYHpX1E5e0IpDOHBZz5kg5l0/fo//Pl2yIIokDHFgRAnY6ounYDfXbDHxVfSgpiZ9W
3fmfZqKq32abYKRoeaqfNlP4pxtJwsubXiRPQlhkfBStxuQjxhoTjz2ty8yTWb8hn8m9iINDgti5
GsJRIZu8t140DiX/84hfsOfzxzbJDWtFhfbOZPeLo3zFxbUqezd2LFTAUFyCE77ZqZbnr0YA5dCZ
7498Ww0z5ElZeVlgG4jbadGzqtEyl2PYCjVsRoT2Rr8jIC8zeuxPtcxY8CNSNod+Io7BBDM/Q7Lb
Nh1Scu+O1uEfTCH/vvueKTO7sXngtdob8IDWuUavZZ9MXZ9BkAUILKYOhuP2tngEpjaWIIIJBr+s
LPdQIAU1v/KaWtcpy3wutNInKUW9cxI4IyGXlxWXc/x0ewG8RcaK9zV4liCl0n+XN4klqSwIeStv
6vj3MRBuOAJp/ueSiTh7TB/t1Pg5YO6MYqnHEDr/pljZZI8GkvguVs92RS/CYzKqvdNL4TKjqMN8
iW29WdigTf5mZ53kviPzLPx3dM2D1dzTqX1EnhzPQKI4utR8ScE7D5Wx3tTgt4RLPZiQeHbpgB4H
7osj/Y1qTHcOYFUP9YVp2F4no6JsQrpLMYBCHrGILZaYVG02gXqSqUUbD9PDmZjossZx7i35fhJh
XTGrkr86PL8CoSJKrwOttmxsLJrTUgkh3pIxC7Bz5YIbP7TbRWXpPNIsd3/G2zZYiq2SskXFtAgS
X+8sosnXBl8y52OWawmQq1Ar5GE+F9YmuMAleniZaaS0O2Z47eGG15sKdNMNdTPB6lexCaSE1gDu
l/8kg9423AUfYUY3eAgR/jpKjxXyeRDhaBDeNCKl4oJvoQaBUR+itMlamyGB2GFRXrd7RwUwdmgX
dycXCXejZt6dAZVFQy8G9OhpFQyctKMVQtFc9CYedROXQIiCupEbR5hUfXOTPVw8/EABkdMKHRck
23scQHH46p6z2EoHPz9Js07+2qxeKdtJJNBWhIXkjHAfjigp3tlYv3gqsi98n8h8arCfgBoGGx8V
dNa0y7pPQ44Y0/9ju4mDf1SF1wZb3m5C1KvVr4rAlaD0DeDCn6vuXjWw8Y3uSaXEivdJ3ObMSsmD
4zQhecu7tSEhsut61uewSSSThP0zV9zIPd/tfXqfS4RvIKU5Gn39v2Y7IJpOsWOA4Opy2GH4gXoi
raVueQykqazrFvlEg30v9E+MIym/JmNuSmnRArdIoa8dHOYab73Pr50Avvveeh+OYIzCw69hZBan
eMsLH2VVI/LbtwKhpZX4hnpiHSo9MsE8ebEfbIH5XPU1l90vsYlbqiZBXcs13T3HvlUNeooZCLyI
Q6zhpImR66xqE0/QSxfJlmMj3I0cH7wP6bBXc2O1kJIYmsDNemRLqhqGI3olDTMGoueML9kYS0eV
mJgWmDFSQxBqMhOEYxmijXugUjTTxAhJi8Kjcv6R5RmhsqSTWvG8kaSOS2XgjO3LRoJ6BJyffWMi
2n9umn4b12NUy8PhvztIqmwRh09PZ0mDWBi+b1jU5X8UfD81tP615al+I8RZzv5K0e7hmaPO9WM/
Zb3fyme5H9dDRxKpOqiISErWww6lBPy4lh50ID7segCeIKh3sVsGCIof+G+H0+hrgApSJ+QMXh7M
Mvnlg3CH9rb41jxmzXtw15fK17/NbH07gLRwE7FTIi56+6EslfkzDhc+Hqz+M7UGJDdtuHfcA/J1
wPNDCGziLYB5eCWWMZtJnlBAddS7RLat6GW+iCYApff5WwyJjjuETPSMdmgLOljJp9GoxvJ9Ikwu
Dii7ZZ4F2Mu4XjwohFW/+rVh6uszgwjBpAd9FJOAJV+zD+InAFstJ/wgcSwL8LILjKoVudmy6G8+
55HXsaddjpryNgpSjvj/xS3itdADMuhwFEWHbyD8GCkN24DMkTUjisrGzwORIlMiQuXzPgt5/5QP
GFZK1944hMuENYP2RedQVuS8s2qQ9GoAEqma5nPSYbhkrdSsZOHjwa+Gr4P09hkmDTGXxFXYxhjO
Bhwhdykd+R4K8hOEQdbCw9jz2lyj2nSCfK1hEM7qsEhQt1AvhS6wcprbVJBuYY0/d3eZ9DUCRxoq
nlZja9Y71JgxN7kWYWVcFEDsaTQlx1hi50Dk6cIuEUiztlZNhkcna1cQPqjZprucOmy7tVjb0oeP
ec/7KokpQ/va7vGpuR0hhEToM4Hd6P3/8YK3Xnqq2VSFb22VaD4wLO9bmQcqntdJJt4L1h7CqQ9I
WnnoacjFByqXCt9q225xZ69YIpbX3VOAqVu78De/6C/soVKOTP0D07yOT59PtUzHODBSJjkeKIPn
3u2nbjodB+H3WmGUwZVRbxNPmWYJYma2CyxzO/EO10QPyNns+138XjSu+bZtrF6Ql0PjCrT0F1gz
KizUnnLIgL3XeiRn0X2NomWGty8GaAdkdMZXb7uHNdN1Z+Y/k661/WwgOqDH8od7egAN7VnU3UbP
jBzPzPjKwJlX3kJBHnPmgnIDadxhn97uDvzgLaiDTJv8DpS8yBb5EUlgdnyGzOz/7n/WIdNsGGZ8
rtP+ZLh8/9AoFWOTw91JBRklucK+qFyOxdWtY56YPadX7bSRn6IQrgo/5SM9+n1utpGyBYiyNN+r
N1PMw3MU240tbSo19vBiDZf2wboeMoVEi463JaTYAMml3c27RRy1PdVvkp68R0TvZX2Fe9jashy3
ARe35o4kMVHWQ/L3u0qSAEFddD6Emcgd/G2UzYWx+hPRqR3DPBU5PiNhO+1aL26dzkvsbZJi27pk
2qvk2wJn84sAOSnYSC05au0ds28tt8ACKKVCSSirP1yobUsCtlXszMD5uziquz22r2PmMSJgtg1O
lumGvTe7zUs6QFjLbuxNHcRO4viAkQfw5GuYIPlp1F00I0LvLIMPxy+KejYAeQK+1bMTT8Y02IB+
Gikn1t43tQ1Rsdejjkij1Bw2ie2PWQY2nryInWNrfX5vUzKUiMy/rUaeUtIzdf82LValkDo48krI
4tlBiUoGusQz3ud2QTB756Fr2BxN2kq03wIHKQMVP8GP0lLxqH0viNWow4rvy6imyOP01i0fpQ7a
uVOghfviAWbyJY/lEcqoR7/ZpYe7uaOSVrZCkyUhyxS4ocuIodwVOpGDj1UuLFq1B2xRvp/i1hIo
enLfHQtU8A0OGJd7jkE1lHYcmSuICTdO9I+bd868d226+THBIK7Ds97lpjjkFok/bj6DO6MGVuex
VepirFIfVLRO+aIPjHlx4j/lqrMXrc155eD1uXp3t90bcq4QwJuJIZIadUKf3ZYynqBoZ7rSIwSt
Q5DBa6sUcWpXs6UmDJad2kAv0gC+ozioDpUV8B5gNusE28lQO+5BU6r4snEIT8l7Feh8D/Pp7wxw
bxOA11fkgkqvbNpmQndbl7IZeD+4SBL206c6nUlEdiy48PA/WLIEZ/3Wt/CB+CKhEmoDbgsthC/X
qF3SQSkADQCDRaWckoqc22G6GG0iZ8ct1cpGyuSTJGRp07PMNYVyqruQDVL+e2q8CvSd8hmBAO+m
GRONMaDOe1RZEe8PUNaaBMdpsxpC8cqpeqhgg/rOoauYP0js1C2BOcpgV6jI0kTw1HC+53KfYHz2
Hu+ZB6TJJXHgDWS0iQMoGBhuouRRhamv/KfSwSN18pGrfDoIjYXKG5O3Dn0/HsZQfTkbRDNR2oNB
WOLSEN3zry8tVXbVjICm2BijK/qrr56q8fo9//qXfWpK0JntQOXfWj38/OJySt9dkYe/HHRHragH
G0NrKPXYegs4mrevRRhtsnk+7WFtlefIAVNL5fX7oo3JPiUHOLyup2fd3iRvVsK4ZEoB7L/5CDvF
fr6op+iPfzkTUor7o4X514A64JQyMf9t92Ox9D8PCTnCDWka01ncjNsEvmrsDbyaPvXl1FKOrwzH
fdHik8AAnknaX8IjTIAnzC+LoY5xaN0pr4V5zpU57j4oS9N9ARmZxD89INrDKNtbs2BB3fGYOq5D
eriJOe7wsB7g+yW10ml+jlwn5ptHsHimxcwo7ikAPr+LQI7P65FlLMgqtkgiNE1ZMQyyrCGmi2xc
AS9BWur5QoIgpXwKlVPYJ6ME+kYHtw60tnkBz+UxEBQcEXW2RArqT1ZvLPkbov7Atx6XcREb/qKm
vgdJ4z90Gw1s0QTBYsHadgcrQfQeuLlpiJHpCQ8QuL2inI6xhGOI8OAw8hQx19NvocHZwoeXmj7x
mUewsCL37cstOFam9mAHwGe7zl2y+OsmhSGTPv2scViJs47j9KBRFlDkmXg7kkgPqf1f96+sYjcO
nfK7u+VbhkBTZqViq6fcXWPpxlVWEihQrtwVh9nh7niwy6qd5+VHwwH103RndIRNg4Tvx6Fd6ck2
39EmClTAcVWiw7Y7AJ5tY86PoV+92CkaQ8n5BKGdFPSqep0FDlVTRFmhrxvdozqlBC/+EsrvgkM6
kNm6JwiFoqGVZC/TjlXGDd8YCKrocv5hPTpn1vIoaxXVZXLrm1/IRISn8r7Qx36f3bQEHc0iQKtv
0jXaSotbV0bbdJOSGGiutEs1iNSlfHVLFNNqziLzVhGq05dB8cFK35mvW4GReN1exdE4c0dNbFrf
gJmArLZMeApFiWeJTDRsBBhNLsA8SFlzEnXKSXE7Pd7FbshdtxF9t908E/76EK8VXnvMBCkLqrvR
FloGerYKn02KZRvhDhst6oMkwOSmaLyWO4JA39ojxDvbCl388zQ8/aHNIcpEfTwHY+/hF13ooGIG
U2faaXf8IUDsYIYw7egmlahR8mkFYr8CmTJeQiFpezAhGww9GDe3Ug0I360VThdssb50xQ6YonKf
y63rdjyeDeSJIkaAQjhaPi0lnGaZnPYiDAU1O0SQNKHWd0H630/K9Oj9TiYp/8uydhZR01jkwRMx
aPP0ouwfLawELKEoP69zvks6q1D4FnZtSr6LnFuJZb261OHtHOCCBObRU8zbUmSVSCSN92rvN3yd
2zC31MM+AkAIqOaWC/TVNf6ssEiHOPF6NtMqocpNkKW+T3reB8GMS8k7OyTIN7MaOlHlrr2ejsbf
qHBqsQ6e0hjnQCt+4UQHZSc2x8jEyjQNyNCbxrj6h36KX84XnPRY7o3Rw/PlC5t/5Rnuz8tJp4SA
6EHeStDmTIu6ofl7Ag5YMby0Uq548VfOldYFzFcgLusXZRf0R7jIHO5Utm3Phsqsd26qOmLX1XGg
xk8JJ6nURf9KAP+YDg0VkJhQc4tx2VqwxMCJ/Iunqm62c7QWnUyCEjuc7D3UaIlrJn0kvc2lQGCh
hNTjx+oGNIE2vban3QCBNXMk+R5IN+nx07E/CG6K1ns1RnrE6OYS6JqD3n3PU1CHnUAArafNgMNt
wnwJMMncg2P2aNFpckkvqlekVgqUe/v3Xe8xXfVh/RQAXnomdwFMPwUUFM4KpOaewM2X45QJKe6y
0oBi7lTCy6FFAzmxsenNjpGA8fV9kKGmIxUHDmRaa2Q8AEMSvW+2Vmism7ataK/y9TNnnvwnHByy
NLxdt7CC7CelvDnEP8Uk7OhF5s26/glIvavgTe1DGcbmhM7Xny4C9jSgoxVsbzP//QP9P2KNAQDH
Psx1DQ+n1lTvzNkfHL2a10YcSgwYgSHkkP3bdefJB0ncjGnnq7uMX6oFU2RHe/tRz415ZmHqnxAY
6zXr5hmg5gxnMahiVpLDOWy3D1+MK8xpUC0ke7Wryz41EDUySNlH3tdGq0YMwxKM/iSONkfeB11p
UKnd/qoOnRBEKNHken1uvzhW0SWsl7ndu4SGr7yQ5zwsHmG9wye9X7v0csbVEE0bOLKMoXs=
`protect end_protected
